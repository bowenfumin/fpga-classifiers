module lut_5level_tree3(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [576:0] data_in,
                       input       data_valid,
                       output      data_out     
                       );
wire    [576:0] InputBits;
wire    gates_1, gates_2, gates_3, gates_4, gates_5, gates_6, gates_7, gates_8, gates_9, gates_10, gates_11, gates_12, gates_13, gates_14, gates_15, gates_16, gates_17, gates_18, gates_19, gates_20, gates_21, gates_22, gates_23, gates_24, gates_25, gates_26, gates_27, gates_28, gates_29, gates_30, gates_31, gates_32, gates_33, gates_34, gates_35, gates_36, gates_37, gates_38, gates_39, gates_40, gates_41, gates_42, gates_43, gates_44, gates_45, gates_46, gates_47, gates_48, gates_49, gates_50, gates_51, gates_52, gates_53, gates_54, gates_55, gates_56, gates_57, gates_58, gates_59, gates_60, gates_61, gates_62, gates_63, gates_64, gates_65, gates_66, gates_67, gates_68, gates_69, gates_70, gates_71, gates_72, gates_73, gates_74, gates_75, gates_76, gates_77, gates_78, gates_79, gates_80, gates_81, gates_82, gates_83, gates_84, gates_85, gates_86, gates_87, gates_88, gates_89, gates_90, gates_91, gates_92, gates_93, gates_94, gates_95, gates_96, gates_97, gates_98, gates_99, gates_100, gates_101, gates_102, gates_103, gates_104, gates_105, gates_106, gates_107, gates_108, gates_109, gates_110, gates_111, gates_112, gates_113, gates_114, gates_115, gates_116, gates_117, gates_118, gates_119, gates_120, gates_121, gates_122, gates_123, gates_124, gates_125, gates_126, gates_127, gates_128, gates_129, gates_130, gates_131, gates_132, gates_133, gates_134, gates_135, gates_136, gates_137, gates_138, gates_139, gates_140, gates_141, gates_142, gates_143, gates_144, gates_145, gates_146, gates_147, gates_148, gates_149, gates_150, gates_151, gates_152, gates_153, gates_154, gates_155, gates_156, gates_157, gates_158, gates_159, gates_160, gates_161, gates_162, gates_163, gates_164, gates_165, gates_166, gates_167, gates_168, gates_169, gates_170, gates_171, gates_172, gates_173, gates_174, gates_175, gates_176, gates_177, gates_178, gates_179, gates_180, gates_181, gates_182, gates_183, gates_184, gates_185, gates_186, gates_187, gates_188, gates_189, gates_190, gates_191, gates_192, gates_193, gates_194, gates_195, gates_196, gates_197, gates_198, gates_199, gates_200, gates_201, gates_202, gates_203, gates_204, gates_205, gates_206, gates_207, gates_208, gates_209, gates_210, gates_211, gates_212, gates_213, gates_214, gates_215, gates_216, gates_217, gates_218, gates_219, gates_220, gates_221, gates_222, gates_223, gates_224, gates_225, gates_226, gates_227, gates_228, gates_229, gates_230, gates_231, gates_232, gates_233, gates_234, gates_235, gates_236, gates_237, gates_238, gates_239, gates_240, gates_241, gates_242, gates_243, gates_244, gates_245, gates_246, gates_247, gates_248, gates_249, gates_250, gates_251, gates_252, gates_253, gates_254, gates_255, gates_256, gates_257, gates_258, gates_259, gates_260, gates_261, gates_262, gates_263, gates_264, gates_265, gates_266, gates_267, gates_268, gates_269, gates_270, gates_271, gates_272, gates_273, gates_274, gates_275, gates_276, gates_277, gates_278, gates_279, gates_280, gates_281, gates_282, gates_283, gates_284, gates_285, gates_286, gates_287, gates_288, gates_289, gates_290, gates_291, gates_292, gates_293, gates_294, gates_295, gates_296, gates_297, gates_298, gates_299, gates_300, gates_301, gates_302, gates_303, gates_304, gates_305, gates_306, gates_307, gates_308, gates_309, gates_310, gates_311, gates_312, gates_313, gates_314, gates_315, gates_316, gates_317, gates_318, gates_319, gates_320, gates_321, gates_322, gates_323, gates_324, gates_325, gates_326, gates_327, gates_328, gates_329, gates_330, gates_331, gates_332, gates_333, gates_334, gates_335, gates_336, gates_337, gates_338, gates_339, gates_340, gates_341, gates_342, gates_343, gates_344, gates_345, gates_346, gates_347, gates_348, gates_349, gates_350, gates_351, gates_352, gates_353, gates_354, gates_355, gates_356, gates_357, gates_358, gates_359, gates_360, gates_361, gates_362, gates_363, gates_364, gates_365, gates_366, gates_367, gates_368, gates_369, gates_370, gates_371, gates_372, gates_373, gates_374, gates_375, gates_376, gates_377, gates_378, gates_379, gates_380, gates_381, gates_382, gates_383, gates_384, gates_385, gates_386, gates_387, gates_388, gates_389, gates_390, gates_391, gates_392, gates_393, gates_394, gates_395, gates_396, gates_397, gates_398, gates_399, gates_400, gates_401, gates_402, gates_403, gates_404, gates_405, gates_406, gates_407, gates_408, gates_409, gates_410, gates_411, gates_412, gates_413, gates_414, gates_415, gates_416, gates_417, gates_418, gates_419, gates_420, gates_421, gates_422, gates_423, gates_424, gates_425, gates_426, gates_427, gates_428, gates_429, gates_430, gates_431, gates_432, gates_433, gates_434, gates_435, gates_436, gates_437, gates_438, gates_439, gates_440, gates_441, gates_442, gates_443, gates_444, gates_445, gates_446, gates_447, gates_448, gates_449, gates_450, gates_451, gates_452, gates_453, gates_454, gates_455, gates_456, gates_457, gates_458, gates_459, gates_460, gates_461, gates_462, gates_463, gates_464, gates_465, gates_466, gates_467, gates_468, gates_469, gates_470, gates_471, gates_472, gates_473, gates_474, gates_475, gates_476, gates_477, gates_478, gates_479, gates_480, gates_481, gates_482, gates_483, gates_484, gates_485, gates_486, gates_487, gates_488, gates_489, gates_490, gates_491, gates_492, gates_493, gates_494, gates_495, gates_496, gates_497, gates_498, gates_499, gates_500, gates_501, gates_502, gates_503, gates_504, gates_505, gates_506, gates_507, gates_508, gates_509, gates_510, gates_511, gates_512, gates_513, gates_514, gates_515, gates_516, gates_517, gates_518, gates_519, gates_520, gates_521, gates_522, gates_523, gates_524, gates_525, gates_526, gates_527, gates_528, gates_529, gates_530, gates_531, gates_532, gates_533, gates_534, gates_535, gates_536, gates_537, gates_538, gates_539, gates_540, gates_541, gates_542, gates_543, gates_544, gates_545, gates_546, gates_547, gates_548, gates_549, gates_550, gates_551, gates_552, gates_553, gates_554, gates_555, gates_556, gates_557, gates_558, gates_559, gates_560, gates_561, gates_562, gates_563, gates_564, gates_565, gates_566, gates_567, gates_568, gates_569, gates_570, gates_571, gates_572, gates_573, gates_574, gates_575, gates_576, gates_577, gates_578, gates_579, gates_580, gates_581, gates_582, gates_583, gates_584, gates_585, gates_586, gates_587, gates_588, gates_589, gates_590, gates_591, gates_592, gates_593, gates_594, gates_595, gates_596, gates_597, gates_598, gates_599, gates_600, gates_601, gates_602, gates_603, gates_604, gates_605, gates_606, gates_607, gates_608, gates_609, gates_610, gates_611, gates_612, gates_613, gates_614, gates_615, gates_616, gates_617, gates_618, gates_619, gates_620, gates_621, gates_622, gates_623, gates_624, gates_625, gates_626, gates_627, gates_628, gates_629, gates_630, gates_631, gates_632, gates_633, gates_634, gates_635, gates_636, gates_637, gates_638, gates_639, gates_640, gates_641, gates_642, gates_643, gates_644, gates_645, gates_646, gates_647, gates_648, gates_649, gates_650, gates_651, gates_652, gates_653, gates_654, gates_655, gates_656, gates_657, gates_658, gates_659, gates_660, gates_661, gates_662, gates_663, gates_664, gates_665, gates_666, gates_667, gates_668, gates_669, gates_670, gates_671, gates_672, gates_673, gates_674, gates_675, gates_676, gates_677, gates_678, gates_679, gates_680, gates_681, gates_682, gates_683, gates_684, gates_685, gates_686, gates_687, gates_688, gates_689, gates_690, gates_691, gates_692, gates_693, gates_694, gates_695, gates_696, gates_697, gates_698, gates_699, gates_700, gates_701, gates_702, gates_703, gates_704, gates_705, gates_706, gates_707, gates_708, gates_709, gates_710, gates_711, gates_712, gates_713, gates_714, gates_715, gates_716, gates_717, gates_718, gates_719, gates_720, gates_721, gates_722, gates_723, gates_724, gates_725, gates_726, gates_727, gates_728, gates_729, gates_730, gates_731, gates_732, gates_733, gates_734, gates_735, gates_736, gates_737, gates_738, gates_739, gates_740, gates_741, gates_742, gates_743, gates_744, gates_745, gates_746, gates_747, gates_748, gates_749, gates_750, gates_751, gates_752, gates_753, gates_754, gates_755, gates_756, gates_757, gates_758, gates_759, gates_760, gates_761, gates_762, gates_763, gates_764, gates_765, gates_766, gates_767, gates_768, gates_769, gates_770, gates_771, gates_772, gates_773, gates_774, gates_775, gates_776, gates_777, gates_778, gates_779, gates_780, gates_781, gates_782, gates_783, gates_784, gates_785, gates_786, gates_787, gates_788, gates_789, gates_790, gates_791, gates_792, gates_793, gates_794, gates_795, gates_796, gates_797, gates_798, gates_799, gates_800, gates_801, gates_802, gates_803, gates_804, gates_805, gates_806, gates_807, gates_808, gates_809, gates_810, gates_811, gates_812, gates_813, gates_814, gates_815, gates_816, gates_817, gates_818, gates_819, gates_820, gates_821, gates_822, gates_823, gates_824, gates_825, gates_826, gates_827, gates_828, gates_829, gates_830, gates_831, gates_832, gates_833, gates_834, gates_835, gates_836, gates_837, gates_838, gates_839, gates_840, gates_841, gates_842, gates_843, gates_844, gates_845, gates_846, gates_847, gates_848, gates_849, gates_850, gates_851, gates_852, gates_853, gates_854, gates_855, gates_856, gates_857, gates_858, gates_859, gates_860, gates_861, gates_862, gates_863, gates_864, gates_865, gates_866, gates_867, gates_868, gates_869, gates_870, gates_871, gates_872, gates_873, gates_874, gates_875, gates_876, gates_877, gates_878, gates_879, gates_880, gates_881, gates_882, gates_883, gates_884, gates_885, gates_886, gates_887, gates_888, gates_889, gates_890, gates_891, gates_892, gates_893, gates_894, gates_895, gates_896, gates_897, gates_898, gates_899, gates_900, gates_901, gates_902, gates_903, gates_904, gates_905, gates_906, gates_907, gates_908, gates_909, gates_910, gates_911, gates_912, gates_913, gates_914, gates_915, gates_916, gates_917, gates_918, gates_919, gates_920, gates_921, gates_922, gates_923, gates_924, gates_925, gates_926, gates_927, gates_928, gates_929, gates_930, gates_931, gates_932, gates_933, gates_934, gates_935, gates_936, gates_937, gates_938, gates_939, gates_940, gates_941, gates_942, gates_943, gates_944, gates_945, gates_946, gates_947, gates_948, gates_949, gates_950, gates_951, gates_952, gates_953, gates_954, gates_955, gates_956, gates_957, gates_958, gates_959, gates_960, gates_961, gates_962, gates_963, gates_964, gates_965, gates_966, gates_967, gates_968, gates_969, gates_970, gates_971, gates_972, gates_973, gates_974, gates_975, gates_976, gates_977, gates_978, gates_979, gates_980, gates_981, gates_982, gates_983, gates_984, gates_985, gates_986, gates_987, gates_988, gates_989, gates_990, gates_991, gates_992, gates_993, gates_994, gates_995, gates_996, gates_997, gates_998, gates_999, gates_1000, gates_1001, gates_1002, gates_1003, gates_1004, gates_1005, gates_1006, gates_1007, gates_1008, gates_1009, gates_1010, gates_1011, gates_1012, gates_1013, gates_1014, gates_1015, gates_1016, gates_1017, gates_1018, gates_1019, gates_1020, gates_1021, gates_1022, gates_1023, gates_1024, gates_1025, gates_1026, gates_1027, gates_1028, gates_1029, gates_1030, gates_1031, gates_1032, gates_1033, gates_1034, gates_1035, gates_1036, gates_1037, gates_1038, gates_1039, gates_1040, gates_1041, gates_1042, gates_1043, gates_1044, gates_1045, gates_1046, gates_1047, gates_1048, gates_1049, gates_1050, gates_1051, gates_1052, gates_1053, gates_1054, gates_1055, gates_1056, gates_1057, gates_1058, gates_1059, gates_1060, gates_1061, gates_1062, gates_1063, gates_1064, gates_1065, gates_1066, gates_1067, gates_1068, gates_1069, gates_1070, gates_1071, gates_1072, gates_1073, gates_1074, gates_1075, gates_1076, gates_1077, gates_1078, gates_1079, gates_1080, gates_1081, gates_1082, gates_1083, gates_1084, gates_1085, gates_1086, gates_1087, gates_1088, gates_1089, gates_1090, gates_1091, gates_1092, gates_1093, gates_1094, gates_1095, gates_1096, gates_1097, gates_1098, gates_1099, gates_1100, gates_1101, gates_1102, gates_1103, gates_1104, gates_1105, gates_1106, gates_1107, gates_1108, gates_1109, gates_1110, gates_1111, gates_1112, gates_1113, gates_1114, gates_1115, gates_1116, gates_1117, gates_1118, gates_1119, gates_1120, gates_1121, gates_1122, gates_1123, gates_1124, gates_1125, gates_1126, gates_1127, gates_1128, gates_1129, gates_1130, gates_1131, gates_1132, gates_1133, gates_1134, gates_1135, gates_1136, gates_1137, gates_1138, gates_1139, gates_1140, gates_1141, gates_1142, gates_1143, gates_1144, gates_1145, gates_1146, gates_1147, gates_1148, gates_1149, gates_1150, gates_1151, gates_1152, gates_1153, gates_1154, gates_1155, gates_1156, gates_1157, gates_1158, gates_1159, gates_1160, gates_1161, gates_1162, gates_1163, gates_1164, gates_1165, gates_1166, gates_1167, gates_1168, gates_1169, gates_1170, gates_1171, gates_1172, gates_1173, gates_1174, gates_1175, gates_1176, gates_1177, gates_1178, gates_1179, gates_1180, gates_1181, gates_1182, gates_1183, gates_1184, gates_1185, gates_1186, gates_1187, gates_1188, gates_1189, gates_1190, gates_1191, gates_1192, gates_1193, gates_1194, gates_1195, gates_1196, gates_1197, gates_1198, gates_1199, gates_1200, gates_1201, gates_1202, gates_1203, gates_1204, gates_1205, gates_1206, gates_1207, gates_1208, gates_1209, gates_1210, gates_1211, gates_1212, gates_1213, gates_1214, gates_1215, gates_1216, gates_1217, gates_1218, gates_1219, gates_1220, gates_1221, gates_1222, gates_1223, gates_1224, gates_1225, gates_1226, gates_1227, gates_1228, gates_1229, gates_1230, gates_1231, gates_1232, gates_1233, gates_1234, gates_1235, gates_1236, gates_1237, gates_1238, gates_1239, gates_1240, gates_1241, gates_1242, gates_1243, gates_1244, gates_1245, gates_1246, gates_1247, gates_1248, gates_1249, gates_1250, gates_1251, gates_1252, gates_1253, gates_1254, gates_1255, gates_1256, gates_1257, gates_1258, gates_1259, gates_1260, gates_1261, gates_1262, gates_1263, gates_1264, gates_1265, gates_1266, gates_1267, gates_1268, gates_1269, gates_1270, gates_1271, gates_1272, gates_1273, gates_1274, gates_1275, gates_1276, gates_1277, gates_1278, gates_1279, gates_1280, gates_1281, gates_1282, gates_1283, gates_1284, gates_1285, gates_1286, gates_1287, gates_1288, gates_1289, gates_1290, gates_1291, gates_1292, gates_1293, gates_1294, gates_1295, gates_1296, gates_1297, gates_1298, gates_1299, gates_1300, gates_1301, gates_1302, gates_1303, gates_1304, gates_1305, gates_1306, gates_1307, gates_1308, gates_1309, gates_1310, gates_1311, gates_1312, gates_1313, gates_1314, gates_1315, gates_1316, gates_1317, gates_1318, gates_1319, gates_1320, gates_1321, gates_1322, gates_1323, gates_1324, gates_1325, gates_1326, gates_1327, gates_1328, gates_1329, gates_1330, gates_1331, gates_1332, gates_1333, gates_1334, gates_1335, gates_1336, gates_1337, gates_1338, gates_1339, gates_1340, gates_1341, gates_1342, gates_1343, gates_1344, gates_1345, gates_1346, gates_1347, gates_1348, gates_1349, gates_1350, gates_1351, gates_1352, gates_1353, gates_1354, gates_1355, gates_1356, gates_1357, gates_1358, gates_1359, gates_1360, gates_1361, gates_1362, gates_1363, gates_1364, gates_1365, gates_1366, gates_1367, gates_1368, gates_1369, gates_1370, gates_1371, gates_1372, gates_1373, gates_1374, gates_1375, gates_1376, gates_1377, gates_1378, gates_1379, gates_1380, gates_1381, gates_1382, gates_1383, gates_1384, gates_1385, gates_1386, gates_1387, gates_1388, gates_1389, gates_1390, gates_1391, gates_1392, gates_1393, gates_1394, gates_1395, gates_1396, gates_1397, gates_1398, gates_1399, gates_1400, gates_1401, gates_1402, gates_1403, gates_1404, gates_1405, gates_1406, gates_1407, gates_1408, gates_1409, gates_1410, gates_1411, gates_1412, gates_1413, gates_1414, gates_1415, gates_1416, gates_1417, gates_1418, gates_1419, gates_1420, gates_1421, gates_1422, gates_1423, gates_1424, gates_1425, gates_1426, gates_1427, gates_1428, gates_1429, gates_1430, gates_1431, gates_1432, gates_1433, gates_1434, gates_1435, gates_1436, gates_1437, gates_1438, gates_1439, gates_1440, gates_1441, gates_1442, gates_1443, gates_1444, gates_1445, gates_1446, gates_1447, gates_1448, gates_1449, gates_1450, gates_1451, gates_1452, gates_1453, gates_1454, gates_1455, gates_1456, gates_1457, gates_1458, gates_1459, gates_1460, gates_1461, gates_1462, gates_1463, gates_1464, gates_1465, gates_1466, gates_1467, gates_1468, gates_1469, gates_1470, gates_1471, gates_1472, gates_1473, gates_1474, gates_1475, gates_1476, gates_1477, gates_1478, gates_1479, gates_1480, gates_1481, gates_1482, gates_1483, gates_1484, gates_1485, gates_1486, gates_1487, gates_1488, gates_1489, gates_1490, gates_1491, gates_1492, gates_1493, gates_1494, gates_1495, gates_1496, gates_1497, gates_1498, gates_1499, gates_1500, gates_1501, gates_1502, gates_1503, gates_1504, gates_1505, gates_1506, gates_1507, gates_1508, gates_1509, gates_1510, gates_1511, gates_1512, gates_1513, gates_1514, gates_1515, gates_1516, gates_1517, gates_1518, gates_1519, gates_1520, gates_1521, gates_1522, gates_1523, gates_1524, gates_1525, gates_1526, gates_1527, gates_1528, gates_1529, gates_1530, gates_1531, gates_1532, gates_1533, gates_1534, gates_1535, gates_1536, gates_1537, gates_1538, gates_1539, gates_1540, gates_1541, gates_1542, gates_1543, gates_1544, gates_1545, gates_1546, gates_1547, gates_1548, gates_1549, gates_1550, gates_1551, gates_1552, gates_1553, gates_1554, gates_1555;

assign  InputBits = data_in;
//assign  data_out = data_valid & gates[807];
assign  data_out = data_valid & gates_1555;

LUT6 #(
   .INIT(64'b0101010001010001010101010101010101010100010101010001010100010101)  
) LUT6_1 (
   .O(gates_1),
   .I0(InputBits[97]),
   .I1(InputBits[131]),
   .I2(InputBits[277]),
   .I3(InputBits[155]),
   .I4(InputBits[408]),
   .I5(InputBits[384])
);
LUT6 #(
   .INIT(64'b0101000101110111001101110101001100100011000100110010011101000000)  
) LUT6_2 (
   .O(gates_2),
   .I0(InputBits[467]),
   .I1(InputBits[570]),
   .I2(InputBits[297]),
   .I3(InputBits[308]),
   .I4(InputBits[244]),
   .I5(InputBits[326])
);
LUT6 #(
   .INIT(64'b0000000100000101000000000000010101000000010000010101010001011101)  
) LUT6_3 (
   .O(gates_3),
   .I0(InputBits[565]),
   .I1(InputBits[138]),
   .I2(InputBits[93]),
   .I3(InputBits[228]),
   .I4(InputBits[230]),
   .I5(InputBits[480])
);
LUT6 #(
   .INIT(64'b0101010100000100010111010000010101010101000001010101011101001111)  
) LUT6_4 (
   .O(gates_4),
   .I0(InputBits[144]),
   .I1(InputBits[284]),
   .I2(InputBits[104]),
   .I3(InputBits[392]),
   .I4(InputBits[474]),
   .I5(InputBits[134])
);
LUT6 #(
   .INIT(64'b0000000000110101000000000001000100000000111101110000000000110001)  
) LUT6_5 (
   .O(gates_5),
   .I0(InputBits[106]),
   .I1(InputBits[386]),
   .I2(InputBits[440]),
   .I3(InputBits[97]),
   .I4(InputBits[236]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0000000000000000000101000100000000000000010000000101000101010000)  
) LUT6_6 (
   .O(gates_6),
   .I0(InputBits[558]),
   .I1(InputBits[375]),
   .I2(InputBits[342]),
   .I3(InputBits[239]),
   .I4(InputBits[52]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0000001100000011000000110000001000110111011101110010001100100111)  
) LUT6_7 (
   .O(gates_7),
   .I0(InputBits[117]),
   .I1(InputBits[9]),
   .I2(InputBits[251]),
   .I3(InputBits[413]),
   .I4(InputBits[443]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0001000100000100000100010000010000000001000001010001000100010101)  
) LUT6_8 (
   .O(gates_8),
   .I0(InputBits[19]),
   .I1(InputBits[384]),
   .I2(InputBits[543]),
   .I3(InputBits[245]),
   .I4(InputBits[133]),
   .I5(InputBits[490])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000010100000001000001110010)  
) LUT6_9 (
   .O(gates_9),
   .I0(InputBits[120]),
   .I1(InputBits[58]),
   .I2(InputBits[372]),
   .I3(InputBits[218]),
   .I4(InputBits[68]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0100010001001000010001010100010001010101010100000100010101010100)  
) LUT6_10 (
   .O(gates_10),
   .I0(InputBits[123]),
   .I1(InputBits[260]),
   .I2(InputBits[118]),
   .I3(InputBits[420]),
   .I4(InputBits[281]),
   .I5(InputBits[401])
);
LUT6 #(
   .INIT(64'b0000010101000101000000000101110100000111000101110000000001000010)  
) LUT6_11 (
   .O(gates_11),
   .I0(InputBits[288]),
   .I1(InputBits[209]),
   .I2(InputBits[569]),
   .I3(InputBits[132]),
   .I4(InputBits[372]),
   .I5(InputBits[176])
);
LUT6 #(
   .INIT(64'b0000111101000000000001010001000100000101000000000000001100110001)  
) LUT6_12 (
   .O(gates_12),
   .I0(InputBits[486]),
   .I1(InputBits[378]),
   .I2(InputBits[30]),
   .I3(InputBits[91]),
   .I4(InputBits[355]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010000101000000000000011110000101000001011)  
) LUT6_13 (
   .O(gates_13),
   .I0(InputBits[372]),
   .I1(InputBits[277]),
   .I2(InputBits[97]),
   .I3(InputBits[508]),
   .I4(InputBits[263]),
   .I5(InputBits[533])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000111011100000000000000000001000111000101)  
) LUT6_14 (
   .O(gates_14),
   .I0(InputBits[485]),
   .I1(InputBits[197]),
   .I2(InputBits[58]),
   .I3(InputBits[17]),
   .I4(InputBits[566]),
   .I5(InputBits[212])
);
LUT6 #(
   .INIT(64'b0000000100000000010101010001010100000000000000000101000000000100)  
) LUT6_15 (
   .O(gates_15),
   .I0(InputBits[51]),
   .I1(InputBits[165]),
   .I2(InputBits[477]),
   .I3(InputBits[139]),
   .I4(InputBits[338]),
   .I5(InputBits[319])
);
LUT6 #(
   .INIT(64'b0000000000001100000000100000011000001110010000000000010100000100)  
) LUT6_16 (
   .O(gates_16),
   .I0(InputBits[447]),
   .I1(InputBits[326]),
   .I2(InputBits[338]),
   .I3(InputBits[243]),
   .I4(InputBits[327]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0000000100000011000000000000001100000010000000110000000000000000)  
) LUT6_17 (
   .O(gates_17),
   .I0(InputBits[93]),
   .I1(InputBits[24]),
   .I2(InputBits[74]),
   .I3(InputBits[302]),
   .I4(InputBits[344]),
   .I5(InputBits[214])
);
LUT6 #(
   .INIT(64'b1000101100001101111111111101111100001010000000111010000001110000)  
) LUT6_18 (
   .O(gates_18),
   .I0(InputBits[346]),
   .I1(InputBits[381]),
   .I2(InputBits[334]),
   .I3(InputBits[347]),
   .I4(InputBits[384]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010101010100010101)  
) LUT6_19 (
   .O(gates_19),
   .I0(InputBits[409]),
   .I1(InputBits[172]),
   .I2(InputBits[331]),
   .I3(InputBits[358]),
   .I4(InputBits[475]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1000100011111111000010000111111100001100101011100000110000101110)  
) LUT6_20 (
   .O(gates_20),
   .I0(InputBits[442]),
   .I1(InputBits[212]),
   .I2(InputBits[257]),
   .I3(InputBits[228]),
   .I4(InputBits[450]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100010001000100010001)  
) LUT6_21 (
   .O(gates_21),
   .I0(InputBits[409]),
   .I1(InputBits[19]),
   .I2(InputBits[90]),
   .I3(InputBits[314]),
   .I4(InputBits[463]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000000000000000000011101111110100000000000010100000111111110100)  
) LUT6_22 (
   .O(gates_22),
   .I0(InputBits[184]),
   .I1(InputBits[375]),
   .I2(InputBits[92]),
   .I3(InputBits[431]),
   .I4(InputBits[570]),
   .I5(InputBits[357])
);
LUT6 #(
   .INIT(64'b0101010101010100010100010101000001110111010001000011011100000110)  
) LUT6_23 (
   .O(gates_23),
   .I0(InputBits[312]),
   .I1(InputBits[142]),
   .I2(InputBits[136]),
   .I3(InputBits[344]),
   .I4(InputBits[307]),
   .I5(InputBits[66])
);
LUT6 #(
   .INIT(64'b0001000000000000110110000001100000000000000100010111001011111111)  
) LUT6_24 (
   .O(gates_24),
   .I0(InputBits[498]),
   .I1(InputBits[503]),
   .I2(InputBits[453]),
   .I3(InputBits[127]),
   .I4(InputBits[12]),
   .I5(InputBits[126])
);
LUT6 #(
   .INIT(64'b0000010100000101010001010101010100000100010001000100010001000100)  
) LUT6_25 (
   .O(gates_25),
   .I0(InputBits[218]),
   .I1(InputBits[395]),
   .I2(InputBits[300]),
   .I3(InputBits[447]),
   .I4(InputBits[484]),
   .I5(InputBits[285])
);
LUT6 #(
   .INIT(64'b0000000000000000010101010101010100000001000000000101010101000000)  
) LUT6_26 (
   .O(gates_26),
   .I0(InputBits[530]),
   .I1(InputBits[227]),
   .I2(InputBits[164]),
   .I3(InputBits[396]),
   .I4(InputBits[18]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010001000100000000000000000000010001010101)  
) LUT6_27 (
   .O(gates_27),
   .I0(InputBits[27]),
   .I1(InputBits[548]),
   .I2(InputBits[233]),
   .I3(InputBits[252]),
   .I4(InputBits[3]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000010100000001000000010000001100000011)  
) LUT6_28 (
   .O(gates_28),
   .I0(InputBits[264]),
   .I1(InputBits[535]),
   .I2(InputBits[122]),
   .I3(InputBits[89]),
   .I4(InputBits[70]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b1100111100001100110111110011101111000001011100010000001010110011)  
) LUT6_29 (
   .O(gates_29),
   .I0(InputBits[157]),
   .I1(InputBits[106]),
   .I2(InputBits[64]),
   .I3(InputBits[83]),
   .I4(InputBits[151]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000100010001000110010000101110111)  
) LUT6_30 (
   .O(gates_30),
   .I0(InputBits[287]),
   .I1(InputBits[546]),
   .I2(InputBits[110]),
   .I3(InputBits[484]),
   .I4(InputBits[84]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0000001100100001000000110010001100000011001000000000001100100011)  
) LUT6_31 (
   .O(gates_31),
   .I0(InputBits[327]),
   .I1(InputBits[3]),
   .I2(InputBits[314]),
   .I3(InputBits[311]),
   .I4(InputBits[448]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110001001100000000000000000000000000000011)  
) LUT6_32 (
   .O(gates_32),
   .I0(InputBits[465]),
   .I1(InputBits[533]),
   .I2(InputBits[568]),
   .I3(InputBits[493]),
   .I4(InputBits[169]),
   .I5(InputBits[291])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000010001000100110000011100100011)  
) LUT6_33 (
   .O(gates_33),
   .I0(InputBits[115]),
   .I1(InputBits[29]),
   .I2(InputBits[128]),
   .I3(InputBits[135]),
   .I4(InputBits[550]),
   .I5(InputBits[537])
);
LUT6 #(
   .INIT(64'b0001000000000000000100000000000011011111010011001111111101111111)  
) LUT6_34 (
   .O(gates_34),
   .I0(InputBits[402]),
   .I1(InputBits[432]),
   .I2(InputBits[449]),
   .I3(InputBits[443]),
   .I4(InputBits[105]),
   .I5(InputBits[508])
);
LUT6 #(
   .INIT(64'b0000000000000001000101100011000000010000000101010001010000110101)  
) LUT6_35 (
   .O(gates_35),
   .I0(InputBits[52]),
   .I1(InputBits[94]),
   .I2(InputBits[478]),
   .I3(InputBits[232]),
   .I4(InputBits[411]),
   .I5(InputBits[172])
);
LUT6 #(
   .INIT(64'b0101010101010111010100010101001100010001000000100001000100000010)  
) LUT6_36 (
   .O(gates_36),
   .I0(InputBits[15]),
   .I1(InputBits[124]),
   .I2(InputBits[476]),
   .I3(InputBits[477]),
   .I4(InputBits[58]),
   .I5(InputBits[374])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010001011100000000000100000000000100010010)  
) LUT6_37 (
   .O(gates_37),
   .I0(InputBits[71]),
   .I1(InputBits[362]),
   .I2(InputBits[550]),
   .I3(InputBits[46]),
   .I4(InputBits[147]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0010000100100011000000010010001100100010001001110010011100110011)  
) LUT6_38 (
   .O(gates_38),
   .I0(InputBits[39]),
   .I1(InputBits[504]),
   .I2(InputBits[299]),
   .I3(InputBits[59]),
   .I4(InputBits[111]),
   .I5(InputBits[357])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011110001111101010101010001010000)  
) LUT6_39 (
   .O(gates_39),
   .I0(InputBits[278]),
   .I1(InputBits[379]),
   .I2(InputBits[317]),
   .I3(InputBits[316]),
   .I4(InputBits[346]),
   .I5(InputBits[507])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011000000110001000100010001)  
) LUT6_40 (
   .O(gates_40),
   .I0(InputBits[564]),
   .I1(InputBits[50]),
   .I2(InputBits[110]),
   .I3(InputBits[137]),
   .I4(InputBits[304]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0000001100000001000001110010000000000011000000110000100100000101)  
) LUT6_41 (
   .O(gates_41),
   .I0(InputBits[305]),
   .I1(InputBits[264]),
   .I2(InputBits[551]),
   .I3(InputBits[89]),
   .I4(InputBits[454]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000010001000000010001000100000000000110011)  
) LUT6_42 (
   .O(gates_42),
   .I0(InputBits[418]),
   .I1(InputBits[19]),
   .I2(InputBits[424]),
   .I3(InputBits[563]),
   .I4(InputBits[281]),
   .I5(InputBits[299])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001010101000000000000000000010000011111110)  
) LUT6_43 (
   .O(gates_43),
   .I0(InputBits[394]),
   .I1(InputBits[201]),
   .I2(InputBits[236]),
   .I3(InputBits[147]),
   .I4(InputBits[26]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0001000100110001000100010011001100000000001100110000000000110011)  
) LUT6_44 (
   .O(gates_44),
   .I0(InputBits[128]),
   .I1(InputBits[554]),
   .I2(InputBits[280]),
   .I3(InputBits[277]),
   .I4(InputBits[474]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0000000000010000000000010010000010010101111101011111110111110101)  
) LUT6_45 (
   .O(gates_45),
   .I0(InputBits[135]),
   .I1(InputBits[161]),
   .I2(InputBits[414]),
   .I3(InputBits[283]),
   .I4(InputBits[197]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011000000000000000000000001001100110011)  
) LUT6_46 (
   .O(gates_46),
   .I0(InputBits[519]),
   .I1(InputBits[337]),
   .I2(InputBits[443]),
   .I3(InputBits[264]),
   .I4(InputBits[481]),
   .I5(InputBits[537])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000001000100000001)  
) LUT6_47 (
   .O(gates_47),
   .I0(InputBits[123]),
   .I1(InputBits[473]),
   .I2(InputBits[483]),
   .I3(InputBits[428]),
   .I4(InputBits[505]),
   .I5(InputBits[147])
);
LUT6 #(
   .INIT(64'b0000001100000011000000110001001100001111000001110000001100111111)  
) LUT6_48 (
   .O(gates_48),
   .I0(InputBits[131]),
   .I1(InputBits[386]),
   .I2(InputBits[253]),
   .I3(InputBits[357]),
   .I4(InputBits[425]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000000011111111111011101)  
) LUT6_49 (
   .O(gates_49),
   .I0(InputBits[539]),
   .I1(InputBits[248]),
   .I2(InputBits[161]),
   .I3(InputBits[268]),
   .I4(InputBits[5]),
   .I5(InputBits[20])
);
LUT6 #(
   .INIT(64'b0000000000000011000000010000001100000001000100110000000100001001)  
) LUT6_50 (
   .O(gates_50),
   .I0(InputBits[486]),
   .I1(InputBits[557]),
   .I2(InputBits[566]),
   .I3(InputBits[14]),
   .I4(InputBits[261]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101010001010000010101010101)  
) LUT6_51 (
   .O(gates_51),
   .I0(InputBits[4]),
   .I1(InputBits[201]),
   .I2(InputBits[517]),
   .I3(InputBits[58]),
   .I4(InputBits[104]),
   .I5(InputBits[530])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000000000011000000110000011100000111)  
) LUT6_52 (
   .O(gates_52),
   .I0(InputBits[89]),
   .I1(InputBits[570]),
   .I2(InputBits[506]),
   .I3(InputBits[188]),
   .I4(InputBits[526]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0000011100000101000000000000000100001111000001010000010100000001)  
) LUT6_53 (
   .O(gates_53),
   .I0(InputBits[251]),
   .I1(InputBits[484]),
   .I2(InputBits[27]),
   .I3(InputBits[159]),
   .I4(InputBits[67]),
   .I5(InputBits[304])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010100000000000000000101010101010000)  
) LUT6_54 (
   .O(gates_54),
   .I0(InputBits[558]),
   .I1(InputBits[185]),
   .I2(InputBits[268]),
   .I3(InputBits[392]),
   .I4(InputBits[48]),
   .I5(InputBits[480])
);
LUT6 #(
   .INIT(64'b1111101011111111001100001111100101111010011110111011001110110010)  
) LUT6_55 (
   .O(gates_55),
   .I0(InputBits[285]),
   .I1(InputBits[496]),
   .I2(InputBits[317]),
   .I3(InputBits[181]),
   .I4(InputBits[200]),
   .I5(InputBits[223])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001010000001000000111000000101)  
) LUT6_56 (
   .O(gates_56),
   .I0(InputBits[96]),
   .I1(InputBits[201]),
   .I2(InputBits[2]),
   .I3(InputBits[280]),
   .I4(InputBits[510]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010000000100000001)  
) LUT6_57 (
   .O(gates_57),
   .I0(InputBits[74]),
   .I1(InputBits[553]),
   .I2(InputBits[146]),
   .I3(InputBits[467]),
   .I4(InputBits[327]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0000010100011100000000000100110000000001000000000001000000000101)  
) LUT6_58 (
   .O(gates_58),
   .I0(InputBits[534]),
   .I1(InputBits[178]),
   .I2(InputBits[314]),
   .I3(InputBits[219]),
   .I4(InputBits[401]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0000111100000111000000110000111100000111000011100000011100000100)  
) LUT6_59 (
   .O(gates_59),
   .I0(InputBits[382]),
   .I1(InputBits[267]),
   .I2(InputBits[313]),
   .I3(InputBits[398]),
   .I4(InputBits[197]),
   .I5(InputBits[419])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000111000010111011101100111111)  
) LUT6_60 (
   .O(gates_60),
   .I0(InputBits[89]),
   .I1(InputBits[206]),
   .I2(InputBits[60]),
   .I3(InputBits[522]),
   .I4(InputBits[549]),
   .I5(InputBits[1])
);
LUT6 #(
   .INIT(64'b0000000000000000001110101111011100000000000000010010101011111111)  
) LUT6_61 (
   .O(gates_61),
   .I0(InputBits[316]),
   .I1(InputBits[536]),
   .I2(InputBits[296]),
   .I3(InputBits[109]),
   .I4(InputBits[29]),
   .I5(InputBits[117])
);
LUT6 #(
   .INIT(64'b0000000000000000000010010000100100000000100010010000111100000100)  
) LUT6_62 (
   .O(gates_62),
   .I0(InputBits[469]),
   .I1(InputBits[468]),
   .I2(InputBits[475]),
   .I3(InputBits[248]),
   .I4(InputBits[408]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0011000000000000001100000011000000010011000000000011001100010000)  
) LUT6_63 (
   .O(gates_63),
   .I0(InputBits[58]),
   .I1(InputBits[24]),
   .I2(InputBits[283]),
   .I3(InputBits[394]),
   .I4(InputBits[257]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100000101011110010011001101111)  
) LUT6_64 (
   .O(gates_64),
   .I0(InputBits[41]),
   .I1(InputBits[178]),
   .I2(InputBits[303]),
   .I3(InputBits[483]),
   .I4(InputBits[113]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b0000000100000001000001010000000000000001000000010000000000000000)  
) LUT6_65 (
   .O(gates_65),
   .I0(InputBits[125]),
   .I1(InputBits[508]),
   .I2(InputBits[560]),
   .I3(InputBits[94]),
   .I4(InputBits[295]),
   .I5(InputBits[323])
);
LUT6 #(
   .INIT(64'b0000000001101111000000000111111100000000111111000000000001010000)  
) LUT6_66 (
   .O(gates_66),
   .I0(InputBits[138]),
   .I1(InputBits[547]),
   .I2(InputBits[267]),
   .I3(InputBits[457]),
   .I4(InputBits[161]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000000000000000000011000100110000000000000000000000000011111100)  
) LUT6_67 (
   .O(gates_67),
   .I0(InputBits[115]),
   .I1(InputBits[345]),
   .I2(InputBits[296]),
   .I3(InputBits[278]),
   .I4(InputBits[385]),
   .I5(InputBits[57])
);
LUT6 #(
   .INIT(64'b0000000000001111000000010000100100101111001110110001011100000000)  
) LUT6_68 (
   .O(gates_68),
   .I0(InputBits[249]),
   .I1(InputBits[157]),
   .I2(InputBits[569]),
   .I3(InputBits[268]),
   .I4(InputBits[200]),
   .I5(InputBits[67])
);
LUT6 #(
   .INIT(64'b0101000001010101000100010101000101000100010101010100010001010000)  
) LUT6_69 (
   .O(gates_69),
   .I0(InputBits[97]),
   .I1(InputBits[446]),
   .I2(InputBits[370]),
   .I3(InputBits[544]),
   .I4(InputBits[178]),
   .I5(InputBits[92])
);
LUT6 #(
   .INIT(64'b0011011101010101011101110010000001010011010101010011001100010111)  
) LUT6_70 (
   .O(gates_70),
   .I0(InputBits[549]),
   .I1(InputBits[66]),
   .I2(InputBits[281]),
   .I3(InputBits[524]),
   .I4(InputBits[367]),
   .I5(InputBits[105])
);
LUT6 #(
   .INIT(64'b0000000000000000000100100000010000000010000000110011001101110011)  
) LUT6_71 (
   .O(gates_71),
   .I0(InputBits[430]),
   .I1(InputBits[565]),
   .I2(InputBits[363]),
   .I3(InputBits[152]),
   .I4(InputBits[12]),
   .I5(InputBits[493])
);
LUT6 #(
   .INIT(64'b0000000000000100000001000000110000000100000011010000010101000101)  
) LUT6_72 (
   .O(gates_72),
   .I0(InputBits[508]),
   .I1(InputBits[199]),
   .I2(InputBits[21]),
   .I3(InputBits[210]),
   .I4(InputBits[460]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001000100010001011111111111111111)  
) LUT6_73 (
   .O(gates_73),
   .I0(InputBits[305]),
   .I1(InputBits[392]),
   .I2(InputBits[429]),
   .I3(InputBits[464]),
   .I4(InputBits[253]),
   .I5(InputBits[529])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010000000000010001000000110011001100000011)  
) LUT6_74 (
   .O(gates_74),
   .I0(InputBits[519]),
   .I1(InputBits[265]),
   .I2(InputBits[106]),
   .I3(InputBits[415]),
   .I4(InputBits[304]),
   .I5(InputBits[534])
);
LUT6 #(
   .INIT(64'b0011000100010001000100100000001100010000000100010000000000000001)  
) LUT6_75 (
   .O(gates_75),
   .I0(InputBits[30]),
   .I1(InputBits[313]),
   .I2(InputBits[380]),
   .I3(InputBits[378]),
   .I4(InputBits[359]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0000001100000010000000110000001100100011000100100000001100110011)  
) LUT6_76 (
   .O(gates_76),
   .I0(InputBits[323]),
   .I1(InputBits[554]),
   .I2(InputBits[480]),
   .I3(InputBits[178]),
   .I4(InputBits[304]),
   .I5(InputBits[339])
);
LUT6 #(
   .INIT(64'b0000001100000000001100110001000000000011000000000011001100110001)  
) LUT6_77 (
   .O(gates_77),
   .I0(InputBits[56]),
   .I1(InputBits[385]),
   .I2(InputBits[325]),
   .I3(InputBits[236]),
   .I4(InputBits[515]),
   .I5(InputBits[329])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000100101000101010001111111111111011)  
) LUT6_78 (
   .O(gates_78),
   .I0(InputBits[269]),
   .I1(InputBits[197]),
   .I2(InputBits[282]),
   .I3(InputBits[437]),
   .I4(InputBits[278]),
   .I5(InputBits[6])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101000001010000010101010111)  
) LUT6_79 (
   .O(gates_79),
   .I0(InputBits[277]),
   .I1(InputBits[299]),
   .I2(InputBits[558]),
   .I3(InputBits[356]),
   .I4(InputBits[60]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000011000000000000000000000010001011111)  
) LUT6_80 (
   .O(gates_80),
   .I0(InputBits[240]),
   .I1(InputBits[261]),
   .I2(InputBits[548]),
   .I3(InputBits[509]),
   .I4(InputBits[169]),
   .I5(InputBits[540])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000111110000000000011111010)  
) LUT6_81 (
   .O(gates_81),
   .I0(InputBits[309]),
   .I1(InputBits[414]),
   .I2(InputBits[395]),
   .I3(InputBits[531]),
   .I4(InputBits[357]),
   .I5(InputBits[573])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010010001000000000000000000001000100100011)  
) LUT6_82 (
   .O(gates_82),
   .I0(InputBits[268]),
   .I1(InputBits[434]),
   .I2(InputBits[327]),
   .I3(InputBits[384]),
   .I4(InputBits[559]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000000000000000010000000110000000000001010011100110011001111)  
) LUT6_83 (
   .O(gates_83),
   .I0(InputBits[464]),
   .I1(InputBits[394]),
   .I2(InputBits[460]),
   .I3(InputBits[494]),
   .I4(InputBits[52]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000100000011)  
) LUT6_84 (
   .O(gates_84),
   .I0(InputBits[21]),
   .I1(InputBits[338]),
   .I2(InputBits[50]),
   .I3(InputBits[428]),
   .I4(InputBits[108]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0000000000000000000011001101110100000001010011101100110111001101)  
) LUT6_85 (
   .O(gates_85),
   .I0(InputBits[300]),
   .I1(InputBits[372]),
   .I2(InputBits[231]),
   .I3(InputBits[356]),
   .I4(InputBits[120]),
   .I5(InputBits[500])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000100000000000000010000000000000001)  
) LUT6_86 (
   .O(gates_86),
   .I0(InputBits[506]),
   .I1(InputBits[276]),
   .I2(InputBits[76]),
   .I3(InputBits[553]),
   .I4(InputBits[567]),
   .I5(InputBits[468])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000111100100000010011110000)  
) LUT6_87 (
   .O(gates_87),
   .I0(InputBits[412]),
   .I1(InputBits[282]),
   .I2(InputBits[370]),
   .I3(InputBits[290]),
   .I4(InputBits[404]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b0000000010000000100011111111111100000000010100101010111111101010)  
) LUT6_88 (
   .O(gates_88),
   .I0(InputBits[364]),
   .I1(InputBits[176]),
   .I2(InputBits[329]),
   .I3(InputBits[467]),
   .I4(InputBits[569]),
   .I5(InputBits[441])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000001000100000000000000010000000000010001)  
) LUT6_89 (
   .O(gates_89),
   .I0(InputBits[74]),
   .I1(InputBits[494]),
   .I2(InputBits[43]),
   .I3(InputBits[50]),
   .I4(InputBits[174]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0000000100000010000000110000001100001111000011100000111100001110)  
) LUT6_90 (
   .O(gates_90),
   .I0(InputBits[396]),
   .I1(InputBits[244]),
   .I2(InputBits[122]),
   .I3(InputBits[200]),
   .I4(InputBits[469]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b1000111100000110001101110100001010101111101111111110011111111010)  
) LUT6_91 (
   .O(gates_91),
   .I0(InputBits[350]),
   .I1(InputBits[118]),
   .I2(InputBits[325]),
   .I3(InputBits[213]),
   .I4(InputBits[212]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000001000111101111111111110000100010101011)  
) LUT6_92 (
   .O(gates_92),
   .I0(InputBits[166]),
   .I1(InputBits[380]),
   .I2(InputBits[435]),
   .I3(InputBits[513]),
   .I4(InputBits[295]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000001001100000000000000010000000100010001)  
) LUT6_93 (
   .O(gates_93),
   .I0(InputBits[275]),
   .I1(InputBits[409]),
   .I2(InputBits[230]),
   .I3(InputBits[459]),
   .I4(InputBits[543]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0000010000000100000001000000010000001111000011100000111100001111)  
) LUT6_94 (
   .O(gates_94),
   .I0(InputBits[502]),
   .I1(InputBits[318]),
   .I2(InputBits[169]),
   .I3(InputBits[399]),
   .I4(InputBits[473]),
   .I5(InputBits[539])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001011000010111010111110111111001110110010)  
) LUT6_95 (
   .O(gates_95),
   .I0(InputBits[369]),
   .I1(InputBits[125]),
   .I2(InputBits[395]),
   .I3(InputBits[479]),
   .I4(InputBits[431]),
   .I5(InputBits[435])
);
LUT6 #(
   .INIT(64'b1111101011111010111111101111111101011100011101111101101011111010)  
) LUT6_96 (
   .O(gates_96),
   .I0(InputBits[393]),
   .I1(InputBits[87]),
   .I2(InputBits[342]),
   .I3(InputBits[500]),
   .I4(InputBits[245]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000000000110010000000000111110000000000001100010000000001111101)  
) LUT6_97 (
   .O(gates_97),
   .I0(InputBits[474]),
   .I1(InputBits[479]),
   .I2(InputBits[247]),
   .I3(InputBits[47]),
   .I4(InputBits[141]),
   .I5(InputBits[86])
);
LUT6 #(
   .INIT(64'b0000011000001000000011110000111110001110100000101100111111101011)  
) LUT6_98 (
   .O(gates_98),
   .I0(InputBits[374]),
   .I1(InputBits[57]),
   .I2(InputBits[31]),
   .I3(InputBits[454]),
   .I4(InputBits[228]),
   .I5(InputBits[153])
);
LUT6 #(
   .INIT(64'b1111111111111111010011101111111100111110111111100000110011001100)  
) LUT6_99 (
   .O(gates_99),
   .I0(InputBits[187]),
   .I1(InputBits[200]),
   .I2(InputBits[324]),
   .I3(InputBits[488]),
   .I4(InputBits[416]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0010001000100000001000100010001000110011001000110011001100100011)  
) LUT6_100 (
   .O(gates_100),
   .I0(InputBits[238]),
   .I1(InputBits[362]),
   .I2(InputBits[492]),
   .I3(InputBits[249]),
   .I4(InputBits[215]),
   .I5(InputBits[105])
);
LUT6 #(
   .INIT(64'b1111000011110000000001010000010011110000111000000000000000000000)  
) LUT6_101 (
   .O(gates_101),
   .I0(InputBits[198]),
   .I1(InputBits[117]),
   .I2(InputBits[270]),
   .I3(InputBits[326]),
   .I4(InputBits[270]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0101010100000000000000000000000001010101010101000101010101110100)  
) LUT6_102 (
   .O(gates_102),
   .I0(InputBits[7]),
   .I1(InputBits[358]),
   .I2(InputBits[445]),
   .I3(InputBits[247]),
   .I4(InputBits[153]),
   .I5(InputBits[255])
);
LUT6 #(
   .INIT(64'b0000010000000100000000000000010000000101001011100101010111101110)  
) LUT6_103 (
   .O(gates_103),
   .I0(InputBits[383]),
   .I1(InputBits[341]),
   .I2(InputBits[232]),
   .I3(InputBits[68]),
   .I4(InputBits[461]),
   .I5(InputBits[386])
);
LUT6 #(
   .INIT(64'b0000000000010100000000000101010101010101010100110101000111010001)  
) LUT6_104 (
   .O(gates_104),
   .I0(InputBits[564]),
   .I1(InputBits[279]),
   .I2(InputBits[373]),
   .I3(InputBits[545]),
   .I4(InputBits[221]),
   .I5(InputBits[408])
);
LUT6 #(
   .INIT(64'b0000000000010111000000000101000100000000000111110000000001011111)  
) LUT6_105 (
   .O(gates_105),
   .I0(InputBits[167]),
   .I1(InputBits[516]),
   .I2(InputBits[455]),
   .I3(InputBits[169]),
   .I4(InputBits[309]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0011001100100010101101110010001100110011001100000011001100001000)  
) LUT6_106 (
   .O(gates_106),
   .I0(InputBits[423]),
   .I1(InputBits[147]),
   .I2(InputBits[413]),
   .I3(InputBits[344]),
   .I4(InputBits[157]),
   .I5(InputBits[477])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000010100000000000000000000001100000010)  
) LUT6_107 (
   .O(gates_107),
   .I0(InputBits[7]),
   .I1(InputBits[531]),
   .I2(InputBits[121]),
   .I3(InputBits[384]),
   .I4(InputBits[434]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1111111101011111111111110001111101010101000001010101011100000101)  
) LUT6_108 (
   .O(gates_108),
   .I0(InputBits[274]),
   .I1(InputBits[156]),
   .I2(InputBits[106]),
   .I3(InputBits[441]),
   .I4(InputBits[466]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010001000000001000101000001111)  
) LUT6_109 (
   .O(gates_109),
   .I0(InputBits[358]),
   .I1(InputBits[156]),
   .I2(InputBits[172]),
   .I3(InputBits[353]),
   .I4(InputBits[219]),
   .I5(InputBits[563])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001000000000000000110000001100100011)  
) LUT6_110 (
   .O(gates_110),
   .I0(InputBits[446]),
   .I1(InputBits[146]),
   .I2(InputBits[6]),
   .I3(InputBits[46]),
   .I4(InputBits[547]),
   .I5(InputBits[54])
);
LUT6 #(
   .INIT(64'b0000010100010101111111111111110100000101000001011111110011111111)  
) LUT6_111 (
   .O(gates_111),
   .I0(InputBits[523]),
   .I1(InputBits[346]),
   .I2(InputBits[200]),
   .I3(InputBits[402]),
   .I4(InputBits[13]),
   .I5(InputBits[341])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000000010100000001010111110000000000001011)  
) LUT6_112 (
   .O(gates_112),
   .I0(InputBits[10]),
   .I1(InputBits[83]),
   .I2(InputBits[485]),
   .I3(InputBits[20]),
   .I4(InputBits[366]),
   .I5(InputBits[14])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000100100000000000100000001001100011111)  
) LUT6_113 (
   .O(gates_113),
   .I0(InputBits[71]),
   .I1(InputBits[513]),
   .I2(InputBits[494]),
   .I3(InputBits[469]),
   .I4(InputBits[568]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000100000000000100110001000100000011)  
) LUT6_114 (
   .O(gates_114),
   .I0(InputBits[517]),
   .I1(InputBits[25]),
   .I2(InputBits[275]),
   .I3(InputBits[36]),
   .I4(InputBits[204]),
   .I5(InputBits[562])
);
LUT6 #(
   .INIT(64'b0000000011001000000000000100010010000000111111000000010011111100)  
) LUT6_115 (
   .O(gates_115),
   .I0(InputBits[203]),
   .I1(InputBits[392]),
   .I2(InputBits[397]),
   .I3(InputBits[531]),
   .I4(InputBits[158]),
   .I5(InputBits[482])
);
LUT6 #(
   .INIT(64'b0000100000000000000000100010000000100000001000000011000000110000)  
) LUT6_116 (
   .O(gates_116),
   .I0(InputBits[442]),
   .I1(InputBits[507]),
   .I2(InputBits[347]),
   .I3(InputBits[429]),
   .I4(InputBits[134]),
   .I5(InputBits[508])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000101010000001100101111)  
) LUT6_117 (
   .O(gates_117),
   .I0(InputBits[114]),
   .I1(InputBits[402]),
   .I2(InputBits[82]),
   .I3(InputBits[567]),
   .I4(InputBits[527]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0000000001000000000000000000000000000000000100000000000001110011)  
) LUT6_118 (
   .O(gates_118),
   .I0(InputBits[185]),
   .I1(InputBits[448]),
   .I2(InputBits[93]),
   .I3(InputBits[571]),
   .I4(InputBits[108]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000001000000000000001010000)  
) LUT6_119 (
   .O(gates_119),
   .I0(InputBits[266]),
   .I1(InputBits[192]),
   .I2(InputBits[325]),
   .I3(InputBits[127]),
   .I4(InputBits[497]),
   .I5(InputBits[561])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001000100000000000000000000000000000000)  
) LUT6_120 (
   .O(gates_120),
   .I0(InputBits[457]),
   .I1(InputBits[193]),
   .I2(InputBits[290]),
   .I3(InputBits[552]),
   .I4(InputBits[60]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b0000000001000101000000000000011100010101010001100101010101010111)  
) LUT6_121 (
   .O(gates_121),
   .I0(InputBits[527]),
   .I1(InputBits[367]),
   .I2(InputBits[203]),
   .I3(InputBits[408]),
   .I4(InputBits[108]),
   .I5(InputBits[524])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000100010100000000000000001101000110100111)  
) LUT6_122 (
   .O(gates_122),
   .I0(InputBits[12]),
   .I1(InputBits[133]),
   .I2(InputBits[448]),
   .I3(InputBits[476]),
   .I4(InputBits[123]),
   .I5(InputBits[45])
);
LUT6 #(
   .INIT(64'b0000000000000000001111111111111100000000000000001111101100100010)  
) LUT6_123 (
   .O(gates_123),
   .I0(InputBits[443]),
   .I1(InputBits[127]),
   .I2(InputBits[90]),
   .I3(InputBits[345]),
   .I4(InputBits[289]),
   .I5(InputBits[190])
);
LUT6 #(
   .INIT(64'b0011101110110011001000000011001010111011101111110010001010111011)  
) LUT6_124 (
   .O(gates_124),
   .I0(InputBits[270]),
   .I1(InputBits[255]),
   .I2(InputBits[114]),
   .I3(InputBits[473]),
   .I4(InputBits[341]),
   .I5(InputBits[436])
);
LUT6 #(
   .INIT(64'b0010000010110010001100011111011100100000011000110111000101110111)  
) LUT6_125 (
   .O(gates_125),
   .I0(InputBits[486]),
   .I1(InputBits[276]),
   .I2(InputBits[270]),
   .I3(InputBits[518]),
   .I4(InputBits[510]),
   .I5(InputBits[159])
);
LUT6 #(
   .INIT(64'b1111110111110001010011110111111111111111111111011111111111111100)  
) LUT6_126 (
   .O(gates_126),
   .I0(InputBits[429]),
   .I1(InputBits[398]),
   .I2(InputBits[392]),
   .I3(InputBits[395]),
   .I4(InputBits[393]),
   .I5(InputBits[213])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001000100000000001000110000000000110011)  
) LUT6_127 (
   .O(gates_127),
   .I0(InputBits[300]),
   .I1(InputBits[555]),
   .I2(InputBits[249]),
   .I3(InputBits[27]),
   .I4(InputBits[549]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0000000000000000000010101010111000001000000011101001111100101100)  
) LUT6_128 (
   .O(gates_128),
   .I0(InputBits[399]),
   .I1(InputBits[348]),
   .I2(InputBits[46]),
   .I3(InputBits[270]),
   .I4(InputBits[32]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0011000000110001011100000101000000110011001100110111001111110100)  
) LUT6_129 (
   .O(gates_129),
   .I0(InputBits[208]),
   .I1(InputBits[167]),
   .I2(InputBits[319]),
   .I3(InputBits[370]),
   .I4(InputBits[334]),
   .I5(InputBits[493])
);
LUT6 #(
   .INIT(64'b0000000000000001000111110000010100000000000001010001111100000001)  
) LUT6_130 (
   .O(gates_130),
   .I0(InputBits[81]),
   .I1(InputBits[462]),
   .I2(InputBits[242]),
   .I3(InputBits[292]),
   .I4(InputBits[192]),
   .I5(InputBits[90])
);
LUT6 #(
   .INIT(64'b0000000000000000010000010100010111111011110111110011001101011011)  
) LUT6_131 (
   .O(gates_131),
   .I0(InputBits[69]),
   .I1(InputBits[207]),
   .I2(InputBits[182]),
   .I3(InputBits[273]),
   .I4(InputBits[68]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0000010011001100110011111100110010100000110011111110011111101111)  
) LUT6_132 (
   .O(gates_132),
   .I0(InputBits[164]),
   .I1(InputBits[365]),
   .I2(InputBits[427]),
   .I3(InputBits[523]),
   .I4(InputBits[249]),
   .I5(InputBits[110])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000000000010110011001100001111011100110000)  
) LUT6_133 (
   .O(gates_133),
   .I0(InputBits[160]),
   .I1(InputBits[300]),
   .I2(InputBits[351]),
   .I3(InputBits[222]),
   .I4(InputBits[88]),
   .I5(InputBits[482])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001111111100000000000000000000000000011101)  
) LUT6_134 (
   .O(gates_134),
   .I0(InputBits[81]),
   .I1(InputBits[244]),
   .I2(InputBits[156]),
   .I3(InputBits[433]),
   .I4(InputBits[575]),
   .I5(InputBits[316])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001101000011010000110000001101)  
) LUT6_135 (
   .O(gates_135),
   .I0(InputBits[494]),
   .I1(InputBits[367]),
   .I2(InputBits[241]),
   .I3(InputBits[512]),
   .I4(InputBits[429]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0000000001011101000000000000000000000000001111110000000000000010)  
) LUT6_136 (
   .O(gates_136),
   .I0(InputBits[119]),
   .I1(InputBits[209]),
   .I2(InputBits[133]),
   .I3(InputBits[192]),
   .I4(InputBits[373]),
   .I5(InputBits[357])
);
LUT6 #(
   .INIT(64'b0000000000000000100010111000111000000000000000001010101010101010)  
) LUT6_137 (
   .O(gates_137),
   .I0(InputBits[397]),
   .I1(InputBits[452]),
   .I2(InputBits[491]),
   .I3(InputBits[177]),
   .I4(InputBits[21]),
   .I5(InputBits[447])
);
LUT6 #(
   .INIT(64'b0011111100001111000000000000110010101111000011011100110001001100)  
) LUT6_138 (
   .O(gates_138),
   .I0(InputBits[113]),
   .I1(InputBits[368]),
   .I2(InputBits[508]),
   .I3(InputBits[413]),
   .I4(InputBits[342]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0000000011111111000000001111111100000000110011110000000001001111)  
) LUT6_139 (
   .O(gates_139),
   .I0(InputBits[157]),
   .I1(InputBits[258]),
   .I2(InputBits[402]),
   .I3(InputBits[481]),
   .I4(InputBits[466]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0111111101101011011100111011001001011111111111111111101111111111)  
) LUT6_140 (
   .O(gates_140),
   .I0(InputBits[375]),
   .I1(InputBits[205]),
   .I2(InputBits[430]),
   .I3(InputBits[174]),
   .I4(InputBits[310]),
   .I5(InputBits[103])
);
LUT6 #(
   .INIT(64'b0000000011001111000000001100111000000000111110111100000011111111)  
) LUT6_141 (
   .O(gates_141),
   .I0(InputBits[283]),
   .I1(InputBits[524]),
   .I2(InputBits[257]),
   .I3(InputBits[242]),
   .I4(InputBits[364]),
   .I5(InputBits[105])
);
LUT6 #(
   .INIT(64'b0000110000001100000011110000110100001000000010000000111111111111)  
) LUT6_142 (
   .O(gates_142),
   .I0(InputBits[151]),
   .I1(InputBits[268]),
   .I2(InputBits[566]),
   .I3(InputBits[64]),
   .I4(InputBits[515]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1011101000000010011100000000001011111111011110101111111011111110)  
) LUT6_143 (
   .O(gates_143),
   .I0(InputBits[335]),
   .I1(InputBits[239]),
   .I2(InputBits[343]),
   .I3(InputBits[247]),
   .I4(InputBits[186]),
   .I5(InputBits[519])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000010111111100100101011111110)  
) LUT6_144 (
   .O(gates_144),
   .I0(InputBits[421]),
   .I1(InputBits[319]),
   .I2(InputBits[285]),
   .I3(InputBits[77]),
   .I4(InputBits[64]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0001001100100010000000100000001000010011001100100010001100100010)  
) LUT6_145 (
   .O(gates_145),
   .I0(InputBits[420]),
   .I1(InputBits[555]),
   .I2(InputBits[65]),
   .I3(InputBits[359]),
   .I4(InputBits[451]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0000000101000000010101010101000000000000000000000001000000010000)  
) LUT6_146 (
   .O(gates_146),
   .I0(InputBits[241]),
   .I1(InputBits[520]),
   .I2(InputBits[418]),
   .I3(InputBits[415]),
   .I4(InputBits[76]),
   .I5(InputBits[211])
);
LUT6 #(
   .INIT(64'b0000110100001100000011010000010000001111000011100000111100001111)  
) LUT6_147 (
   .O(gates_147),
   .I0(InputBits[405]),
   .I1(InputBits[391]),
   .I2(InputBits[553]),
   .I3(InputBits[358]),
   .I4(InputBits[490]),
   .I5(InputBits[495])
);
LUT6 #(
   .INIT(64'b0000000000010001000001000001001101010101001000110101010101110111)  
) LUT6_148 (
   .O(gates_148),
   .I0(InputBits[11]),
   .I1(InputBits[515]),
   .I2(InputBits[462]),
   .I3(InputBits[262]),
   .I4(InputBits[278]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0100000001010101111101111110111100000000000101001111011101100111)  
) LUT6_149 (
   .O(gates_149),
   .I0(InputBits[286]),
   .I1(InputBits[38]),
   .I2(InputBits[426]),
   .I3(InputBits[211]),
   .I4(InputBits[11]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b1111111011111111001100110101010110111111111111111011001101110101)  
) LUT6_150 (
   .O(gates_150),
   .I0(InputBits[354]),
   .I1(InputBits[493]),
   .I2(InputBits[116]),
   .I3(InputBits[376]),
   .I4(InputBits[261]),
   .I5(InputBits[64])
);
LUT6 #(
   .INIT(64'b0000010100000101000001000000010111010111010001100101111101011110)  
) LUT6_151 (
   .O(gates_151),
   .I0(InputBits[360]),
   .I1(InputBits[200]),
   .I2(InputBits[454]),
   .I3(InputBits[397]),
   .I4(InputBits[297]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b0101010101000100010101010100010100010101000000000101010101000111)  
) LUT6_152 (
   .O(gates_152),
   .I0(InputBits[574]),
   .I1(InputBits[320]),
   .I2(InputBits[520]),
   .I3(InputBits[317]),
   .I4(InputBits[490]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0000101000110011001100110010101111001111000100111111101100000111)  
) LUT6_153 (
   .O(gates_153),
   .I0(InputBits[306]),
   .I1(InputBits[491]),
   .I2(InputBits[520]),
   .I3(InputBits[291]),
   .I4(InputBits[469]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0001111100011111000111110001101100001100000001000000010000011110)  
) LUT6_154 (
   .O(gates_154),
   .I0(InputBits[476]),
   .I1(InputBits[244]),
   .I2(InputBits[13]),
   .I3(InputBits[328]),
   .I4(InputBits[307]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0001010001000101000000000000000000010101010101010100010000000100)  
) LUT6_155 (
   .O(gates_155),
   .I0(InputBits[97]),
   .I1(InputBits[220]),
   .I2(InputBits[183]),
   .I3(InputBits[448]),
   .I4(InputBits[395]),
   .I5(InputBits[172])
);
LUT6 #(
   .INIT(64'b0100010001010101010001000101010100000100010101010000010101010101)  
) LUT6_156 (
   .O(gates_156),
   .I0(InputBits[557]),
   .I1(InputBits[406]),
   .I2(InputBits[461]),
   .I3(InputBits[230]),
   .I4(InputBits[56]),
   .I5(InputBits[59])
);
LUT6 #(
   .INIT(64'b0000000000000000000011110000111100000000000000000000011100000000)  
) LUT6_157 (
   .O(gates_157),
   .I0(InputBits[182]),
   .I1(InputBits[209]),
   .I2(InputBits[146]),
   .I3(InputBits[398]),
   .I4(InputBits[122]),
   .I5(InputBits[286])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001011111011111110111011101111111011)  
) LUT6_158 (
   .O(gates_158),
   .I0(InputBits[268]),
   .I1(InputBits[495]),
   .I2(InputBits[415]),
   .I3(InputBits[226]),
   .I4(InputBits[157]),
   .I5(InputBits[573])
);
LUT6 #(
   .INIT(64'b0010000100000000001100100001000000000011001101110011001000110011)  
) LUT6_159 (
   .O(gates_159),
   .I0(InputBits[175]),
   .I1(InputBits[251]),
   .I2(InputBits[57]),
   .I3(InputBits[102]),
   .I4(InputBits[92]),
   .I5(InputBits[77])
);
LUT6 #(
   .INIT(64'b0010000000010000001100110001001110101011101000110010001100011100)  
) LUT6_160 (
   .O(gates_160),
   .I0(InputBits[89]),
   .I1(InputBits[544]),
   .I2(InputBits[468]),
   .I3(InputBits[440]),
   .I4(InputBits[522]),
   .I5(InputBits[479])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000000001000000010000000000000000)  
) LUT6_161 (
   .O(gates_161),
   .I0(InputBits[1]),
   .I1(InputBits[555]),
   .I2(InputBits[433]),
   .I3(InputBits[487]),
   .I4(InputBits[394]),
   .I5(InputBits[527])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000000000000001101110000000000111110)  
) LUT6_162 (
   .O(gates_162),
   .I0(InputBits[224]),
   .I1(InputBits[43]),
   .I2(InputBits[268]),
   .I3(InputBits[507]),
   .I4(InputBits[37]),
   .I5(InputBits[362])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000101010100110010111100110100000011111010)  
) LUT6_163 (
   .O(gates_163),
   .I0(InputBits[295]),
   .I1(InputBits[59]),
   .I2(InputBits[347]),
   .I3(InputBits[518]),
   .I4(InputBits[271]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000100000101000000010101111100010111)  
) LUT6_164 (
   .O(gates_164),
   .I0(InputBits[353]),
   .I1(InputBits[539]),
   .I2(InputBits[513]),
   .I3(InputBits[114]),
   .I4(InputBits[531]),
   .I5(InputBits[534])
);
LUT6 #(
   .INIT(64'b0000000000001001000000000000111100000000000000100000000000001010)  
) LUT6_165 (
   .O(gates_165),
   .I0(InputBits[201]),
   .I1(InputBits[135]),
   .I2(InputBits[100]),
   .I3(InputBits[51]),
   .I4(InputBits[257]),
   .I5(InputBits[38])
);
LUT6 #(
   .INIT(64'b0000010000100101101001011010010100000101000000000000000100000101)  
) LUT6_166 (
   .O(gates_166),
   .I0(InputBits[472]),
   .I1(InputBits[158]),
   .I2(InputBits[472]),
   .I3(InputBits[257]),
   .I4(InputBits[57]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001000001001100010011)  
) LUT6_167 (
   .O(gates_167),
   .I0(InputBits[168]),
   .I1(InputBits[574]),
   .I2(InputBits[185]),
   .I3(InputBits[188]),
   .I4(InputBits[255]),
   .I5(InputBits[27])
);
LUT6 #(
   .INIT(64'b0101010100010000000100010001000001010101000100000101000000010001)  
) LUT6_168 (
   .O(gates_168),
   .I0(InputBits[98]),
   .I1(InputBits[171]),
   .I2(InputBits[368]),
   .I3(InputBits[501]),
   .I4(InputBits[162]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000100010100000000111101110000000011110011)  
) LUT6_169 (
   .O(gates_169),
   .I0(InputBits[203]),
   .I1(InputBits[108]),
   .I2(InputBits[178]),
   .I3(InputBits[49]),
   .I4(InputBits[312]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000001000110111011101110111100111111011111)  
) LUT6_170 (
   .O(gates_170),
   .I0(InputBits[60]),
   .I1(InputBits[38]),
   .I2(InputBits[472]),
   .I3(InputBits[301]),
   .I4(InputBits[431]),
   .I5(InputBits[266])
);
LUT6 #(
   .INIT(64'b0000001100000000000011110000010000001111000001010000111100000100)  
) LUT6_171 (
   .O(gates_171),
   .I0(InputBits[300]),
   .I1(InputBits[143]),
   .I2(InputBits[193]),
   .I3(InputBits[397]),
   .I4(InputBits[309]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1000110000100000111111011111111100010000110100010111110111111111)  
) LUT6_172 (
   .O(gates_172),
   .I0(InputBits[150]),
   .I1(InputBits[523]),
   .I2(InputBits[442]),
   .I3(InputBits[299]),
   .I4(InputBits[253]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b0000000000001000000010100000000000001111000011000000101000001010)  
) LUT6_173 (
   .O(gates_173),
   .I0(InputBits[294]),
   .I1(InputBits[212]),
   .I2(InputBits[338]),
   .I3(InputBits[387]),
   .I4(InputBits[452]),
   .I5(InputBits[231])
);
LUT6 #(
   .INIT(64'b0000000010111111000000001010111010000000101110110000000011101111)  
) LUT6_174 (
   .O(gates_174),
   .I0(InputBits[200]),
   .I1(InputBits[199]),
   .I2(InputBits[160]),
   .I3(InputBits[507]),
   .I4(InputBits[180]),
   .I5(InputBits[462])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000101010100000000000000000101010100010101)  
) LUT6_175 (
   .O(gates_175),
   .I0(InputBits[507]),
   .I1(InputBits[183]),
   .I2(InputBits[355]),
   .I3(InputBits[287]),
   .I4(InputBits[507]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b0000000000000101000000001000101000000000001101010000010100110110)  
) LUT6_176 (
   .O(gates_176),
   .I0(InputBits[383]),
   .I1(InputBits[282]),
   .I2(InputBits[406]),
   .I3(InputBits[9]),
   .I4(InputBits[190]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0000001100010011000000110100010100000001001100110000000101000101)  
) LUT6_177 (
   .O(gates_177),
   .I0(InputBits[485]),
   .I1(InputBits[288]),
   .I2(InputBits[540]),
   .I3(InputBits[548]),
   .I4(InputBits[259]),
   .I5(InputBits[303])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000010000001001001111101110)  
) LUT6_178 (
   .O(gates_178),
   .I0(InputBits[223]),
   .I1(InputBits[398]),
   .I2(InputBits[464]),
   .I3(InputBits[527]),
   .I4(InputBits[51]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0000000000000000010101110101010100000000000100011111000001011000)  
) LUT6_179 (
   .O(gates_179),
   .I0(InputBits[43]),
   .I1(InputBits[211]),
   .I2(InputBits[369]),
   .I3(InputBits[92]),
   .I4(InputBits[384]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0000100000001000000010100000100000001000110010001100110011001110)  
) LUT6_180 (
   .O(gates_180),
   .I0(InputBits[296]),
   .I1(InputBits[370]),
   .I2(InputBits[62]),
   .I3(InputBits[160]),
   .I4(InputBits[519]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0010001000110111000000000000010000100010001101110000000000010101)  
) LUT6_181 (
   .O(gates_181),
   .I0(InputBits[436]),
   .I1(InputBits[550]),
   .I2(InputBits[464]),
   .I3(InputBits[483]),
   .I4(InputBits[294]),
   .I5(InputBits[450])
);
LUT6 #(
   .INIT(64'b0000000001011101000000000101010000000001010101000000000101010000)  
) LUT6_182 (
   .O(gates_182),
   .I0(InputBits[564]),
   .I1(InputBits[165]),
   .I2(InputBits[245]),
   .I3(InputBits[10]),
   .I4(InputBits[320]),
   .I5(InputBits[283])
);
LUT6 #(
   .INIT(64'b0000000001010001000000000101000000000000110101010000000001011101)  
) LUT6_183 (
   .O(gates_183),
   .I0(InputBits[314]),
   .I1(InputBits[185]),
   .I2(InputBits[200]),
   .I3(InputBits[560]),
   .I4(InputBits[91]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0000000000000100011111111111111100000000000101001101111111001101)  
) LUT6_184 (
   .O(gates_184),
   .I0(InputBits[81]),
   .I1(InputBits[199]),
   .I2(InputBits[303]),
   .I3(InputBits[261]),
   .I4(InputBits[264]),
   .I5(InputBits[311])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010101000000001101111110101111)  
) LUT6_185 (
   .O(gates_185),
   .I0(InputBits[525]),
   .I1(InputBits[160]),
   .I2(InputBits[541]),
   .I3(InputBits[445]),
   .I4(InputBits[563]),
   .I5(InputBits[557])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000011100000000000010100000010100001011)  
) LUT6_186 (
   .O(gates_186),
   .I0(InputBits[340]),
   .I1(InputBits[495]),
   .I2(InputBits[575]),
   .I3(InputBits[432]),
   .I4(InputBits[434]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010010001100110111011101011101)  
) LUT6_187 (
   .O(gates_187),
   .I0(InputBits[229]),
   .I1(InputBits[116]),
   .I2(InputBits[132]),
   .I3(InputBits[383]),
   .I4(InputBits[479]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0000000000000111000000000100110011101100110111011100110011001100)  
) LUT6_188 (
   .O(gates_188),
   .I0(InputBits[158]),
   .I1(InputBits[341]),
   .I2(InputBits[165]),
   .I3(InputBits[85]),
   .I4(InputBits[296]),
   .I5(InputBits[243])
);
LUT6 #(
   .INIT(64'b0000010001001111000100101111110000000000010011110000000011110011)  
) LUT6_189 (
   .O(gates_189),
   .I0(InputBits[160]),
   .I1(InputBits[402]),
   .I2(InputBits[35]),
   .I3(InputBits[434]),
   .I4(InputBits[141]),
   .I5(InputBits[380])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000100011100000000010101000000000001010010)  
) LUT6_190 (
   .O(gates_190),
   .I0(InputBits[480]),
   .I1(InputBits[196]),
   .I2(InputBits[293]),
   .I3(InputBits[481]),
   .I4(InputBits[339]),
   .I5(InputBits[478])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001000000000000000010101011010000010101111)  
) LUT6_191 (
   .O(gates_191),
   .I0(InputBits[268]),
   .I1(InputBits[321]),
   .I2(InputBits[403]),
   .I3(InputBits[78]),
   .I4(InputBits[17]),
   .I5(InputBits[242])
);
LUT6 #(
   .INIT(64'b0000000001010111000000010101111100000000000000000000000001010000)  
) LUT6_192 (
   .O(gates_192),
   .I0(InputBits[102]),
   .I1(InputBits[448]),
   .I2(InputBits[118]),
   .I3(InputBits[564]),
   .I4(InputBits[90]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0111111100111111000101011111111100001111000000110011111100001000)  
) LUT6_193 (
   .O(gates_193),
   .I0(InputBits[138]),
   .I1(InputBits[428]),
   .I2(InputBits[231]),
   .I3(InputBits[260]),
   .I4(InputBits[283]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001000110010001000101011101011110)  
) LUT6_194 (
   .O(gates_194),
   .I0(InputBits[312]),
   .I1(InputBits[396]),
   .I2(InputBits[94]),
   .I3(InputBits[271]),
   .I4(InputBits[451]),
   .I5(InputBits[572])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100000001100111011101100001001)  
) LUT6_195 (
   .O(gates_195),
   .I0(InputBits[449]),
   .I1(InputBits[544]),
   .I2(InputBits[131]),
   .I3(InputBits[117]),
   .I4(InputBits[525]),
   .I5(InputBits[554])
);
LUT6 #(
   .INIT(64'b0000000010000000000000001111101000000000100110010000000011111101)  
) LUT6_196 (
   .O(gates_196),
   .I0(InputBits[522]),
   .I1(InputBits[446]),
   .I2(InputBits[187]),
   .I3(InputBits[217]),
   .I4(InputBits[488]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0000000001001111000000001001110000000000010101010000000001010100)  
) LUT6_197 (
   .O(gates_197),
   .I0(InputBits[538]),
   .I1(InputBits[368]),
   .I2(InputBits[384]),
   .I3(InputBits[193]),
   .I4(InputBits[342]),
   .I5(InputBits[248])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000011100100000000111111110000000010101010)  
) LUT6_198 (
   .O(gates_198),
   .I0(InputBits[261]),
   .I1(InputBits[381]),
   .I2(InputBits[113]),
   .I3(InputBits[28]),
   .I4(InputBits[407]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110101001000000000000000001111001101010000)  
) LUT6_199 (
   .O(gates_199),
   .I0(InputBits[282]),
   .I1(InputBits[538]),
   .I2(InputBits[308]),
   .I3(InputBits[199]),
   .I4(InputBits[552]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0111000110110001110001001100110100011111001110111100110111011101)  
) LUT6_200 (
   .O(gates_200),
   .I0(InputBits[126]),
   .I1(InputBits[407]),
   .I2(InputBits[377]),
   .I3(InputBits[112]),
   .I4(InputBits[244]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0000010000000100010001000100010000000000000000000001000100010001)  
) LUT6_201 (
   .O(gates_201),
   .I0(InputBits[433]),
   .I1(InputBits[432]),
   .I2(InputBits[162]),
   .I3(InputBits[79]),
   .I4(InputBits[251]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110010001100110011000000110000)  
) LUT6_202 (
   .O(gates_202),
   .I0(InputBits[477]),
   .I1(InputBits[313]),
   .I2(InputBits[525]),
   .I3(InputBits[160]),
   .I4(InputBits[375]),
   .I5(InputBits[574])
);
LUT6 #(
   .INIT(64'b0000000010101010000000001011101100000000111111100000000011111111)  
) LUT6_203 (
   .O(gates_203),
   .I0(InputBits[237]),
   .I1(InputBits[471]),
   .I2(InputBits[188]),
   .I3(InputBits[265]),
   .I4(InputBits[519]),
   .I5(InputBits[515])
);
LUT6 #(
   .INIT(64'b0000011100000101001111110101111100001000000011010010110000010101)  
) LUT6_204 (
   .O(gates_204),
   .I0(InputBits[104]),
   .I1(InputBits[310]),
   .I2(InputBits[70]),
   .I3(InputBits[128]),
   .I4(InputBits[545]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000010000000100000001001101111110100010)  
) LUT6_205 (
   .O(gates_205),
   .I0(InputBits[430]),
   .I1(InputBits[305]),
   .I2(InputBits[435]),
   .I3(InputBits[317]),
   .I4(InputBits[570]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0000001000100010100000100010101100000000000000110010101100110011)  
) LUT6_206 (
   .O(gates_206),
   .I0(InputBits[164]),
   .I1(InputBits[52]),
   .I2(InputBits[447]),
   .I3(InputBits[485]),
   .I4(InputBits[110]),
   .I5(InputBits[425])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010100000000110011001000110011101110)  
) LUT6_207 (
   .O(gates_207),
   .I0(InputBits[249]),
   .I1(InputBits[347]),
   .I2(InputBits[159]),
   .I3(InputBits[151]),
   .I4(InputBits[229]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b0000000001010111000000010001010100000000011101110000000000010011)  
) LUT6_208 (
   .O(gates_208),
   .I0(InputBits[515]),
   .I1(InputBits[386]),
   .I2(InputBits[471]),
   .I3(InputBits[28]),
   .I4(InputBits[319]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000001100000101000101000000000100000010)  
) LUT6_209 (
   .O(gates_209),
   .I0(InputBits[30]),
   .I1(InputBits[332]),
   .I2(InputBits[362]),
   .I3(InputBits[43]),
   .I4(InputBits[296]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b0000010100000101000000000000010000000100000001010000000000000000)  
) LUT6_210 (
   .O(gates_210),
   .I0(InputBits[504]),
   .I1(InputBits[235]),
   .I2(InputBits[48]),
   .I3(InputBits[404]),
   .I4(InputBits[293]),
   .I5(InputBits[358])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000001100110011000010110000)  
) LUT6_211 (
   .O(gates_211),
   .I0(InputBits[442]),
   .I1(InputBits[30]),
   .I2(InputBits[372]),
   .I3(InputBits[386]),
   .I4(InputBits[549]),
   .I5(InputBits[533])
);
LUT6 #(
   .INIT(64'b0000000000001011000000000000000100000000001111110000001000000000)  
) LUT6_212 (
   .O(gates_212),
   .I0(InputBits[351]),
   .I1(InputBits[540]),
   .I2(InputBits[10]),
   .I3(InputBits[266]),
   .I4(InputBits[396]),
   .I5(InputBits[165])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001010100000000000000010000000000000011)  
) LUT6_213 (
   .O(gates_213),
   .I0(InputBits[566]),
   .I1(InputBits[527]),
   .I2(InputBits[511]),
   .I3(InputBits[505]),
   .I4(InputBits[519]),
   .I5(InputBits[451])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000000010011000100100011101100011111)  
) LUT6_214 (
   .O(gates_214),
   .I0(InputBits[36]),
   .I1(InputBits[8]),
   .I2(InputBits[141]),
   .I3(InputBits[37]),
   .I4(InputBits[497]),
   .I5(InputBits[99])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011111111000000111111111100000000)  
) LUT6_215 (
   .O(gates_215),
   .I0(InputBits[159]),
   .I1(InputBits[388]),
   .I2(InputBits[304]),
   .I3(InputBits[366]),
   .I4(InputBits[416]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b1100000000000000010011000000000011111111111011001011111111111111)  
) LUT6_216 (
   .O(gates_216),
   .I0(InputBits[151]),
   .I1(InputBits[272]),
   .I2(InputBits[307]),
   .I3(InputBits[268]),
   .I4(InputBits[355]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0101010100000000010101010000000001010101010101010101010100010101)  
) LUT6_217 (
   .O(gates_217),
   .I0(InputBits[48]),
   .I1(InputBits[405]),
   .I2(InputBits[330]),
   .I3(InputBits[350]),
   .I4(InputBits[162]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010111001100000000000000000000000000010011)  
) LUT6_218 (
   .O(gates_218),
   .I0(InputBits[568]),
   .I1(InputBits[380]),
   .I2(InputBits[546]),
   .I3(InputBits[110]),
   .I4(InputBits[338]),
   .I5(InputBits[283])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000000000001)  
) LUT6_219 (
   .O(gates_219),
   .I0(InputBits[328]),
   .I1(InputBits[534]),
   .I2(InputBits[121]),
   .I3(InputBits[54]),
   .I4(InputBits[552]),
   .I5(InputBits[505])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000100000000000101000000000001010000)  
) LUT6_220 (
   .O(gates_220),
   .I0(InputBits[39]),
   .I1(InputBits[91]),
   .I2(InputBits[311]),
   .I3(InputBits[50]),
   .I4(InputBits[220]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000000100010011000000000001000100000001000000000000000000000000)  
) LUT6_221 (
   .O(gates_221),
   .I0(InputBits[195]),
   .I1(InputBits[97]),
   .I2(InputBits[460]),
   .I3(InputBits[6]),
   .I4(InputBits[375]),
   .I5(InputBits[393])
);
LUT6 #(
   .INIT(64'b0000000000000000010101010001000100000000000000010110010101100101)  
) LUT6_222 (
   .O(gates_222),
   .I0(InputBits[9]),
   .I1(InputBits[239]),
   .I2(InputBits[425]),
   .I3(InputBits[160]),
   .I4(InputBits[566]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000000000000000000100110000001100000001)  
) LUT6_223 (
   .O(gates_223),
   .I0(InputBits[132]),
   .I1(InputBits[147]),
   .I2(InputBits[148]),
   .I3(InputBits[14]),
   .I4(InputBits[119]),
   .I5(InputBits[558])
);
LUT6 #(
   .INIT(64'b0000110000001001110010000000101100000000000010001100111110011011)  
) LUT6_224 (
   .O(gates_224),
   .I0(InputBits[326]),
   .I1(InputBits[257]),
   .I2(InputBits[496]),
   .I3(InputBits[376]),
   .I4(InputBits[527]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0000101100001000000011110000110000001111000011000000111100001100)  
) LUT6_225 (
   .O(gates_225),
   .I0(InputBits[161]),
   .I1(InputBits[244]),
   .I2(InputBits[48]),
   .I3(InputBits[397]),
   .I4(InputBits[497]),
   .I5(InputBits[134])
);
LUT6 #(
   .INIT(64'b0001011111110111001100111100110000110001011111110011001111011011)  
) LUT6_226 (
   .O(gates_226),
   .I0(InputBits[281]),
   .I1(InputBits[502]),
   .I2(InputBits[88]),
   .I3(InputBits[383]),
   .I4(InputBits[236]),
   .I5(InputBits[82])
);
LUT6 #(
   .INIT(64'b0011111000011111001110000011101011111010111110101111101010100010)  
) LUT6_227 (
   .O(gates_227),
   .I0(InputBits[366]),
   .I1(InputBits[440]),
   .I2(InputBits[292]),
   .I3(InputBits[153]),
   .I4(InputBits[202]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010100000000000000000000000000001000)  
) LUT6_228 (
   .O(gates_228),
   .I0(InputBits[35]),
   .I1(InputBits[498]),
   .I2(InputBits[147]),
   .I3(InputBits[4]),
   .I4(InputBits[72]),
   .I5(InputBits[200])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010000011101110000000000100000)  
) LUT6_229 (
   .O(gates_229),
   .I0(InputBits[10]),
   .I1(InputBits[173]),
   .I2(InputBits[423]),
   .I3(InputBits[542]),
   .I4(InputBits[371]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010001000100010000000001010001)  
) LUT6_230 (
   .O(gates_230),
   .I0(InputBits[557]),
   .I1(InputBits[205]),
   .I2(InputBits[116]),
   .I3(InputBits[301]),
   .I4(InputBits[547]),
   .I5(InputBits[529])
);
LUT6 #(
   .INIT(64'b1011101110111010011110101011101100011111101010100011111110101011)  
) LUT6_231 (
   .O(gates_231),
   .I0(InputBits[261]),
   .I1(InputBits[519]),
   .I2(InputBits[452]),
   .I3(InputBits[399]),
   .I4(InputBits[151]),
   .I5(InputBits[466])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000100000000000000010000001100000111)  
) LUT6_232 (
   .O(gates_232),
   .I0(InputBits[517]),
   .I1(InputBits[573]),
   .I2(InputBits[72]),
   .I3(InputBits[360]),
   .I4(InputBits[514]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1111010111110111000101011111111110100110101011111011111110101111)  
) LUT6_233 (
   .O(gates_233),
   .I0(InputBits[444]),
   .I1(InputBits[339]),
   .I2(InputBits[468]),
   .I3(InputBits[475]),
   .I4(InputBits[428]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000110000000100000111)  
) LUT6_234 (
   .O(gates_234),
   .I0(InputBits[43]),
   .I1(InputBits[567]),
   .I2(InputBits[124]),
   .I3(InputBits[288]),
   .I4(InputBits[154]),
   .I5(InputBits[97])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000000000000000000000001010000000000000000)  
) LUT6_235 (
   .O(gates_235),
   .I0(InputBits[505]),
   .I1(InputBits[301]),
   .I2(InputBits[530]),
   .I3(InputBits[19]),
   .I4(InputBits[317]),
   .I5(InputBits[67])
);
LUT6 #(
   .INIT(64'b0000000100000000010111111111101000000001000000101110111111111010)  
) LUT6_236 (
   .O(gates_236),
   .I0(InputBits[373]),
   .I1(InputBits[196]),
   .I2(InputBits[431]),
   .I3(InputBits[285]),
   .I4(InputBits[483]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0000001100000011000000100000000000000010000000110000000000000010)  
) LUT6_237 (
   .O(gates_237),
   .I0(InputBits[445]),
   .I1(InputBits[527]),
   .I2(InputBits[575]),
   .I3(InputBits[273]),
   .I4(InputBits[198]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000111100001011000011110000111100000001000000000000010100000101)  
) LUT6_238 (
   .O(gates_238),
   .I0(InputBits[511]),
   .I1(InputBits[303]),
   .I2(InputBits[25]),
   .I3(InputBits[162]),
   .I4(InputBits[489]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000100000001)  
) LUT6_239 (
   .O(gates_239),
   .I0(InputBits[4]),
   .I1(InputBits[59]),
   .I2(InputBits[72]),
   .I3(InputBits[20]),
   .I4(InputBits[134]),
   .I5(InputBits[123])
);
LUT6 #(
   .INIT(64'b0000000000000000000111010000110000000000000101110000111100111111)  
) LUT6_240 (
   .O(gates_240),
   .I0(InputBits[412]),
   .I1(InputBits[167]),
   .I2(InputBits[10]),
   .I3(InputBits[228]),
   .I4(InputBits[104]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0000000000010001011111110101011100000001000000011000100010001000)  
) LUT6_241 (
   .O(gates_241),
   .I0(InputBits[62]),
   .I1(InputBits[500]),
   .I2(InputBits[412]),
   .I3(InputBits[86]),
   .I4(InputBits[143]),
   .I5(InputBits[261])
);
LUT6 #(
   .INIT(64'b0111000011110111111111011111011100110000101110101111000011110011)  
) LUT6_242 (
   .O(gates_242),
   .I0(InputBits[64]),
   .I1(InputBits[209]),
   .I2(InputBits[237]),
   .I3(InputBits[227]),
   .I4(InputBits[151]),
   .I5(InputBits[286])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000000001000000000011011101)  
) LUT6_243 (
   .O(gates_243),
   .I0(InputBits[52]),
   .I1(InputBits[89]),
   .I2(InputBits[466]),
   .I3(InputBits[565]),
   .I4(InputBits[361]),
   .I5(InputBits[434])
);
LUT6 #(
   .INIT(64'b0000010111011111100011111101111100000000000011000000100011011101)  
) LUT6_244 (
   .O(gates_244),
   .I0(InputBits[330]),
   .I1(InputBits[319]),
   .I2(InputBits[229]),
   .I3(InputBits[102]),
   .I4(InputBits[491]),
   .I5(InputBits[222])
);
LUT6 #(
   .INIT(64'b0000010100000101010101010100010100000000000001010001010101000100)  
) LUT6_245 (
   .O(gates_245),
   .I0(InputBits[433]),
   .I1(InputBits[418]),
   .I2(InputBits[56]),
   .I3(InputBits[268]),
   .I4(InputBits[70]),
   .I5(InputBits[294])
);
LUT6 #(
   .INIT(64'b0000011100000011000000110000001100000011000010110000000100000011)  
) LUT6_246 (
   .O(gates_246),
   .I0(InputBits[154]),
   .I1(InputBits[252]),
   .I2(InputBits[47]),
   .I3(InputBits[112]),
   .I4(InputBits[319]),
   .I5(InputBits[523])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000111111110000000011110011)  
) LUT6_247 (
   .O(gates_247),
   .I0(InputBits[173]),
   .I1(InputBits[497]),
   .I2(InputBits[524]),
   .I3(InputBits[576]),
   .I4(InputBits[259]),
   .I5(InputBits[554])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000001000011010100000101001111)  
) LUT6_248 (
   .O(gates_248),
   .I0(InputBits[460]),
   .I1(InputBits[351]),
   .I2(InputBits[279]),
   .I3(InputBits[240]),
   .I4(InputBits[173]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0000001100000000000000110000000000000001000000000001000100000101)  
) LUT6_249 (
   .O(gates_249),
   .I0(InputBits[509]),
   .I1(InputBits[8]),
   .I2(InputBits[170]),
   .I3(InputBits[246]),
   .I4(InputBits[535]),
   .I5(InputBits[461])
);
LUT6 #(
   .INIT(64'b0000010101010101000000000101010101000101000101010101010100000101)  
) LUT6_250 (
   .O(gates_250),
   .I0(InputBits[123]),
   .I1(InputBits[379]),
   .I2(InputBits[254]),
   .I3(InputBits[383]),
   .I4(InputBits[223]),
   .I5(InputBits[239])
);
LUT6 #(
   .INIT(64'b0010011101100010001000100011011001110000110010000101001111011101)  
) LUT6_251 (
   .O(gates_251),
   .I0(InputBits[184]),
   .I1(InputBits[165]),
   .I2(InputBits[351]),
   .I3(InputBits[243]),
   .I4(InputBits[148]),
   .I5(InputBits[547])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010001010001011101010101011101110)  
) LUT6_252 (
   .O(gates_252),
   .I0(InputBits[394]),
   .I1(InputBits[444]),
   .I2(InputBits[151]),
   .I3(InputBits[184]),
   .I4(InputBits[297]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1101111101010101000100000001000001011101010101010101010001010100)  
) LUT6_253 (
   .O(gates_253),
   .I0(InputBits[100]),
   .I1(InputBits[115]),
   .I2(InputBits[178]),
   .I3(InputBits[476]),
   .I4(InputBits[347]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0101110001010110010101100101110001011100010101100101010001011100)  
) LUT6_254 (
   .O(gates_254),
   .I0(InputBits[10]),
   .I1(InputBits[349]),
   .I2(InputBits[223]),
   .I3(InputBits[209]),
   .I4(InputBits[355]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0100111100001101000011110000111100000000000001000000001000000101)  
) LUT6_255 (
   .O(gates_255),
   .I0(InputBits[485]),
   .I1(InputBits[89]),
   .I2(InputBits[409]),
   .I3(InputBits[411]),
   .I4(InputBits[426]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000010100000000000000000000001100001101)  
) LUT6_256 (
   .O(gates_256),
   .I0(InputBits[149]),
   .I1(InputBits[411]),
   .I2(InputBits[433]),
   .I3(InputBits[526]),
   .I4(InputBits[146]),
   .I5(InputBits[160])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100010011100000000000000000001001000010011)  
) LUT6_257 (
   .O(gates_257),
   .I0(InputBits[383]),
   .I1(InputBits[52]),
   .I2(InputBits[6]),
   .I3(InputBits[232]),
   .I4(InputBits[98]),
   .I5(InputBits[323])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001111000010000000111100001100)  
) LUT6_258 (
   .O(gates_258),
   .I0(InputBits[154]),
   .I1(InputBits[311]),
   .I2(InputBits[531]),
   .I3(InputBits[261]),
   .I4(InputBits[485]),
   .I5(InputBits[530])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000001000000000000000100000001000000010001)  
) LUT6_259 (
   .O(gates_259),
   .I0(InputBits[434]),
   .I1(InputBits[409]),
   .I2(InputBits[157]),
   .I3(InputBits[558]),
   .I4(InputBits[6]),
   .I5(InputBits[135])
);
LUT6 #(
   .INIT(64'b0011010100110100001101010001010000010101000000000101011100010100)  
) LUT6_260 (
   .O(gates_260),
   .I0(InputBits[123]),
   .I1(InputBits[312]),
   .I2(InputBits[245]),
   .I3(InputBits[342]),
   .I4(InputBits[257]),
   .I5(InputBits[321])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110101111100000000000000000000001000011010)  
) LUT6_261 (
   .O(gates_261),
   .I0(InputBits[118]),
   .I1(InputBits[131]),
   .I2(InputBits[478]),
   .I3(InputBits[535]),
   .I4(InputBits[458]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0000000000010011000000000001001100000000001100110001100000010011)  
) LUT6_262 (
   .O(gates_262),
   .I0(InputBits[468]),
   .I1(InputBits[150]),
   .I2(InputBits[411]),
   .I3(InputBits[82]),
   .I4(InputBits[44]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000000000011001100010011001100010000000100010001001100010001)  
) LUT6_263 (
   .O(gates_263),
   .I0(InputBits[277]),
   .I1(InputBits[409]),
   .I2(InputBits[160]),
   .I3(InputBits[183]),
   .I4(InputBits[498]),
   .I5(InputBits[94])
);
LUT6 #(
   .INIT(64'b0101000101010101010100000101000001010101010101010101000101010001)  
) LUT6_264 (
   .O(gates_264),
   .I0(InputBits[554]),
   .I1(InputBits[279]),
   .I2(InputBits[393]),
   .I3(InputBits[403]),
   .I4(InputBits[221]),
   .I5(InputBits[128])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000111100000000000000000000010100000000)  
) LUT6_265 (
   .O(gates_265),
   .I0(InputBits[400]),
   .I1(InputBits[468]),
   .I2(InputBits[506]),
   .I3(InputBits[120]),
   .I4(InputBits[241]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000000111011100000000111101110)  
) LUT6_266 (
   .O(gates_266),
   .I0(InputBits[397]),
   .I1(InputBits[456]),
   .I2(InputBits[208]),
   .I3(InputBits[572]),
   .I4(InputBits[59]),
   .I5(InputBits[21])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000100010100000000000001000000010101000100)  
) LUT6_267 (
   .O(gates_267),
   .I0(InputBits[98]),
   .I1(InputBits[342]),
   .I2(InputBits[37]),
   .I3(InputBits[45]),
   .I4(InputBits[568]),
   .I5(InputBits[261])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100000011000000000000001000000000000001110)  
) LUT6_268 (
   .O(gates_268),
   .I0(InputBits[455]),
   .I1(InputBits[271]),
   .I2(InputBits[482]),
   .I3(InputBits[508]),
   .I4(InputBits[559]),
   .I5(InputBits[133])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001111011100000000000000000000001010100010)  
) LUT6_269 (
   .O(gates_269),
   .I0(InputBits[324]),
   .I1(InputBits[132]),
   .I2(InputBits[42]),
   .I3(InputBits[528]),
   .I4(InputBits[361]),
   .I5(InputBits[235])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000101100000000001100110000000001110111)  
) LUT6_270 (
   .O(gates_270),
   .I0(InputBits[328]),
   .I1(InputBits[516]),
   .I2(InputBits[550]),
   .I3(InputBits[96]),
   .I4(InputBits[427]),
   .I5(InputBits[119])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000111000000010000000000000000)  
) LUT6_271 (
   .O(gates_271),
   .I0(InputBits[297]),
   .I1(InputBits[561]),
   .I2(InputBits[313]),
   .I3(InputBits[179]),
   .I4(InputBits[318]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000000100000000000100010000001000000101000101110001010100010111)  
) LUT6_272 (
   .O(gates_272),
   .I0(InputBits[7]),
   .I1(InputBits[16]),
   .I2(InputBits[46]),
   .I3(InputBits[187]),
   .I4(InputBits[321]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001011100010000000100000011001000010001)  
) LUT6_273 (
   .O(gates_273),
   .I0(InputBits[101]),
   .I1(InputBits[571]),
   .I2(InputBits[381]),
   .I3(InputBits[58]),
   .I4(InputBits[518]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0011111111101111001111111111110100000101000011010000000000000000)  
) LUT6_274 (
   .O(gates_274),
   .I0(InputBits[281]),
   .I1(InputBits[296]),
   .I2(InputBits[484]),
   .I3(InputBits[476]),
   .I4(InputBits[212]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000010000000100000001000000000000000100000001000000000100000011)  
) LUT6_275 (
   .O(gates_275),
   .I0(InputBits[495]),
   .I1(InputBits[424]),
   .I2(InputBits[409]),
   .I3(InputBits[378]),
   .I4(InputBits[150]),
   .I5(InputBits[99])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010000000100010011001100100011)  
) LUT6_276 (
   .O(gates_276),
   .I0(InputBits[89]),
   .I1(InputBits[122]),
   .I2(InputBits[427]),
   .I3(InputBits[430]),
   .I4(InputBits[7]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0000001111111110111110101111100000000001111111111111101011111010)  
) LUT6_277 (
   .O(gates_277),
   .I0(InputBits[345]),
   .I1(InputBits[66]),
   .I2(InputBits[394]),
   .I3(InputBits[40]),
   .I4(InputBits[202]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0001000000000000000000000100000000010000100111110000000010001101)  
) LUT6_278 (
   .O(gates_278),
   .I0(InputBits[105]),
   .I1(InputBits[549]),
   .I2(InputBits[149]),
   .I3(InputBits[218]),
   .I4(InputBits[164]),
   .I5(InputBits[123])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100010001111110001000000111011)  
) LUT6_279 (
   .O(gates_279),
   .I0(InputBits[270]),
   .I1(InputBits[538]),
   .I2(InputBits[454]),
   .I3(InputBits[254]),
   .I4(InputBits[292]),
   .I5(InputBits[99])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001000100000000000000000000000000000101)  
) LUT6_280 (
   .O(gates_280),
   .I0(InputBits[554]),
   .I1(InputBits[566]),
   .I2(InputBits[195]),
   .I3(InputBits[564]),
   .I4(InputBits[512]),
   .I5(InputBits[524])
);
LUT6 #(
   .INIT(64'b0000000100000101000000000000110100000001000011010000000101111101)  
) LUT6_281 (
   .O(gates_281),
   .I0(InputBits[95]),
   .I1(InputBits[141]),
   .I2(InputBits[276]),
   .I3(InputBits[52]),
   .I4(InputBits[485]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000010100000100010101001100)  
) LUT6_282 (
   .O(gates_282),
   .I0(InputBits[567]),
   .I1(InputBits[141]),
   .I2(InputBits[413]),
   .I3(InputBits[120]),
   .I4(InputBits[405]),
   .I5(InputBits[527])
);
LUT6 #(
   .INIT(64'b0000000000010001000000010010001100000000000000010000000000100011)  
) LUT6_283 (
   .O(gates_283),
   .I0(InputBits[221]),
   .I1(InputBits[19]),
   .I2(InputBits[274]),
   .I3(InputBits[504]),
   .I4(InputBits[10]),
   .I5(InputBits[426])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000010000011011100011111111111111111)  
) LUT6_284 (
   .O(gates_284),
   .I0(InputBits[207]),
   .I1(InputBits[477]),
   .I2(InputBits[292]),
   .I3(InputBits[524]),
   .I4(InputBits[250]),
   .I5(InputBits[533])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010000001100010011)  
) LUT6_285 (
   .O(gates_285),
   .I0(InputBits[536]),
   .I1(InputBits[55]),
   .I2(InputBits[86]),
   .I3(InputBits[144]),
   .I4(InputBits[470]),
   .I5(InputBits[122])
);
LUT6 #(
   .INIT(64'b0000011000010111000000000001011100010101000101010001011000010111)  
) LUT6_286 (
   .O(gates_286),
   .I0(InputBits[243]),
   .I1(InputBits[215]),
   .I2(InputBits[70]),
   .I3(InputBits[83]),
   .I4(InputBits[438]),
   .I5(InputBits[184])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000000000010110000101100001011)  
) LUT6_287 (
   .O(gates_287),
   .I0(InputBits[294]),
   .I1(InputBits[299]),
   .I2(InputBits[552]),
   .I3(InputBits[192]),
   .I4(InputBits[548]),
   .I5(InputBits[561])
);
LUT6 #(
   .INIT(64'b0011001101110011101110101111011100110111101100101011101011110010)  
) LUT6_288 (
   .O(gates_288),
   .I0(InputBits[343]),
   .I1(InputBits[149]),
   .I2(InputBits[261]),
   .I3(InputBits[248]),
   .I4(InputBits[142]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b1101111100001010011110110000111100000000000011000011000100011111)  
) LUT6_289 (
   .O(gates_289),
   .I0(InputBits[356]),
   .I1(InputBits[157]),
   .I2(InputBits[521]),
   .I3(InputBits[497]),
   .I4(InputBits[109]),
   .I5(InputBits[165])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000110000000000000110100001000)  
) LUT6_290 (
   .O(gates_290),
   .I0(InputBits[113]),
   .I1(InputBits[35]),
   .I2(InputBits[552]),
   .I3(InputBits[296]),
   .I4(InputBits[356]),
   .I5(InputBits[409])
);
LUT6 #(
   .INIT(64'b1111100011111111111111001111111110000000101110101111110010111110)  
) LUT6_291 (
   .O(gates_291),
   .I0(InputBits[333]),
   .I1(InputBits[325]),
   .I2(InputBits[211]),
   .I3(InputBits[305]),
   .I4(InputBits[380]),
   .I5(InputBits[441])
);
LUT6 #(
   .INIT(64'b0011001100110011000100110010000000110011001000110000001100100000)  
) LUT6_292 (
   .O(gates_292),
   .I0(InputBits[190]),
   .I1(InputBits[532]),
   .I2(InputBits[226]),
   .I3(InputBits[245]),
   .I4(InputBits[223]),
   .I5(InputBits[376])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001000100000000001100010000000010110011)  
) LUT6_293 (
   .O(gates_293),
   .I0(InputBits[207]),
   .I1(InputBits[361]),
   .I2(InputBits[315]),
   .I3(InputBits[122]),
   .I4(InputBits[402]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0101000001000000010101010101010001000000010100000101010101010101)  
) LUT6_294 (
   .O(gates_294),
   .I0(InputBits[73]),
   .I1(InputBits[348]),
   .I2(InputBits[392]),
   .I3(InputBits[429]),
   .I4(InputBits[275]),
   .I5(InputBits[86])
);
LUT6 #(
   .INIT(64'b0000000000110000000000000011000000000000001100000000000000110000)  
) LUT6_295 (
   .O(gates_295),
   .I0(InputBits[459]),
   .I1(InputBits[98]),
   .I2(InputBits[366]),
   .I3(InputBits[3]),
   .I4(InputBits[175]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000001100000000000001000010001100111101)  
) LUT6_296 (
   .O(gates_296),
   .I0(InputBits[57]),
   .I1(InputBits[119]),
   .I2(InputBits[30]),
   .I3(InputBits[430]),
   .I4(InputBits[558]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010011110100000000000000000000000001011000)  
) LUT6_297 (
   .O(gates_297),
   .I0(InputBits[172]),
   .I1(InputBits[66]),
   .I2(InputBits[359]),
   .I3(InputBits[28]),
   .I4(InputBits[3]),
   .I5(InputBits[348])
);
LUT6 #(
   .INIT(64'b0000000100000001000000010000000000000001000000000000000100000000)  
) LUT6_298 (
   .O(gates_298),
   .I0(InputBits[54]),
   .I1(InputBits[337]),
   .I2(InputBits[551]),
   .I3(InputBits[310]),
   .I4(InputBits[188]),
   .I5(InputBits[357])
);
LUT6 #(
   .INIT(64'b0000001000000011000000110000001100000000000100010001001100010101)  
) LUT6_299 (
   .O(gates_299),
   .I0(InputBits[133]),
   .I1(InputBits[410]),
   .I2(InputBits[195]),
   .I3(InputBits[87]),
   .I4(InputBits[230]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000011100100000000000100001111110011111101)  
) LUT6_300 (
   .O(gates_300),
   .I0(InputBits[149]),
   .I1(InputBits[502]),
   .I2(InputBits[423]),
   .I3(InputBits[77]),
   .I4(InputBits[565]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000001110111000000000000010100000000111111110000001010001101)  
) LUT6_301 (
   .O(gates_301),
   .I0(InputBits[403]),
   .I1(InputBits[44]),
   .I2(InputBits[86]),
   .I3(InputBits[528]),
   .I4(InputBits[370]),
   .I5(InputBits[469])
);
LUT6 #(
   .INIT(64'b0000000000000000111111111111111100000000100000001010101110101011)  
) LUT6_302 (
   .O(gates_302),
   .I0(InputBits[419]),
   .I1(InputBits[304]),
   .I2(InputBits[160]),
   .I3(InputBits[302]),
   .I4(InputBits[51]),
   .I5(InputBits[248])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000010110000000000001011)  
) LUT6_303 (
   .O(gates_303),
   .I0(InputBits[263]),
   .I1(InputBits[58]),
   .I2(InputBits[147]),
   .I3(InputBits[265]),
   .I4(InputBits[412]),
   .I5(InputBits[410])
);
LUT6 #(
   .INIT(64'b0000001100000011001100110010000000000011000000110000001000000010)  
) LUT6_304 (
   .O(gates_304),
   .I0(InputBits[224]),
   .I1(InputBits[4]),
   .I2(InputBits[434]),
   .I3(InputBits[114]),
   .I4(InputBits[238]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0000000000000000000001001000101000000000101010101010111011111111)  
) LUT6_305 (
   .O(gates_305),
   .I0(InputBits[319]),
   .I1(InputBits[398]),
   .I2(InputBits[185]),
   .I3(InputBits[495]),
   .I4(InputBits[144]),
   .I5(InputBits[508])
);
LUT6 #(
   .INIT(64'b1111111101010000111110110000000110111111010101011011011101010101)  
) LUT6_306 (
   .O(gates_306),
   .I0(InputBits[495]),
   .I1(InputBits[59]),
   .I2(InputBits[160]),
   .I3(InputBits[222]),
   .I4(InputBits[440]),
   .I5(InputBits[469])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000001100010001)  
) LUT6_307 (
   .O(gates_307),
   .I0(InputBits[512]),
   .I1(InputBits[250]),
   .I2(InputBits[508]),
   .I3(InputBits[548]),
   .I4(InputBits[56]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000110000000000000000000000000000011100)  
) LUT6_308 (
   .O(gates_308),
   .I0(InputBits[307]),
   .I1(InputBits[284]),
   .I2(InputBits[218]),
   .I3(InputBits[289]),
   .I4(InputBits[534]),
   .I5(InputBits[174])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000001000111000001110)  
) LUT6_309 (
   .O(gates_309),
   .I0(InputBits[164]),
   .I1(InputBits[186]),
   .I2(InputBits[99]),
   .I3(InputBits[282]),
   .I4(InputBits[231]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0000110100010001111100101110000010101111010111111111111111111101)  
) LUT6_310 (
   .O(gates_310),
   .I0(InputBits[413]),
   .I1(InputBits[327]),
   .I2(InputBits[309]),
   .I3(InputBits[139]),
   .I4(InputBits[501]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000010110000000000011100)  
) LUT6_311 (
   .O(gates_311),
   .I0(InputBits[31]),
   .I1(InputBits[501]),
   .I2(InputBits[288]),
   .I3(InputBits[573]),
   .I4(InputBits[430]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0000000000000101010100000000000001000000000001011101000000000010)  
) LUT6_312 (
   .O(gates_312),
   .I0(InputBits[550]),
   .I1(InputBits[327]),
   .I2(InputBits[501]),
   .I3(InputBits[501]),
   .I4(InputBits[223]),
   .I5(InputBits[64])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000001000000000000011110000000000001111)  
) LUT6_313 (
   .O(gates_313),
   .I0(InputBits[476]),
   .I1(InputBits[516]),
   .I2(InputBits[533]),
   .I3(InputBits[28]),
   .I4(InputBits[158]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100000001000000000000000000000111000101110)  
) LUT6_314 (
   .O(gates_314),
   .I0(InputBits[343]),
   .I1(InputBits[408]),
   .I2(InputBits[544]),
   .I3(InputBits[463]),
   .I4(InputBits[553]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b0010000000000000011101100111001000110011000100000110001101110111)  
) LUT6_315 (
   .O(gates_315),
   .I0(InputBits[235]),
   .I1(InputBits[10]),
   .I2(InputBits[399]),
   .I3(InputBits[463]),
   .I4(InputBits[16]),
   .I5(InputBits[355])
);
LUT6 #(
   .INIT(64'b0000000100000111000000110000111100000000000000000000000100000111)  
) LUT6_316 (
   .O(gates_316),
   .I0(InputBits[485]),
   .I1(InputBits[491]),
   .I2(InputBits[74]),
   .I3(InputBits[279]),
   .I4(InputBits[149]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0101000000010000010001000101000000010000010100000100010001010000)  
) LUT6_317 (
   .O(gates_317),
   .I0(InputBits[124]),
   .I1(InputBits[180]),
   .I2(InputBits[340]),
   .I3(InputBits[89]),
   .I4(InputBits[323]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000001000000000000000010000000001010011)  
) LUT6_318 (
   .O(gates_318),
   .I0(InputBits[10]),
   .I1(InputBits[482]),
   .I2(InputBits[42]),
   .I3(InputBits[409]),
   .I4(InputBits[118]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0001000000110001000100010001000100000000000100010001000100010011)  
) LUT6_319 (
   .O(gates_319),
   .I0(InputBits[540]),
   .I1(InputBits[313]),
   .I2(InputBits[501]),
   .I3(InputBits[219]),
   .I4(InputBits[131]),
   .I5(InputBits[174])
);
LUT6 #(
   .INIT(64'b0000000000000000011101011111111100000000000000001111110011111100)  
) LUT6_320 (
   .O(gates_320),
   .I0(InputBits[450]),
   .I1(InputBits[286]),
   .I2(InputBits[268]),
   .I3(InputBits[496]),
   .I4(InputBits[22]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0000111101001111101011110110111100101110011011101010101011101110)  
) LUT6_321 (
   .O(gates_321),
   .I0(InputBits[396]),
   .I1(InputBits[391]),
   .I2(InputBits[538]),
   .I3(InputBits[328]),
   .I4(InputBits[477]),
   .I5(InputBits[370])
);
LUT6 #(
   .INIT(64'b0000011100011111011111111111110101001101010011011110110011101100)  
) LUT6_322 (
   .O(gates_322),
   .I0(InputBits[204]),
   .I1(InputBits[345]),
   .I2(InputBits[141]),
   .I3(InputBits[162]),
   .I4(InputBits[454]),
   .I5(InputBits[222])
);
LUT6 #(
   .INIT(64'b0000000000000111000000101000001000000000110010100000000000001010)  
) LUT6_323 (
   .O(gates_323),
   .I0(InputBits[224]),
   .I1(InputBits[196]),
   .I2(InputBits[149]),
   .I3(InputBits[314]),
   .I4(InputBits[442]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010111010100010001)  
) LUT6_324 (
   .O(gates_324),
   .I0(InputBits[229]),
   .I1(InputBits[100]),
   .I2(InputBits[320]),
   .I3(InputBits[210]),
   .I4(InputBits[192]),
   .I5(InputBits[277])
);
LUT6 #(
   .INIT(64'b0000000000001100000000010000111100000010000011000000001100001111)  
) LUT6_325 (
   .O(gates_325),
   .I0(InputBits[306]),
   .I1(InputBits[285]),
   .I2(InputBits[556]),
   .I3(InputBits[527]),
   .I4(InputBits[275]),
   .I5(InputBits[175])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000101111101010001)  
) LUT6_326 (
   .O(gates_326),
   .I0(InputBits[354]),
   .I1(InputBits[489]),
   .I2(InputBits[480]),
   .I3(InputBits[415]),
   .I4(InputBits[433]),
   .I5(InputBits[385])
);
LUT6 #(
   .INIT(64'b0000000000001110000000000000110000000010000011100000000000000100)  
) LUT6_327 (
   .O(gates_327),
   .I0(InputBits[211]),
   .I1(InputBits[69]),
   .I2(InputBits[530]),
   .I3(InputBits[53]),
   .I4(InputBits[283]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b0000000010000100000000000100000000000000110100000100000101010001)  
) LUT6_328 (
   .O(gates_328),
   .I0(InputBits[79]),
   .I1(InputBits[233]),
   .I2(InputBits[326]),
   .I3(InputBits[71]),
   .I4(InputBits[58]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0000001100000011000000000001000000000010000011110000000000010000)  
) LUT6_329 (
   .O(gates_329),
   .I0(InputBits[204]),
   .I1(InputBits[144]),
   .I2(InputBits[17]),
   .I3(InputBits[159]),
   .I4(InputBits[212]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b1000010110101111011101110001111100100101001011110111010100110000)  
) LUT6_330 (
   .O(gates_330),
   .I0(InputBits[474]),
   .I1(InputBits[380]),
   .I2(InputBits[476]),
   .I3(InputBits[325]),
   .I4(InputBits[383]),
   .I5(InputBits[247])
);
LUT6 #(
   .INIT(64'b0000001100001111000000110000011100000000000001010000000000010101)  
) LUT6_331 (
   .O(gates_331),
   .I0(InputBits[251]),
   .I1(InputBits[243]),
   .I2(InputBits[29]),
   .I3(InputBits[509]),
   .I4(InputBits[115]),
   .I5(InputBits[222])
);
LUT6 #(
   .INIT(64'b0001000000000000000100010001000100010001000000000001000100000000)  
) LUT6_332 (
   .O(gates_332),
   .I0(InputBits[169]),
   .I1(InputBits[433]),
   .I2(InputBits[197]),
   .I3(InputBits[420]),
   .I4(InputBits[231]),
   .I5(InputBits[440])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000000000000000100100011)  
) LUT6_333 (
   .O(gates_333),
   .I0(InputBits[440]),
   .I1(InputBits[22]),
   .I2(InputBits[512]),
   .I3(InputBits[571]),
   .I4(InputBits[193]),
   .I5(InputBits[69])
);
LUT6 #(
   .INIT(64'b1010001000111110000010100010001101111111110011110010001100100011)  
) LUT6_334 (
   .O(gates_334),
   .I0(InputBits[476]),
   .I1(InputBits[498]),
   .I2(InputBits[56]),
   .I3(InputBits[466]),
   .I4(InputBits[187]),
   .I5(InputBits[435])
);
LUT6 #(
   .INIT(64'b0011011100010000111111111111111111001110010011001100111011011111)  
) LUT6_335 (
   .O(gates_335),
   .I0(InputBits[63]),
   .I1(InputBits[421]),
   .I2(InputBits[209]),
   .I3(InputBits[131]),
   .I4(InputBits[518]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000101010100000000010001010000000001010100)  
) LUT6_336 (
   .O(gates_336),
   .I0(InputBits[24]),
   .I1(InputBits[309]),
   .I2(InputBits[406]),
   .I3(InputBits[21]),
   .I4(InputBits[476]),
   .I5(InputBits[248])
);
LUT6 #(
   .INIT(64'b0101111101011111110001011111111100010011000111100101111111101010)  
) LUT6_337 (
   .O(gates_337),
   .I0(InputBits[525]),
   .I1(InputBits[347]),
   .I2(InputBits[220]),
   .I3(InputBits[364]),
   .I4(InputBits[441]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0000000000011110000000000010010000000000001011110000000000110100)  
) LUT6_338 (
   .O(gates_338),
   .I0(InputBits[210]),
   .I1(InputBits[141]),
   .I2(InputBits[503]),
   .I3(InputBits[25]),
   .I4(InputBits[295]),
   .I5(InputBits[403])
);
LUT6 #(
   .INIT(64'b0000000000000000111111111100110100000000000000001111111111001111)  
) LUT6_339 (
   .O(gates_339),
   .I0(InputBits[87]),
   .I1(InputBits[246]),
   .I2(InputBits[401]),
   .I3(InputBits[392]),
   .I4(InputBits[556]),
   .I5(InputBits[186])
);
LUT6 #(
   .INIT(64'b0101010011011011110111111101111100000000101010100000100000001010)  
) LUT6_340 (
   .O(gates_340),
   .I0(InputBits[383]),
   .I1(InputBits[400]),
   .I2(InputBits[61]),
   .I3(InputBits[436]),
   .I4(InputBits[472]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0100000000010001000000000100010001110000111101110101001101110101)  
) LUT6_341 (
   .O(gates_341),
   .I0(InputBits[16]),
   .I1(InputBits[111]),
   .I2(InputBits[394]),
   .I3(InputBits[254]),
   .I4(InputBits[425]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b0000000001111111000000000001110100001100101111110000110001111111)  
) LUT6_342 (
   .O(gates_342),
   .I0(InputBits[136]),
   .I1(InputBits[261]),
   .I2(InputBits[42]),
   .I3(InputBits[536]),
   .I4(InputBits[439]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000000000000000000010011)  
) LUT6_343 (
   .O(gates_343),
   .I0(InputBits[184]),
   .I1(InputBits[409]),
   .I2(InputBits[300]),
   .I3(InputBits[481]),
   .I4(InputBits[560]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000100000011110010011011101111101100110000)  
) LUT6_344 (
   .O(gates_344),
   .I0(InputBits[161]),
   .I1(InputBits[79]),
   .I2(InputBits[417]),
   .I3(InputBits[419]),
   .I4(InputBits[480]),
   .I5(InputBits[194])
);
LUT6 #(
   .INIT(64'b0001010001000001010101010001010101010001010110110001000001010010)  
) LUT6_345 (
   .O(gates_345),
   .I0(InputBits[266]),
   .I1(InputBits[521]),
   .I2(InputBits[418]),
   .I3(InputBits[440]),
   .I4(InputBits[522]),
   .I5(InputBits[190])
);
LUT6 #(
   .INIT(64'b0000000011101110100000101100111000000000111111110000010011011111)  
) LUT6_346 (
   .O(gates_346),
   .I0(InputBits[210]),
   .I1(InputBits[340]),
   .I2(InputBits[112]),
   .I3(InputBits[218]),
   .I4(InputBits[64]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0000001000000001001100110001001100000000000000000000001100000011)  
) LUT6_347 (
   .O(gates_347),
   .I0(InputBits[163]),
   .I1(InputBits[433]),
   .I2(InputBits[125]),
   .I3(InputBits[283]),
   .I4(InputBits[29]),
   .I5(InputBits[375])
);
LUT6 #(
   .INIT(64'b0010110011101010001010111000101111111010111110101011001011111011)  
) LUT6_348 (
   .O(gates_348),
   .I0(InputBits[343]),
   .I1(InputBits[354]),
   .I2(InputBits[246]),
   .I3(InputBits[108]),
   .I4(InputBits[283]),
   .I5(InputBits[477])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000101000000010000000000011100000001010001)  
) LUT6_349 (
   .O(gates_349),
   .I0(InputBits[124]),
   .I1(InputBits[522]),
   .I2(InputBits[223]),
   .I3(InputBits[148]),
   .I4(InputBits[527]),
   .I5(InputBits[207])
);
LUT6 #(
   .INIT(64'b0000000001011101000000000000110000000000110011110000000001001101)  
) LUT6_350 (
   .O(gates_350),
   .I0(InputBits[435]),
   .I1(InputBits[342]),
   .I2(InputBits[538]),
   .I3(InputBits[145]),
   .I4(InputBits[225]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0011000000100000000000000000000100110011001100110111111000000011)  
) LUT6_351 (
   .O(gates_351),
   .I0(InputBits[297]),
   .I1(InputBits[6]),
   .I2(InputBits[327]),
   .I3(InputBits[375]),
   .I4(InputBits[283]),
   .I5(InputBits[278])
);
LUT6 #(
   .INIT(64'b0001000000100000000100010010011111010000000000000101011100100010)  
) LUT6_352 (
   .O(gates_352),
   .I0(InputBits[524]),
   .I1(InputBits[429]),
   .I2(InputBits[512]),
   .I3(InputBits[334]),
   .I4(InputBits[536]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0000000000000000010100010000000000000000000000000101000101010111)  
) LUT6_353 (
   .O(gates_353),
   .I0(InputBits[537]),
   .I1(InputBits[58]),
   .I2(InputBits[174]),
   .I3(InputBits[471]),
   .I4(InputBits[289]),
   .I5(InputBits[520])
);
LUT6 #(
   .INIT(64'b0001001100010000001100010001000000110011001110110011001100001011)  
) LUT6_354 (
   .O(gates_354),
   .I0(InputBits[90]),
   .I1(InputBits[520]),
   .I2(InputBits[37]),
   .I3(InputBits[39]),
   .I4(InputBits[155]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001001100000000000000000000000000010000)  
) LUT6_355 (
   .O(gates_355),
   .I0(InputBits[196]),
   .I1(InputBits[529]),
   .I2(InputBits[336]),
   .I3(InputBits[553]),
   .I4(InputBits[540]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000000000000001000000110011001100000000000000000000000000000001)  
) LUT6_356 (
   .O(gates_356),
   .I0(InputBits[83]),
   .I1(InputBits[529]),
   .I2(InputBits[104]),
   .I3(InputBits[300]),
   .I4(InputBits[29]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0000000001010101010000000101010100010001010101010101000101010101)  
) LUT6_357 (
   .O(gates_357),
   .I0(InputBits[25]),
   .I1(InputBits[57]),
   .I2(InputBits[382]),
   .I3(InputBits[205]),
   .I4(InputBits[186]),
   .I5(InputBits[56])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000111000000111000101111110111111111)  
) LUT6_358 (
   .O(gates_358),
   .I0(InputBits[445]),
   .I1(InputBits[439]),
   .I2(InputBits[200]),
   .I3(InputBits[512]),
   .I4(InputBits[514]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0000000000000000101111111010111100000000000000000010101010101011)  
) LUT6_359 (
   .O(gates_359),
   .I0(InputBits[221]),
   .I1(InputBits[129]),
   .I2(InputBits[173]),
   .I3(InputBits[330]),
   .I4(InputBits[532]),
   .I5(InputBits[258])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000110011000001111111111111)  
) LUT6_360 (
   .O(gates_360),
   .I0(InputBits[233]),
   .I1(InputBits[153]),
   .I2(InputBits[157]),
   .I3(InputBits[300]),
   .I4(InputBits[107]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b1010000010110000111110111111101110100001101000001111111111111011)  
) LUT6_361 (
   .O(gates_361),
   .I0(InputBits[375]),
   .I1(InputBits[81]),
   .I2(InputBits[406]),
   .I3(InputBits[444]),
   .I4(InputBits[277]),
   .I5(InputBits[388])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000111111000000000000000000000000011111110)  
) LUT6_362 (
   .O(gates_362),
   .I0(InputBits[295]),
   .I1(InputBits[246]),
   .I2(InputBits[478]),
   .I3(InputBits[193]),
   .I4(InputBits[146]),
   .I5(InputBits[436])
);
LUT6 #(
   .INIT(64'b0000000000100011000000000010001100000000001100110000000000101011)  
) LUT6_363 (
   .O(gates_363),
   .I0(InputBits[246]),
   .I1(InputBits[574]),
   .I2(InputBits[126]),
   .I3(InputBits[409]),
   .I4(InputBits[467]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000001010000000000000001)  
) LUT6_364 (
   .O(gates_364),
   .I0(InputBits[489]),
   .I1(InputBits[544]),
   .I2(InputBits[482]),
   .I3(InputBits[484]),
   .I4(InputBits[569]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0000000111011101000001010101110100000100010011110000010001001101)  
) LUT6_365 (
   .O(gates_365),
   .I0(InputBits[10]),
   .I1(InputBits[374]),
   .I2(InputBits[251]),
   .I3(InputBits[147]),
   .I4(InputBits[206]),
   .I5(InputBits[319])
);
LUT6 #(
   .INIT(64'b0100000000010001111111111111111100010000010101001111100011111100)  
) LUT6_366 (
   .O(gates_366),
   .I0(InputBits[339]),
   .I1(InputBits[325]),
   .I2(InputBits[374]),
   .I3(InputBits[298]),
   .I4(InputBits[78]),
   .I5(InputBits[261])
);
LUT6 #(
   .INIT(64'b0000010000000001111111111111111100001110000000001111001011110011)  
) LUT6_367 (
   .O(gates_367),
   .I0(InputBits[364]),
   .I1(InputBits[207]),
   .I2(InputBits[261]),
   .I3(InputBits[451]),
   .I4(InputBits[9]),
   .I5(InputBits[393])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010001100001101100011100001111110111111)  
) LUT6_368 (
   .O(gates_368),
   .I0(InputBits[261]),
   .I1(InputBits[165]),
   .I2(InputBits[278]),
   .I3(InputBits[68]),
   .I4(InputBits[104]),
   .I5(InputBits[218])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110010001000000010000000100010001000100010)  
) LUT6_369 (
   .O(gates_369),
   .I0(InputBits[342]),
   .I1(InputBits[48]),
   .I2(InputBits[87]),
   .I3(InputBits[365]),
   .I4(InputBits[564]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b0000001000001010000000100000101000000101000000010000000000000000)  
) LUT6_370 (
   .O(gates_370),
   .I0(InputBits[478]),
   .I1(InputBits[126]),
   .I2(InputBits[555]),
   .I3(InputBits[33]),
   .I4(InputBits[368]),
   .I5(InputBits[478])
);
LUT6 #(
   .INIT(64'b0000000100000011000000000000001100100011001000100011001100110011)  
) LUT6_371 (
   .O(gates_371),
   .I0(InputBits[244]),
   .I1(InputBits[559]),
   .I2(InputBits[387]),
   .I3(InputBits[438]),
   .I4(InputBits[130]),
   .I5(InputBits[548])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011000000110000000000000000)  
) LUT6_372 (
   .O(gates_372),
   .I0(InputBits[475]),
   .I1(InputBits[505]),
   .I2(InputBits[289]),
   .I3(InputBits[427]),
   .I4(InputBits[286]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0000000100000011000100100000001000000001000000110000000000101111)  
) LUT6_373 (
   .O(gates_373),
   .I0(InputBits[370]),
   .I1(InputBits[562]),
   .I2(InputBits[338]),
   .I3(InputBits[541]),
   .I4(InputBits[311]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000001000001010000000000000101)  
) LUT6_374 (
   .O(gates_374),
   .I0(InputBits[47]),
   .I1(InputBits[55]),
   .I2(InputBits[289]),
   .I3(InputBits[469]),
   .I4(InputBits[157]),
   .I5(InputBits[498])
);
LUT6 #(
   .INIT(64'b0011000100100000001100111011101100100011001000100011101110101011)  
) LUT6_375 (
   .O(gates_375),
   .I0(InputBits[166]),
   .I1(InputBits[534]),
   .I2(InputBits[401]),
   .I3(InputBits[176]),
   .I4(InputBits[83]),
   .I5(InputBits[162])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000001100000000000000000001001100000011)  
) LUT6_376 (
   .O(gates_376),
   .I0(InputBits[213]),
   .I1(InputBits[47]),
   .I2(InputBits[100]),
   .I3(InputBits[175]),
   .I4(InputBits[276]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0000000001000000000000010000000100000101010100010000010101000101)  
) LUT6_377 (
   .O(gates_377),
   .I0(InputBits[26]),
   .I1(InputBits[519]),
   .I2(InputBits[568]),
   .I3(InputBits[89]),
   .I4(InputBits[473]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0000000100000000000001110010011000000001000000010000010100100010)  
) LUT6_378 (
   .O(gates_378),
   .I0(InputBits[431]),
   .I1(InputBits[315]),
   .I2(InputBits[33]),
   .I3(InputBits[247]),
   .I4(InputBits[526]),
   .I5(InputBits[404])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000101011100000000000100000000000001010110)  
) LUT6_379 (
   .O(gates_379),
   .I0(InputBits[480]),
   .I1(InputBits[292]),
   .I2(InputBits[340]),
   .I3(InputBits[193]),
   .I4(InputBits[483]),
   .I5(InputBits[431])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000100000001000010101)  
) LUT6_380 (
   .O(gates_380),
   .I0(InputBits[173]),
   .I1(InputBits[95]),
   .I2(InputBits[45]),
   .I3(InputBits[573]),
   .I4(InputBits[59]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b0000001100100010000111110011111100000100001100000001111100110001)  
) LUT6_381 (
   .O(gates_381),
   .I0(InputBits[513]),
   .I1(InputBits[54]),
   .I2(InputBits[68]),
   .I3(InputBits[454]),
   .I4(InputBits[228]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b0000000001000100000000000000000001010100010100001101011111111110)  
) LUT6_382 (
   .O(gates_382),
   .I0(InputBits[95]),
   .I1(InputBits[421]),
   .I2(InputBits[345]),
   .I3(InputBits[388]),
   .I4(InputBits[161]),
   .I5(InputBits[170])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000000000000000000000100)  
) LUT6_383 (
   .O(gates_383),
   .I0(InputBits[482]),
   .I1(InputBits[374]),
   .I2(InputBits[560]),
   .I3(InputBits[553]),
   .I4(InputBits[561]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010001000100000000000000000011001111110110)  
) LUT6_384 (
   .O(gates_384),
   .I0(InputBits[239]),
   .I1(InputBits[384]),
   .I2(InputBits[343]),
   .I3(InputBits[143]),
   .I4(InputBits[76]),
   .I5(InputBits[119])
);
LUT6 #(
   .INIT(64'b0000000100000001000011110101111100000001000100100000011101111111)  
) LUT6_385 (
   .O(gates_385),
   .I0(InputBits[38]),
   .I1(InputBits[492]),
   .I2(InputBits[267]),
   .I3(InputBits[43]),
   .I4(InputBits[251]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0000101000001010000000100001101000001010000010100000001100000011)  
) LUT6_386 (
   .O(gates_386),
   .I0(InputBits[247]),
   .I1(InputBits[127]),
   .I2(InputBits[266]),
   .I3(InputBits[87]),
   .I4(InputBits[423]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0000000000000000010001010001000101000101010001010101110111010111)  
) LUT6_387 (
   .O(gates_387),
   .I0(InputBits[569]),
   .I1(InputBits[364]),
   .I2(InputBits[105]),
   .I3(InputBits[388]),
   .I4(InputBits[515]),
   .I5(InputBits[54])
);
LUT6 #(
   .INIT(64'b0100110010111111111111001111111100000000011110110110110011111101)  
) LUT6_388 (
   .O(gates_388),
   .I0(InputBits[331]),
   .I1(InputBits[350]),
   .I2(InputBits[238]),
   .I3(InputBits[279]),
   .I4(InputBits[173]),
   .I5(InputBits[319])
);
LUT6 #(
   .INIT(64'b0000000100000101010101010101010100010001010100010101000001010101)  
) LUT6_389 (
   .O(gates_389),
   .I0(InputBits[482]),
   .I1(InputBits[134]),
   .I2(InputBits[334]),
   .I3(InputBits[448]),
   .I4(InputBits[288]),
   .I5(InputBits[272])
);
LUT6 #(
   .INIT(64'b0101010101010001010101010101010101010101010101110000010001010110)  
) LUT6_390 (
   .O(gates_390),
   .I0(InputBits[360]),
   .I1(InputBits[142]),
   .I2(InputBits[212]),
   .I3(InputBits[139]),
   .I4(InputBits[393]),
   .I5(InputBits[269])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000100110100000100010001000000000001001110)  
) LUT6_391 (
   .O(gates_391),
   .I0(InputBits[168]),
   .I1(InputBits[398]),
   .I2(InputBits[195]),
   .I3(InputBits[484]),
   .I4(InputBits[100]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010110000100100001111011111010111)  
) LUT6_392 (
   .O(gates_392),
   .I0(InputBits[207]),
   .I1(InputBits[470]),
   .I2(InputBits[525]),
   .I3(InputBits[233]),
   .I4(InputBits[299]),
   .I5(InputBits[573])
);
LUT6 #(
   .INIT(64'b0000000010111111001000100000000100000000111111110101000100010001)  
) LUT6_393 (
   .O(gates_393),
   .I0(InputBits[377]),
   .I1(InputBits[81]),
   .I2(InputBits[161]),
   .I3(InputBits[16]),
   .I4(InputBits[285]),
   .I5(InputBits[376])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000100010000000000000100010000000001000101)  
) LUT6_394 (
   .O(gates_394),
   .I0(InputBits[560]),
   .I1(InputBits[503]),
   .I2(InputBits[125]),
   .I3(InputBits[73]),
   .I4(InputBits[314]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0000000010101111000000000011001100000000111111110000001110110011)  
) LUT6_395 (
   .O(gates_395),
   .I0(InputBits[114]),
   .I1(InputBits[129]),
   .I2(InputBits[191]),
   .I3(InputBits[16]),
   .I4(InputBits[223]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000100001111000011100001111100011111)  
) LUT6_396 (
   .O(gates_396),
   .I0(InputBits[259]),
   .I1(InputBits[287]),
   .I2(InputBits[10]),
   .I3(InputBits[375]),
   .I4(InputBits[127]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1001010011110000110101001111110111100100111101001101010011111100)  
) LUT6_397 (
   .O(gates_397),
   .I0(InputBits[299]),
   .I1(InputBits[319]),
   .I2(InputBits[421]),
   .I3(InputBits[111]),
   .I4(InputBits[204]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b0000000100000000000111000000110100000001000000000000111100001101)  
) LUT6_398 (
   .O(gates_398),
   .I0(InputBits[516]),
   .I1(InputBits[263]),
   .I2(InputBits[171]),
   .I3(InputBits[422]),
   .I4(InputBits[124]),
   .I5(InputBits[488])
);
LUT6 #(
   .INIT(64'b0010001000000000011101010001000110100011000000001111111101010011)  
) LUT6_399 (
   .O(gates_399),
   .I0(InputBits[545]),
   .I1(InputBits[355]),
   .I2(InputBits[161]),
   .I3(InputBits[295]),
   .I4(InputBits[275]),
   .I5(InputBits[462])
);
LUT6 #(
   .INIT(64'b0000001101010101000001111111111000001101000010000000110101010000)  
) LUT6_400 (
   .O(gates_400),
   .I0(InputBits[63]),
   .I1(InputBits[351]),
   .I2(InputBits[384]),
   .I3(InputBits[364]),
   .I4(InputBits[151]),
   .I5(InputBits[383])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000100000000000000000000001100001111)  
) LUT6_401 (
   .O(gates_401),
   .I0(InputBits[104]),
   .I1(InputBits[277]),
   .I2(InputBits[27]),
   .I3(InputBits[492]),
   .I4(InputBits[265]),
   .I5(InputBits[517])
);
LUT6 #(
   .INIT(64'b0111001100000010001100110011001000110011001000100011001100010010)  
) LUT6_402 (
   .O(gates_402),
   .I0(InputBits[392]),
   .I1(InputBits[242]),
   .I2(InputBits[316]),
   .I3(InputBits[294]),
   .I4(InputBits[302]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0000000100000001000000010000000100010001010100000001000101010101)  
) LUT6_403 (
   .O(gates_403),
   .I0(InputBits[553]),
   .I1(InputBits[96]),
   .I2(InputBits[143]),
   .I3(InputBits[388]),
   .I4(InputBits[330]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0000010100000101000000010000000100000101001001110111010100100111)  
) LUT6_404 (
   .O(gates_404),
   .I0(InputBits[526]),
   .I1(InputBits[68]),
   .I2(InputBits[127]),
   .I3(InputBits[117]),
   .I4(InputBits[179]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0000000001010101000000000011011100010000011111010000000110111101)  
) LUT6_405 (
   .O(gates_405),
   .I0(InputBits[515]),
   .I1(InputBits[68]),
   .I2(InputBits[292]),
   .I3(InputBits[266]),
   .I4(InputBits[330]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000000011111111001100111111111101000000111110100011000111111011)  
) LUT6_406 (
   .O(gates_406),
   .I0(InputBits[187]),
   .I1(InputBits[449]),
   .I2(InputBits[334]),
   .I3(InputBits[278]),
   .I4(InputBits[474]),
   .I5(InputBits[309])
);
LUT6 #(
   .INIT(64'b0000000001000000010001000100000000000000000000000000010000000101)  
) LUT6_407 (
   .O(gates_407),
   .I0(InputBits[193]),
   .I1(InputBits[453]),
   .I2(InputBits[330]),
   .I3(InputBits[152]),
   .I4(InputBits[28]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001010001111111011111010111000010001)  
) LUT6_408 (
   .O(gates_408),
   .I0(InputBits[474]),
   .I1(InputBits[80]),
   .I2(InputBits[55]),
   .I3(InputBits[500]),
   .I4(InputBits[341]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001001010010111000001101000111000)  
) LUT6_409 (
   .O(gates_409),
   .I0(InputBits[523]),
   .I1(InputBits[89]),
   .I2(InputBits[93]),
   .I3(InputBits[423]),
   .I4(InputBits[157]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0000000001100011000000000111001000000000011111110000000011110010)  
) LUT6_410 (
   .O(gates_410),
   .I0(InputBits[224]),
   .I1(InputBits[55]),
   .I2(InputBits[324]),
   .I3(InputBits[385]),
   .I4(InputBits[235]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0011001111111111001100110011011100100000010100100001001100010011)  
) LUT6_411 (
   .O(gates_411),
   .I0(InputBits[499]),
   .I1(InputBits[514]),
   .I2(InputBits[156]),
   .I3(InputBits[435]),
   .I4(InputBits[465]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000010100000110)  
) LUT6_412 (
   .O(gates_412),
   .I0(InputBits[572]),
   .I1(InputBits[44]),
   .I2(InputBits[73]),
   .I3(InputBits[202]),
   .I4(InputBits[122]),
   .I5(InputBits[123])
);
LUT6 #(
   .INIT(64'b0101010101010101000000000001100000010111011101110000001100011011)  
) LUT6_413 (
   .O(gates_413),
   .I0(InputBits[312]),
   .I1(InputBits[515]),
   .I2(InputBits[477]),
   .I3(InputBits[355]),
   .I4(InputBits[419]),
   .I5(InputBits[512])
);
LUT6 #(
   .INIT(64'b0000010100000101000001010000111100000000000000001000111100000101)  
) LUT6_414 (
   .O(gates_414),
   .I0(InputBits[483]),
   .I1(InputBits[154]),
   .I2(InputBits[482]),
   .I3(InputBits[499]),
   .I4(InputBits[127]),
   .I5(InputBits[339])
);
LUT6 #(
   .INIT(64'b0000000001110101000001110110011100000000000000110000000100011111)  
) LUT6_415 (
   .O(gates_415),
   .I0(InputBits[255]),
   .I1(InputBits[354]),
   .I2(InputBits[533]),
   .I3(InputBits[81]),
   .I4(InputBits[230]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000110011000000000010000000000000000100110)  
) LUT6_416 (
   .O(gates_416),
   .I0(InputBits[455]),
   .I1(InputBits[165]),
   .I2(InputBits[87]),
   .I3(InputBits[146]),
   .I4(InputBits[362]),
   .I5(InputBits[466])
);
LUT6 #(
   .INIT(64'b0100001000000000010101000101011000001000000100001101101001011111)  
) LUT6_417 (
   .O(gates_417),
   .I0(InputBits[360]),
   .I1(InputBits[156]),
   .I2(InputBits[213]),
   .I3(InputBits[133]),
   .I4(InputBits[78]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b0001000101010001000101111111011100000001000000010001011100000000)  
) LUT6_418 (
   .O(gates_418),
   .I0(InputBits[535]),
   .I1(InputBits[510]),
   .I2(InputBits[468]),
   .I3(InputBits[324]),
   .I4(InputBits[376]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100110011000100110011011110010111)  
) LUT6_419 (
   .O(gates_419),
   .I0(InputBits[536]),
   .I1(InputBits[194]),
   .I2(InputBits[130]),
   .I3(InputBits[357]),
   .I4(InputBits[459]),
   .I5(InputBits[255])
);
LUT6 #(
   .INIT(64'b0001000100010001010000000100010000010001000100010100010001001100)  
) LUT6_420 (
   .O(gates_420),
   .I0(InputBits[123]),
   .I1(InputBits[245]),
   .I2(InputBits[468]),
   .I3(InputBits[58]),
   .I4(InputBits[384]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000101010100000000000000000000010100001000)  
) LUT6_421 (
   .O(gates_421),
   .I0(InputBits[31]),
   .I1(InputBits[233]),
   .I2(InputBits[561]),
   .I3(InputBits[45]),
   .I4(InputBits[1]),
   .I5(InputBits[246])
);
LUT6 #(
   .INIT(64'b0000000000000011000000110011011100000000000000100000001100110010)  
) LUT6_422 (
   .O(gates_422),
   .I0(InputBits[325]),
   .I1(InputBits[409]),
   .I2(InputBits[69]),
   .I3(InputBits[8]),
   .I4(InputBits[569]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000000000010101000000111111000000000000000101010000010101110101)  
) LUT6_423 (
   .O(gates_423),
   .I0(InputBits[56]),
   .I1(InputBits[89]),
   .I2(InputBits[316]),
   .I3(InputBits[11]),
   .I4(InputBits[70]),
   .I5(InputBits[299])
);
LUT6 #(
   .INIT(64'b0000000000000001001100110011001100000001000000000011000000100010)  
) LUT6_424 (
   .O(gates_424),
   .I0(InputBits[166]),
   .I1(InputBits[74]),
   .I2(InputBits[308]),
   .I3(InputBits[114]),
   .I4(InputBits[290]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b0010001100100000001100110010001110110011001000111111111110100001)  
) LUT6_425 (
   .O(gates_425),
   .I0(InputBits[332]),
   .I1(InputBits[128]),
   .I2(InputBits[376]),
   .I3(InputBits[295]),
   .I4(InputBits[539]),
   .I5(InputBits[537])
);
LUT6 #(
   .INIT(64'b1010011000100001011101110011011110111111011101110011011101110111)  
) LUT6_426 (
   .O(gates_426),
   .I0(InputBits[492]),
   .I1(InputBits[255]),
   .I2(InputBits[135]),
   .I3(InputBits[197]),
   .I4(InputBits[64]),
   .I5(InputBits[244])
);
LUT6 #(
   .INIT(64'b0000111100001111000001000010010000010111000001110001011000010110)  
) LUT6_427 (
   .O(gates_427),
   .I0(InputBits[357]),
   .I1(InputBits[431]),
   .I2(InputBits[549]),
   .I3(InputBits[350]),
   .I4(InputBits[420]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0000001000010010001100100011001100110011001100110010001100000010)  
) LUT6_428 (
   .O(gates_428),
   .I0(InputBits[259]),
   .I1(InputBits[21]),
   .I2(InputBits[207]),
   .I3(InputBits[272]),
   .I4(InputBits[315]),
   .I5(InputBits[524])
);
LUT6 #(
   .INIT(64'b1011111110111000111111111111111011110001101000001111000011110001)  
) LUT6_429 (
   .O(gates_429),
   .I0(InputBits[186]),
   .I1(InputBits[328]),
   .I2(InputBits[318]),
   .I3(InputBits[423]),
   .I4(InputBits[149]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0000000100000000000000000000000011110011111100111111111111110111)  
) LUT6_430 (
   .O(gates_430),
   .I0(InputBits[232]),
   .I1(InputBits[493]),
   .I2(InputBits[261]),
   .I3(InputBits[180]),
   .I4(InputBits[448]),
   .I5(InputBits[409])
);
LUT6 #(
   .INIT(64'b0000000100000001000100010000010100000001000100000001000100000100)  
) LUT6_431 (
   .O(gates_431),
   .I0(InputBits[25]),
   .I1(InputBits[550]),
   .I2(InputBits[33]),
   .I3(InputBits[237]),
   .I4(InputBits[91]),
   .I5(InputBits[268])
);
LUT6 #(
   .INIT(64'b0101010101010001000000000001000101010100011101110000010001000111)  
) LUT6_432 (
   .O(gates_432),
   .I0(InputBits[16]),
   .I1(InputBits[153]),
   .I2(InputBits[413]),
   .I3(InputBits[129]),
   .I4(InputBits[389]),
   .I5(InputBits[150])
);
LUT6 #(
   .INIT(64'b0000000000000000000000111111010100000000000000011111001011111111)  
) LUT6_433 (
   .O(gates_433),
   .I0(InputBits[498]),
   .I1(InputBits[129]),
   .I2(InputBits[282]),
   .I3(InputBits[483]),
   .I4(InputBits[229]),
   .I5(InputBits[355])
);
LUT6 #(
   .INIT(64'b0000000000000001010001010101011100000000000000001111010001111111)  
) LUT6_434 (
   .O(gates_434),
   .I0(InputBits[101]),
   .I1(InputBits[452]),
   .I2(InputBits[65]),
   .I3(InputBits[103]),
   .I4(InputBits[565]),
   .I5(InputBits[333])
);
LUT6 #(
   .INIT(64'b0000000000000001010100000000000100000000000001010001000000000001)  
) LUT6_435 (
   .O(gates_435),
   .I0(InputBits[22]),
   .I1(InputBits[541]),
   .I2(InputBits[549]),
   .I3(InputBits[549]),
   .I4(InputBits[363]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000011100000000000001011)  
) LUT6_436 (
   .O(gates_436),
   .I0(InputBits[167]),
   .I1(InputBits[144]),
   .I2(InputBits[73]),
   .I3(InputBits[76]),
   .I4(InputBits[489]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b0000011101011111000000000001111100000010010111110000000010000010)  
) LUT6_437 (
   .O(gates_437),
   .I0(InputBits[525]),
   .I1(InputBits[405]),
   .I2(InputBits[459]),
   .I3(InputBits[99]),
   .I4(InputBits[370]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b0100010000000000000000000100010000000100000000000000000001001100)  
) LUT6_438 (
   .O(gates_438),
   .I0(InputBits[242]),
   .I1(InputBits[269]),
   .I2(InputBits[152]),
   .I3(InputBits[226]),
   .I4(InputBits[226]),
   .I5(InputBits[468])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001000100000000000000100010111011111111101)  
) LUT6_439 (
   .O(gates_439),
   .I0(InputBits[135]),
   .I1(InputBits[358]),
   .I2(InputBits[234]),
   .I3(InputBits[45]),
   .I4(InputBits[16]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0001000100010101000100010101010100010001000000000011000100010110)  
) LUT6_440 (
   .O(gates_440),
   .I0(InputBits[6]),
   .I1(InputBits[196]),
   .I2(InputBits[380]),
   .I3(InputBits[432]),
   .I4(InputBits[302]),
   .I5(InputBits[349])
);
LUT6 #(
   .INIT(64'b0001000101010111000100011101010000010001010101010001000101000100)  
) LUT6_441 (
   .O(gates_441),
   .I0(InputBits[537]),
   .I1(InputBits[291]),
   .I2(InputBits[160]),
   .I3(InputBits[478]),
   .I4(InputBits[373]),
   .I5(InputBits[211])
);
LUT6 #(
   .INIT(64'b0000010100100011000001000000101100000101101010110000010110111111)  
) LUT6_442 (
   .O(gates_442),
   .I0(InputBits[286]),
   .I1(InputBits[276]),
   .I2(InputBits[509]),
   .I3(InputBits[456]),
   .I4(InputBits[448]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b0000001000000010101100110011001100000011000000100011000000110010)  
) LUT6_443 (
   .O(gates_443),
   .I0(InputBits[442]),
   .I1(InputBits[228]),
   .I2(InputBits[222]),
   .I3(InputBits[400]),
   .I4(InputBits[36]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0001000100000000000100010011001100010001000100000001111100010001)  
) LUT6_444 (
   .O(gates_444),
   .I0(InputBits[298]),
   .I1(InputBits[99]),
   .I2(InputBits[445]),
   .I3(InputBits[244]),
   .I4(InputBits[81]),
   .I5(InputBits[179])
);
LUT6 #(
   .INIT(64'b0000001100000011001100110010001101010011000000000011011100100010)  
) LUT6_445 (
   .O(gates_445),
   .I0(InputBits[248]),
   .I1(InputBits[29]),
   .I2(InputBits[460]),
   .I3(InputBits[397]),
   .I4(InputBits[55]),
   .I5(InputBits[198])
);
LUT6 #(
   .INIT(64'b0000001100011010000000000100101000000001000110100000000101111010)  
) LUT6_446 (
   .O(gates_446),
   .I0(InputBits[262]),
   .I1(InputBits[520]),
   .I2(InputBits[68]),
   .I3(InputBits[431]),
   .I4(InputBits[161]),
   .I5(InputBits[186])
);
LUT6 #(
   .INIT(64'b0000001100000001000000110000011100000000000000010000001000001111)  
) LUT6_447 (
   .O(gates_447),
   .I0(InputBits[496]),
   .I1(InputBits[205]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[124]),
   .I5(InputBits[473])
);
LUT6 #(
   .INIT(64'b0000000000000000001110100010111100110011001100111010111010101110)  
) LUT6_448 (
   .O(gates_448),
   .I0(InputBits[373]),
   .I1(InputBits[364]),
   .I2(InputBits[208]),
   .I3(InputBits[440]),
   .I4(InputBits[384]),
   .I5(InputBits[94])
);
LUT6 #(
   .INIT(64'b0000100100000000001011010000000000001000000001000000110000001101)  
) LUT6_449 (
   .O(gates_449),
   .I0(InputBits[305]),
   .I1(InputBits[333]),
   .I2(InputBits[52]),
   .I3(InputBits[400]),
   .I4(InputBits[541]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010101111111011110001100001010001)  
) LUT6_450 (
   .O(gates_450),
   .I0(InputBits[111]),
   .I1(InputBits[424]),
   .I2(InputBits[154]),
   .I3(InputBits[502]),
   .I4(InputBits[501]),
   .I5(InputBits[457])
);
LUT6 #(
   .INIT(64'b0000000000100100000100110011000100000000000000000001011100010001)  
) LUT6_451 (
   .O(gates_451),
   .I0(InputBits[472]),
   .I1(InputBits[77]),
   .I2(InputBits[70]),
   .I3(InputBits[179]),
   .I4(InputBits[126]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0111011101111111111100110110111111010111011101110100010000000101)  
) LUT6_452 (
   .O(gates_452),
   .I0(InputBits[227]),
   .I1(InputBits[40]),
   .I2(InputBits[110]),
   .I3(InputBits[405]),
   .I4(InputBits[394]),
   .I5(InputBits[164])
);
LUT6 #(
   .INIT(64'b0010000100100101101100001010000000000101001101111011101011111011)  
) LUT6_453 (
   .O(gates_453),
   .I0(InputBits[271]),
   .I1(InputBits[331]),
   .I2(InputBits[200]),
   .I3(InputBits[462]),
   .I4(InputBits[384]),
   .I5(InputBits[82])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011110011111100011111110011110011)  
) LUT6_454 (
   .O(gates_454),
   .I0(InputBits[153]),
   .I1(InputBits[475]),
   .I2(InputBits[316]),
   .I3(InputBits[112]),
   .I4(InputBits[521]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000000100000000000100010000011000000000000000000001011100010111)  
) LUT6_455 (
   .O(gates_455),
   .I0(InputBits[46]),
   .I1(InputBits[192]),
   .I2(InputBits[58]),
   .I3(InputBits[372]),
   .I4(InputBits[433]),
   .I5(InputBits[229])
);
LUT6 #(
   .INIT(64'b0101111101011111110100110100111101110111010111110101001001010110)  
) LUT6_456 (
   .O(gates_456),
   .I0(InputBits[214]),
   .I1(InputBits[324]),
   .I2(InputBits[478]),
   .I3(InputBits[107]),
   .I4(InputBits[367]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b0000000001010000000000000101000001010000010100000101010001010100)  
) LUT6_457 (
   .O(gates_457),
   .I0(InputBits[575]),
   .I1(InputBits[222]),
   .I2(InputBits[341]),
   .I3(InputBits[382]),
   .I4(InputBits[499]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1111111100000111111111110001000000110111000111011111010101010000)  
) LUT6_458 (
   .O(gates_458),
   .I0(InputBits[520]),
   .I1(InputBits[462]),
   .I2(InputBits[268]),
   .I3(InputBits[317]),
   .I4(InputBits[368]),
   .I5(InputBits[176])
);
LUT6 #(
   .INIT(64'b0011001100010001001100110011001100010011000001010011001100110011)  
) LUT6_459 (
   .O(gates_459),
   .I0(InputBits[411]),
   .I1(InputBits[122]),
   .I2(InputBits[228]),
   .I3(InputBits[316]),
   .I4(InputBits[448]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000100000000101000001010100010100000111)  
) LUT6_460 (
   .O(gates_460),
   .I0(InputBits[504]),
   .I1(InputBits[468]),
   .I2(InputBits[561]),
   .I3(InputBits[203]),
   .I4(InputBits[356]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0101010101001111010101010101010101011101010001000101110101011101)  
) LUT6_461 (
   .O(gates_461),
   .I0(InputBits[101]),
   .I1(InputBits[284]),
   .I2(InputBits[227]),
   .I3(InputBits[238]),
   .I4(InputBits[109]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b0011001000110011001100100011101000110011101100110011001010111010)  
) LUT6_462 (
   .O(gates_462),
   .I0(InputBits[373]),
   .I1(InputBits[96]),
   .I2(InputBits[343]),
   .I3(InputBits[91]),
   .I4(InputBits[293]),
   .I5(InputBits[208])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000001000000000000000000000101000001110000)  
) LUT6_463 (
   .O(gates_463),
   .I0(InputBits[75]),
   .I1(InputBits[45]),
   .I2(InputBits[319]),
   .I3(InputBits[157]),
   .I4(InputBits[79]),
   .I5(InputBits[152])
);
LUT6 #(
   .INIT(64'b0000010011101110010000001110011000000100111011100000010111111110)  
) LUT6_464 (
   .O(gates_464),
   .I0(InputBits[268]),
   .I1(InputBits[418]),
   .I2(InputBits[114]),
   .I3(InputBits[384]),
   .I4(InputBits[209]),
   .I5(InputBits[88])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010101010101010101001100010101011101011111)  
) LUT6_465 (
   .O(gates_465),
   .I0(InputBits[515]),
   .I1(InputBits[462]),
   .I2(InputBits[129]),
   .I3(InputBits[184]),
   .I4(InputBits[360]),
   .I5(InputBits[520])
);
LUT6 #(
   .INIT(64'b0000000000000000000010100101001100000010110000010011111100010011)  
) LUT6_466 (
   .O(gates_466),
   .I0(InputBits[354]),
   .I1(InputBits[276]),
   .I2(InputBits[277]),
   .I3(InputBits[190]),
   .I4(InputBits[240]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0111000001111011000000000000010010111111111111110111011110001101)  
) LUT6_467 (
   .O(gates_467),
   .I0(InputBits[322]),
   .I1(InputBits[248]),
   .I2(InputBits[280]),
   .I3(InputBits[407]),
   .I4(InputBits[393]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0011000100110011000100000000000101010000001101110000000000000001)  
) LUT6_468 (
   .O(gates_468),
   .I0(InputBits[540]),
   .I1(InputBits[77]),
   .I2(InputBits[462]),
   .I3(InputBits[511]),
   .I4(InputBits[189]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0000000000000101000011111111111100000000000001000000000000110101)  
) LUT6_469 (
   .O(gates_469),
   .I0(InputBits[133]),
   .I1(InputBits[258]),
   .I2(InputBits[363]),
   .I3(InputBits[59]),
   .I4(InputBits[545]),
   .I5(InputBits[199])
);
LUT6 #(
   .INIT(64'b0000000000000100000101010001010000000100000100000000010100010000)  
) LUT6_470 (
   .O(gates_470),
   .I0(InputBits[22]),
   .I1(InputBits[36]),
   .I2(InputBits[267]),
   .I3(InputBits[501]),
   .I4(InputBits[156]),
   .I5(InputBits[321])
);
LUT6 #(
   .INIT(64'b0000000000000101000001010001101100000000000001010000011111111011)  
) LUT6_471 (
   .O(gates_471),
   .I0(InputBits[477]),
   .I1(InputBits[304]),
   .I2(InputBits[31]),
   .I3(InputBits[13]),
   .I4(InputBits[45]),
   .I5(InputBits[388])
);
LUT6 #(
   .INIT(64'b0101010101000000010111110101110101010101000100000101110100010101)  
) LUT6_472 (
   .O(gates_472),
   .I0(InputBits[508]),
   .I1(InputBits[464]),
   .I2(InputBits[291]),
   .I3(InputBits[212]),
   .I4(InputBits[515]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0000010100000000010101010000000100010101000100010001010100000001)  
) LUT6_473 (
   .O(gates_473),
   .I0(InputBits[97]),
   .I1(InputBits[514]),
   .I2(InputBits[149]),
   .I3(InputBits[394]),
   .I4(InputBits[331]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0011001110110000111100000111000000110011111100000111001111110000)  
) LUT6_474 (
   .O(gates_474),
   .I0(InputBits[161]),
   .I1(InputBits[540]),
   .I2(InputBits[342]),
   .I3(InputBits[347]),
   .I4(InputBits[440]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b0000000100010100001111111111111000000000000000100010000010111100)  
) LUT6_475 (
   .O(gates_475),
   .I0(InputBits[90]),
   .I1(InputBits[324]),
   .I2(InputBits[175]),
   .I3(InputBits[437]),
   .I4(InputBits[240]),
   .I5(InputBits[333])
);
LUT6 #(
   .INIT(64'b0101010001010100011101010101010101010101010101010101010100010011)  
) LUT6_476 (
   .O(gates_476),
   .I0(InputBits[218]),
   .I1(InputBits[105]),
   .I2(InputBits[185]),
   .I3(InputBits[421]),
   .I4(InputBits[479]),
   .I5(InputBits[201])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000100011100000000000100010000000001000111)  
) LUT6_477 (
   .O(gates_477),
   .I0(InputBits[29]),
   .I1(InputBits[67]),
   .I2(InputBits[228]),
   .I3(InputBits[97]),
   .I4(InputBits[12]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0101010101010101000000000000010001010101010101010100101001011010)  
) LUT6_478 (
   .O(gates_478),
   .I0(InputBits[479]),
   .I1(InputBits[399]),
   .I2(InputBits[263]),
   .I3(InputBits[463]),
   .I4(InputBits[238]),
   .I5(InputBits[226])
);
LUT6 #(
   .INIT(64'b1111001101110000111111111111001111111111011100111111111101110111)  
) LUT6_479 (
   .O(gates_479),
   .I0(InputBits[109]),
   .I1(InputBits[253]),
   .I2(InputBits[367]),
   .I3(InputBits[373]),
   .I4(InputBits[250]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0000000000110001000000000001000100000000011100010000000000110001)  
) LUT6_480 (
   .O(gates_480),
   .I0(InputBits[514]),
   .I1(InputBits[458]),
   .I2(InputBits[271]),
   .I3(InputBits[74]),
   .I4(InputBits[159]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000010101011100000001010101111)  
) LUT6_481 (
   .O(gates_481),
   .I0(InputBits[236]),
   .I1(InputBits[31]),
   .I2(InputBits[380]),
   .I3(InputBits[557]),
   .I4(InputBits[299]),
   .I5(InputBits[562])
);
LUT6 #(
   .INIT(64'b0000000000001100000010110000100000000001000011100000111110001000)  
) LUT6_482 (
   .O(gates_482),
   .I0(InputBits[417]),
   .I1(InputBits[346]),
   .I2(InputBits[386]),
   .I3(InputBits[238]),
   .I4(InputBits[431]),
   .I5(InputBits[56])
);
LUT6 #(
   .INIT(64'b0000101000001011000010110000111100001000000010100000100000001111)  
) LUT6_483 (
   .O(gates_483),
   .I0(InputBits[442]),
   .I1(InputBits[321]),
   .I2(InputBits[26]),
   .I3(InputBits[402]),
   .I4(InputBits[475]),
   .I5(InputBits[155])
);
LUT6 #(
   .INIT(64'b1100110011011111101111111011111100001110001011110000111100011111)  
) LUT6_484 (
   .O(gates_484),
   .I0(InputBits[436]),
   .I1(InputBits[449]),
   .I2(InputBits[230]),
   .I3(InputBits[273]),
   .I4(InputBits[427]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001010101000100010011010000110111)  
) LUT6_485 (
   .O(gates_485),
   .I0(InputBits[497]),
   .I1(InputBits[12]),
   .I2(InputBits[477]),
   .I3(InputBits[426]),
   .I4(InputBits[157]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0000000001000001000000000101010100000000010101010000001000011010)  
) LUT6_486 (
   .O(gates_486),
   .I0(InputBits[236]),
   .I1(InputBits[231]),
   .I2(InputBits[232]),
   .I3(InputBits[565]),
   .I4(InputBits[384]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000001100000011000000100000000000000011000101110000001100010011)  
) LUT6_487 (
   .O(gates_487),
   .I0(InputBits[179]),
   .I1(InputBits[266]),
   .I2(InputBits[71]),
   .I3(InputBits[437]),
   .I4(InputBits[346]),
   .I5(InputBits[229])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010001000101010000010100000101010001110110)  
) LUT6_488 (
   .O(gates_488),
   .I0(InputBits[360]),
   .I1(InputBits[453]),
   .I2(InputBits[368]),
   .I3(InputBits[235]),
   .I4(InputBits[498]),
   .I5(InputBits[215])
);
LUT6 #(
   .INIT(64'b0000000011110000000000000001010000000000011100010000010101110101)  
) LUT6_489 (
   .O(gates_489),
   .I0(InputBits[535]),
   .I1(InputBits[302]),
   .I2(InputBits[262]),
   .I3(InputBits[290]),
   .I4(InputBits[462]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b0000000010010000000100000000000000000000111110110001110100000011)  
) LUT6_490 (
   .O(gates_490),
   .I0(InputBits[380]),
   .I1(InputBits[403]),
   .I2(InputBits[134]),
   .I3(InputBits[523]),
   .I4(InputBits[239]),
   .I5(InputBits[508])
);
LUT6 #(
   .INIT(64'b0010001000110011001000100011001100110011001100110000101000100010)  
) LUT6_491 (
   .O(gates_491),
   .I0(InputBits[398]),
   .I1(InputBits[566]),
   .I2(InputBits[406]),
   .I3(InputBits[250]),
   .I4(InputBits[390]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0000111100001000000011110000100000001111000001010000111100001001)  
) LUT6_492 (
   .O(gates_492),
   .I0(InputBits[475]),
   .I1(InputBits[423]),
   .I2(InputBits[217]),
   .I3(InputBits[366]),
   .I4(InputBits[204]),
   .I5(InputBits[376])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000011011100000000000010100010000000101010)  
) LUT6_493 (
   .O(gates_493),
   .I0(InputBits[420]),
   .I1(InputBits[486]),
   .I2(InputBits[444]),
   .I3(InputBits[543]),
   .I4(InputBits[461]),
   .I5(InputBits[119])
);
LUT6 #(
   .INIT(64'b0000000001010100000001010100010100000000000101010000010101010100)  
) LUT6_494 (
   .O(gates_494),
   .I0(InputBits[361]),
   .I1(InputBits[258]),
   .I2(InputBits[37]),
   .I3(InputBits[94]),
   .I4(InputBits[15]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0000000000000000000101110000000100000000000000000001001100000001)  
) LUT6_495 (
   .O(gates_495),
   .I0(InputBits[510]),
   .I1(InputBits[458]),
   .I2(InputBits[148]),
   .I3(InputBits[66]),
   .I4(InputBits[576]),
   .I5(InputBits[303])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000000011100000010000000110001000100010001)  
) LUT6_496 (
   .O(gates_496),
   .I0(InputBits[232]),
   .I1(InputBits[148]),
   .I2(InputBits[43]),
   .I3(InputBits[205]),
   .I4(InputBits[568]),
   .I5(InputBits[197])
);
LUT6 #(
   .INIT(64'b0000000000000111000000000000011100000010000100010000000000111111)  
) LUT6_497 (
   .O(gates_497),
   .I0(InputBits[85]),
   .I1(InputBits[496]),
   .I2(InputBits[276]),
   .I3(InputBits[504]),
   .I4(InputBits[231]),
   .I5(InputBits[299])
);
LUT6 #(
   .INIT(64'b0000101100001000000111110000101000000010000011000011111100001110)  
) LUT6_498 (
   .O(gates_498),
   .I0(InputBits[398]),
   .I1(InputBits[477]),
   .I2(InputBits[314]),
   .I3(InputBits[318]),
   .I4(InputBits[510]),
   .I5(InputBits[132])
);
LUT6 #(
   .INIT(64'b0000000000001000000000000000000000000000000010100000000011111010)  
) LUT6_499 (
   .O(gates_499),
   .I0(InputBits[224]),
   .I1(InputBits[352]),
   .I2(InputBits[407]),
   .I3(InputBits[530]),
   .I4(InputBits[141]),
   .I5(InputBits[557])
);
LUT6 #(
   .INIT(64'b1010111100101010000000000000000000000000000000001111111010101110)  
) LUT6_500 (
   .O(gates_500),
   .I0(InputBits[419]),
   .I1(InputBits[469]),
   .I2(InputBits[489]),
   .I3(InputBits[176]),
   .I4(InputBits[328]),
   .I5(InputBits[328])
);
LUT6 #(
   .INIT(64'b0000010100000101000011010000110110011100000101011100110101011101)  
) LUT6_501 (
   .O(gates_501),
   .I0(InputBits[514]),
   .I1(InputBits[393]),
   .I2(InputBits[540]),
   .I3(InputBits[131]),
   .I4(InputBits[387]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0000000000110011000000000011001100110011110111110011001101010101)  
) LUT6_502 (
   .O(gates_502),
   .I0(InputBits[490]),
   .I1(InputBits[477]),
   .I2(InputBits[154]),
   .I3(InputBits[167]),
   .I4(InputBits[347]),
   .I5(InputBits[69])
);
LUT6 #(
   .INIT(64'b0011000111110111000001000101000000000001110101110000000000000001)  
) LUT6_503 (
   .O(gates_503),
   .I0(InputBits[127]),
   .I1(InputBits[464]),
   .I2(InputBits[428]),
   .I3(InputBits[195]),
   .I4(InputBits[270]),
   .I5(InputBits[426])
);
LUT6 #(
   .INIT(64'b0000000100000000001100110011000000000001000000110011001100110001)  
) LUT6_504 (
   .O(gates_504),
   .I0(InputBits[107]),
   .I1(InputBits[50]),
   .I2(InputBits[291]),
   .I3(InputBits[394]),
   .I4(InputBits[120]),
   .I5(InputBits[448])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001001100000000000000010001000000110011)  
) LUT6_505 (
   .O(gates_505),
   .I0(InputBits[518]),
   .I1(InputBits[121]),
   .I2(InputBits[281]),
   .I3(InputBits[559]),
   .I4(InputBits[278]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0000000010000001110111010101110100000000001010000000110011101111)  
) LUT6_506 (
   .O(gates_506),
   .I0(InputBits[191]),
   .I1(InputBits[214]),
   .I2(InputBits[298]),
   .I3(InputBits[128]),
   .I4(InputBits[192]),
   .I5(InputBits[245])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000111011100000001011101110101000101110101)  
) LUT6_507 (
   .O(gates_507),
   .I0(InputBits[535]),
   .I1(InputBits[501]),
   .I2(InputBits[442]),
   .I3(InputBits[70]),
   .I4(InputBits[244]),
   .I5(InputBits[286])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101000000010000010100010101)  
) LUT6_508 (
   .O(gates_508),
   .I0(InputBits[49]),
   .I1(InputBits[492]),
   .I2(InputBits[52]),
   .I3(InputBits[336]),
   .I4(InputBits[280]),
   .I5(InputBits[552])
);
LUT6 #(
   .INIT(64'b0000010000000101000011010000010000001011000000110000011100000001)  
) LUT6_509 (
   .O(gates_509),
   .I0(InputBits[429]),
   .I1(InputBits[328]),
   .I2(InputBits[73]),
   .I3(InputBits[326]),
   .I4(InputBits[136]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0000111100111111000000000011001100011111000111110001000100111011)  
) LUT6_510 (
   .O(gates_510),
   .I0(InputBits[157]),
   .I1(InputBits[492]),
   .I2(InputBits[300]),
   .I3(InputBits[543]),
   .I4(InputBits[213]),
   .I5(InputBits[427])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010000101101000011111111111110110)  
) LUT6_511 (
   .O(gates_511),
   .I0(InputBits[189]),
   .I1(InputBits[324]),
   .I2(InputBits[118]),
   .I3(InputBits[345]),
   .I4(InputBits[45]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000100001000000010111)  
) LUT6_512 (
   .O(gates_512),
   .I0(InputBits[136]),
   .I1(InputBits[273]),
   .I2(InputBits[469]),
   .I3(InputBits[151]),
   .I4(InputBits[52]),
   .I5(InputBits[554])
);
LUT6 #(
   .INIT(64'b0000000100000001000101111001000100000000000000000000010110110001)  
) LUT6_513 (
   .O(gates_513),
   .I0(InputBits[434]),
   .I1(InputBits[299]),
   .I2(InputBits[43]),
   .I3(InputBits[222]),
   .I4(InputBits[51]),
   .I5(InputBits[138])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100000001100000000000100110001)  
) LUT6_514 (
   .O(gates_514),
   .I0(InputBits[173]),
   .I1(InputBits[74]),
   .I2(InputBits[423]),
   .I3(InputBits[510]),
   .I4(InputBits[111]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000001010100000000010101000001000011111110)  
) LUT6_515 (
   .O(gates_515),
   .I0(InputBits[244]),
   .I1(InputBits[222]),
   .I2(InputBits[416]),
   .I3(InputBits[533]),
   .I4(InputBits[37]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010101010000000000000100010001000101010101)  
) LUT6_516 (
   .O(gates_516),
   .I0(InputBits[2]),
   .I1(InputBits[455]),
   .I2(InputBits[524]),
   .I3(InputBits[213]),
   .I4(InputBits[550]),
   .I5(InputBits[486])
);
LUT6 #(
   .INIT(64'b0000000000000000001111000000100000000000000100001111111111110010)  
) LUT6_517 (
   .O(gates_517),
   .I0(InputBits[341]),
   .I1(InputBits[378]),
   .I2(InputBits[393]),
   .I3(InputBits[318]),
   .I4(InputBits[481]),
   .I5(InputBits[362])
);
LUT6 #(
   .INIT(64'b0011100010100000001011111010101000011001001000001011111111111010)  
) LUT6_518 (
   .O(gates_518),
   .I0(InputBits[294]),
   .I1(InputBits[332]),
   .I2(InputBits[547]),
   .I3(InputBits[395]),
   .I4(InputBits[100]),
   .I5(InputBits[297])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001100001001100001110)  
) LUT6_519 (
   .O(gates_519),
   .I0(InputBits[272]),
   .I1(InputBits[45]),
   .I2(InputBits[451]),
   .I3(InputBits[312]),
   .I4(InputBits[282]),
   .I5(InputBits[150])
);
LUT6 #(
   .INIT(64'b0000000000110011000000000011000000010000111101110001000000000000)  
) LUT6_520 (
   .O(gates_520),
   .I0(InputBits[356]),
   .I1(InputBits[535]),
   .I2(InputBits[249]),
   .I3(InputBits[565]),
   .I4(InputBits[395]),
   .I5(InputBits[67])
);
LUT6 #(
   .INIT(64'b0000001000111111000000110011111100000010001011110000001100001010)  
) LUT6_521 (
   .O(gates_521),
   .I0(InputBits[296]),
   .I1(InputBits[243]),
   .I2(InputBits[512]),
   .I3(InputBits[13]),
   .I4(InputBits[212]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0011000000010000001100111011001100110110001100000011111111111011)  
) LUT6_522 (
   .O(gates_522),
   .I0(InputBits[245]),
   .I1(InputBits[565]),
   .I2(InputBits[310]),
   .I3(InputBits[235]),
   .I4(InputBits[252]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000000000000000000001000000010)  
) LUT6_523 (
   .O(gates_523),
   .I0(InputBits[395]),
   .I1(InputBits[553]),
   .I2(InputBits[22]),
   .I3(InputBits[154]),
   .I4(InputBits[555]),
   .I5(InputBits[409])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100000011001100110011)  
) LUT6_524 (
   .O(gates_524),
   .I0(InputBits[378]),
   .I1(InputBits[575]),
   .I2(InputBits[69]),
   .I3(InputBits[156]),
   .I4(InputBits[276]),
   .I5(InputBits[529])
);
LUT6 #(
   .INIT(64'b0101010100010101000101010001010100000101000000000000010100010011)  
) LUT6_525 (
   .O(gates_525),
   .I0(InputBits[531]),
   .I1(InputBits[81]),
   .I2(InputBits[278]),
   .I3(InputBits[162]),
   .I4(InputBits[126]),
   .I5(InputBits[244])
);
LUT6 #(
   .INIT(64'b0000000100000001000001010000010100000000000000000000010000000101)  
) LUT6_526 (
   .O(gates_526),
   .I0(InputBits[22]),
   .I1(InputBits[15]),
   .I2(InputBits[560]),
   .I3(InputBits[328]),
   .I4(InputBits[174]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0100000000000000000000100000001100010010000101100000001100000011)  
) LUT6_527 (
   .O(gates_527),
   .I0(InputBits[288]),
   .I1(InputBits[571]),
   .I2(InputBits[545]),
   .I3(InputBits[327]),
   .I4(InputBits[473]),
   .I5(InputBits[159])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011110111011100011111000000000000)  
) LUT6_528 (
   .O(gates_528),
   .I0(InputBits[511]),
   .I1(InputBits[209]),
   .I2(InputBits[200]),
   .I3(InputBits[295]),
   .I4(InputBits[421]),
   .I5(InputBits[27])
);
LUT6 #(
   .INIT(64'b0011000100010010111111111111001100010000000100001101010101010000)  
) LUT6_529 (
   .O(gates_529),
   .I0(InputBits[354]),
   .I1(InputBits[379]),
   .I2(InputBits[394]),
   .I3(InputBits[419]),
   .I4(InputBits[95]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0000110000000000000011000100100000011111000100011000111100011011)  
) LUT6_530 (
   .O(gates_530),
   .I0(InputBits[233]),
   .I1(InputBits[297]),
   .I2(InputBits[240]),
   .I3(InputBits[393]),
   .I4(InputBits[132]),
   .I5(InputBits[250])
);
LUT6 #(
   .INIT(64'b0000000101011111000100000101101100000000010101110000000010111010)  
) LUT6_531 (
   .O(gates_531),
   .I0(InputBits[548]),
   .I1(InputBits[207]),
   .I2(InputBits[422]),
   .I3(InputBits[483]),
   .I4(InputBits[334]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b0101010100000100000001000000010011111111111111110000010100000001)  
) LUT6_532 (
   .O(gates_532),
   .I0(InputBits[128]),
   .I1(InputBits[161]),
   .I2(InputBits[487]),
   .I3(InputBits[89]),
   .I4(InputBits[247]),
   .I5(InputBits[250])
);
LUT6 #(
   .INIT(64'b0011001100110111001100110011011100111011000111110011001100010101)  
) LUT6_533 (
   .O(gates_533),
   .I0(InputBits[83]),
   .I1(InputBits[77]),
   .I2(InputBits[519]),
   .I3(InputBits[286]),
   .I4(InputBits[414]),
   .I5(InputBits[268])
);
LUT6 #(
   .INIT(64'b0101010100000001000001010001010101010001000000000101010100000011)  
) LUT6_534 (
   .O(gates_534),
   .I0(InputBits[551]),
   .I1(InputBits[128]),
   .I2(InputBits[62]),
   .I3(InputBits[415]),
   .I4(InputBits[86]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010101111101111111010111111101111)  
) LUT6_535 (
   .O(gates_535),
   .I0(InputBits[236]),
   .I1(InputBits[308]),
   .I2(InputBits[492]),
   .I3(InputBits[464]),
   .I4(InputBits[182]),
   .I5(InputBits[217])
);
LUT6 #(
   .INIT(64'b0000000000000000000001110000001000000011000000010000001000001011)  
) LUT6_536 (
   .O(gates_536),
   .I0(InputBits[176]),
   .I1(InputBits[172]),
   .I2(InputBits[48]),
   .I3(InputBits[280]),
   .I4(InputBits[46]),
   .I5(InputBits[569])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000000001101)  
) LUT6_537 (
   .O(gates_537),
   .I0(InputBits[298]),
   .I1(InputBits[44]),
   .I2(InputBits[241]),
   .I3(InputBits[56]),
   .I4(InputBits[481]),
   .I5(InputBits[448])
);
LUT6 #(
   .INIT(64'b0100000000000000110100011100101111010101110101011111011111111111)  
) LUT6_538 (
   .O(gates_538),
   .I0(InputBits[207]),
   .I1(InputBits[132]),
   .I2(InputBits[383]),
   .I3(InputBits[161]),
   .I4(InputBits[517]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0101000100000000010101010001000101010011000010001111111100110011)  
) LUT6_539 (
   .O(gates_539),
   .I0(InputBits[15]),
   .I1(InputBits[109]),
   .I2(InputBits[186]),
   .I3(InputBits[366]),
   .I4(InputBits[228]),
   .I5(InputBits[153])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010001000000000001000000000001000100010011)  
) LUT6_540 (
   .O(gates_540),
   .I0(InputBits[572]),
   .I1(InputBits[3]),
   .I2(InputBits[436]),
   .I3(InputBits[526]),
   .I4(InputBits[255]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1000000000010000000000000010000000000101000001110000001100000111)  
) LUT6_541 (
   .O(gates_541),
   .I0(InputBits[243]),
   .I1(InputBits[489]),
   .I2(InputBits[519]),
   .I3(InputBits[86]),
   .I4(InputBits[248]),
   .I5(InputBits[519])
);
LUT6 #(
   .INIT(64'b0000110100001111000101110101111100000100000000000000010100000000)  
) LUT6_542 (
   .O(gates_542),
   .I0(InputBits[79]),
   .I1(InputBits[487]),
   .I2(InputBits[537]),
   .I3(InputBits[295]),
   .I4(InputBits[486]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100010001000101011001100110011)  
) LUT6_543 (
   .O(gates_543),
   .I0(InputBits[212]),
   .I1(InputBits[507]),
   .I2(InputBits[138]),
   .I3(InputBits[182]),
   .I4(InputBits[132]),
   .I5(InputBits[19])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001111001111110000001101100000)  
) LUT6_544 (
   .O(gates_544),
   .I0(InputBits[376]),
   .I1(InputBits[435]),
   .I2(InputBits[17]),
   .I3(InputBits[165]),
   .I4(InputBits[391]),
   .I5(InputBits[554])
);
LUT6 #(
   .INIT(64'b0000001000001011000000001001001100000000000000110000000000110111)  
) LUT6_545 (
   .O(gates_545),
   .I0(InputBits[134]),
   .I1(InputBits[518]),
   .I2(InputBits[76]),
   .I3(InputBits[482]),
   .I4(InputBits[404]),
   .I5(InputBits[88])
);
LUT6 #(
   .INIT(64'b0000111101000111000011110101111110001010000000000000111100000000)  
) LUT6_546 (
   .O(gates_546),
   .I0(InputBits[400]),
   .I1(InputBits[466]),
   .I2(InputBits[144]),
   .I3(InputBits[309]),
   .I4(InputBits[205]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0000000000000010000011010000111000000001000011110000110100001111)  
) LUT6_547 (
   .O(gates_547),
   .I0(InputBits[94]),
   .I1(InputBits[350]),
   .I2(InputBits[122]),
   .I3(InputBits[500]),
   .I4(InputBits[541]),
   .I5(InputBits[105])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010101010000000000000000000000010101010110)  
) LUT6_548 (
   .O(gates_548),
   .I0(InputBits[29]),
   .I1(InputBits[247]),
   .I2(InputBits[549]),
   .I3(InputBits[191]),
   .I4(InputBits[28]),
   .I5(InputBits[403])
);
LUT6 #(
   .INIT(64'b0000000001000001000000000101110100000101010001010101000001010101)  
) LUT6_549 (
   .O(gates_549),
   .I0(InputBits[28]),
   .I1(InputBits[87]),
   .I2(InputBits[548]),
   .I3(InputBits[514]),
   .I4(InputBits[249]),
   .I5(InputBits[305])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001111111011111110010011100010011)  
) LUT6_550 (
   .O(gates_550),
   .I0(InputBits[282]),
   .I1(InputBits[274]),
   .I2(InputBits[56]),
   .I3(InputBits[283]),
   .I4(InputBits[366]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010001011111010001010001111111)  
) LUT6_551 (
   .O(gates_551),
   .I0(InputBits[253]),
   .I1(InputBits[267]),
   .I2(InputBits[392]),
   .I3(InputBits[565]),
   .I4(InputBits[255]),
   .I5(InputBits[573])
);
LUT6 #(
   .INIT(64'b0000000000110010000000000011001000000011001100110001000101110111)  
) LUT6_552 (
   .O(gates_552),
   .I0(InputBits[131]),
   .I1(InputBits[126]),
   .I2(InputBits[324]),
   .I3(InputBits[536]),
   .I4(InputBits[437]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010000000100010001000100000001)  
) LUT6_553 (
   .O(gates_553),
   .I0(InputBits[506]),
   .I1(InputBits[533]),
   .I2(InputBits[353]),
   .I3(InputBits[120]),
   .I4(InputBits[175]),
   .I5(InputBits[565])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000000100010000000000000001010101010101)  
) LUT6_554 (
   .O(gates_554),
   .I0(InputBits[146]),
   .I1(InputBits[201]),
   .I2(InputBits[243]),
   .I3(InputBits[522]),
   .I4(InputBits[253]),
   .I5(InputBits[386])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010001000000000000000000100001000100110001)  
) LUT6_555 (
   .O(gates_555),
   .I0(InputBits[504]),
   .I1(InputBits[19]),
   .I2(InputBits[232]),
   .I3(InputBits[320]),
   .I4(InputBits[254]),
   .I5(InputBits[6])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000000000111010111110000000000000001)  
) LUT6_556 (
   .O(gates_556),
   .I0(InputBits[274]),
   .I1(InputBits[82]),
   .I2(InputBits[76]),
   .I3(InputBits[540]),
   .I4(InputBits[394]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000001001100110001001100110001001000100010)  
) LUT6_557 (
   .O(gates_557),
   .I0(InputBits[267]),
   .I1(InputBits[562]),
   .I2(InputBits[375]),
   .I3(InputBits[430]),
   .I4(InputBits[398]),
   .I5(InputBits[569])
);
LUT6 #(
   .INIT(64'b0011000000110010010101010110000000110011001100110110010001110110)  
) LUT6_558 (
   .O(gates_558),
   .I0(InputBits[202]),
   .I1(InputBits[13]),
   .I2(InputBits[113]),
   .I3(InputBits[87]),
   .I4(InputBits[309]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000100000001010100010000010111111101)  
) LUT6_559 (
   .O(gates_559),
   .I0(InputBits[450]),
   .I1(InputBits[358]),
   .I2(InputBits[292]),
   .I3(InputBits[240]),
   .I4(InputBits[143]),
   .I5(InputBits[51])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000100111111110111111101101100011111110)  
) LUT6_560 (
   .O(gates_560),
   .I0(InputBits[392]),
   .I1(InputBits[367]),
   .I2(InputBits[245]),
   .I3(InputBits[498]),
   .I4(InputBits[259]),
   .I5(InputBits[6])
);
LUT6 #(
   .INIT(64'b0100010001010101010101000101010100000100000011010001010000000100)  
) LUT6_561 (
   .O(gates_561),
   .I0(InputBits[507]),
   .I1(InputBits[165]),
   .I2(InputBits[233]),
   .I3(InputBits[118]),
   .I4(InputBits[284]),
   .I5(InputBits[293])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000010011010101000)  
) LUT6_562 (
   .O(gates_562),
   .I0(InputBits[321]),
   .I1(InputBits[43]),
   .I2(InputBits[38]),
   .I3(InputBits[248]),
   .I4(InputBits[576]),
   .I5(InputBits[170])
);
LUT6 #(
   .INIT(64'b0000000000000100001100001100010100000000000001010001111011011111)  
) LUT6_563 (
   .O(gates_563),
   .I0(InputBits[448]),
   .I1(InputBits[186]),
   .I2(InputBits[312]),
   .I3(InputBits[79]),
   .I4(InputBits[46]),
   .I5(InputBits[490])
);
LUT6 #(
   .INIT(64'b0010001000100010001110110010001000100010001000100011011100100010)  
) LUT6_564 (
   .O(gates_564),
   .I0(InputBits[341]),
   .I1(InputBits[30]),
   .I2(InputBits[151]),
   .I3(InputBits[443]),
   .I4(InputBits[470]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1000111111111111100011011111110010001110111111110000110011011100)  
) LUT6_565 (
   .O(gates_565),
   .I0(InputBits[450]),
   .I1(InputBits[396]),
   .I2(InputBits[427]),
   .I3(InputBits[498]),
   .I4(InputBits[319]),
   .I5(InputBits[398])
);
LUT6 #(
   .INIT(64'b0000111100001010010110100101111000001110000011110000101011011110)  
) LUT6_566 (
   .O(gates_566),
   .I0(InputBits[235]),
   .I1(InputBits[444]),
   .I2(InputBits[432]),
   .I3(InputBits[331]),
   .I4(InputBits[67]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0000010011010100000000001101010100000000010001000000000001110101)  
) LUT6_567 (
   .O(gates_567),
   .I0(InputBits[251]),
   .I1(InputBits[442]),
   .I2(InputBits[222]),
   .I3(InputBits[28]),
   .I4(InputBits[488]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000010100000010000110110000000000011011)  
) LUT6_568 (
   .O(gates_568),
   .I0(InputBits[188]),
   .I1(InputBits[496]),
   .I2(InputBits[10]),
   .I3(InputBits[28]),
   .I4(InputBits[322]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0000000100010000000000010000100000000000000100000000000100011111)  
) LUT6_569 (
   .O(gates_569),
   .I0(InputBits[363]),
   .I1(InputBits[458]),
   .I2(InputBits[143]),
   .I3(InputBits[8]),
   .I4(InputBits[279]),
   .I5(InputBits[231])
);
LUT6 #(
   .INIT(64'b0000000100000010000000010000001100000001000100110000000100000011)  
) LUT6_570 (
   .O(gates_570),
   .I0(InputBits[287]),
   .I1(InputBits[24]),
   .I2(InputBits[75]),
   .I3(InputBits[363]),
   .I4(InputBits[150]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001010101000000000000000000011101110101010)  
) LUT6_571 (
   .O(gates_571),
   .I0(InputBits[370]),
   .I1(InputBits[80]),
   .I2(InputBits[183]),
   .I3(InputBits[93]),
   .I4(InputBits[568]),
   .I5(InputBits[79])
);
LUT6 #(
   .INIT(64'b0010000000100010111111111010111001110111011001101111111111101111)  
) LUT6_572 (
   .O(gates_572),
   .I0(InputBits[370]),
   .I1(InputBits[270]),
   .I2(InputBits[402]),
   .I3(InputBits[367]),
   .I4(InputBits[508]),
   .I5(InputBits[105])
);
LUT6 #(
   .INIT(64'b0000100100000010000011010100101100001010000010101100111110001011)  
) LUT6_573 (
   .O(gates_573),
   .I0(InputBits[444]),
   .I1(InputBits[475]),
   .I2(InputBits[482]),
   .I3(InputBits[500]),
   .I4(InputBits[159]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0011000110110011000000000010000000111011101110110000001010001011)  
) LUT6_574 (
   .O(gates_574),
   .I0(InputBits[272]),
   .I1(InputBits[256]),
   .I2(InputBits[153]),
   .I3(InputBits[510]),
   .I4(InputBits[236]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0000000001000001000000000100111000000000010001100000000011101111)  
) LUT6_575 (
   .O(gates_575),
   .I0(InputBits[143]),
   .I1(InputBits[263]),
   .I2(InputBits[111]),
   .I3(InputBits[55]),
   .I4(InputBits[475]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1110011100110011110111111111111100000000001100110000000000100011)  
) LUT6_576 (
   .O(gates_576),
   .I0(InputBits[114]),
   .I1(InputBits[232]),
   .I2(InputBits[128]),
   .I3(InputBits[279]),
   .I4(InputBits[387]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000000100010001010101010100010100010000000100010001010101000111)  
) LUT6_577 (
   .O(gates_577),
   .I0(InputBits[17]),
   .I1(InputBits[116]),
   .I2(InputBits[227]),
   .I3(InputBits[221]),
   .I4(InputBits[384]),
   .I5(InputBits[159])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000111111110010011000000011)  
) LUT6_578 (
   .O(gates_578),
   .I0(InputBits[322]),
   .I1(InputBits[173]),
   .I2(InputBits[492]),
   .I3(InputBits[290]),
   .I4(InputBits[213]),
   .I5(InputBits[574])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000101000000011000000000000111101011011)  
) LUT6_579 (
   .O(gates_579),
   .I0(InputBits[429]),
   .I1(InputBits[411]),
   .I2(InputBits[46]),
   .I3(InputBits[502]),
   .I4(InputBits[100]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0000000011010101000100110101010100000000110011000001001101011111)  
) LUT6_580 (
   .O(gates_580),
   .I0(InputBits[131]),
   .I1(InputBits[92]),
   .I2(InputBits[137]),
   .I3(InputBits[12]),
   .I4(InputBits[521]),
   .I5(InputBits[161])
);
LUT6 #(
   .INIT(64'b0000000100000000000000110000001000000111000000000000111100001111)  
) LUT6_581 (
   .O(gates_581),
   .I0(InputBits[467]),
   .I1(InputBits[160]),
   .I2(InputBits[553]),
   .I3(InputBits[375]),
   .I4(InputBits[484]),
   .I5(InputBits[109])
);
LUT6 #(
   .INIT(64'b0011110100001101000001010000110000011101000011000001010100001100)  
) LUT6_582 (
   .O(gates_582),
   .I0(InputBits[250]),
   .I1(InputBits[239]),
   .I2(InputBits[411]),
   .I3(InputBits[417]),
   .I4(InputBits[439]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000000000000000000000001001100110011)  
) LUT6_583 (
   .O(gates_583),
   .I0(InputBits[56]),
   .I1(InputBits[194]),
   .I2(InputBits[473]),
   .I3(InputBits[305]),
   .I4(InputBits[275]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000100000000000000000001001000010011)  
) LUT6_584 (
   .O(gates_584),
   .I0(InputBits[336]),
   .I1(InputBits[531]),
   .I2(InputBits[339]),
   .I3(InputBits[427]),
   .I4(InputBits[481]),
   .I5(InputBits[215])
);
LUT6 #(
   .INIT(64'b0010110000111100100111101011111001110100011111001111110011111100)  
) LUT6_585 (
   .O(gates_585),
   .I0(InputBits[113]),
   .I1(InputBits[396]),
   .I2(InputBits[340]),
   .I3(InputBits[83]),
   .I4(InputBits[495]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000100000101000001000000010100010110)  
) LUT6_586 (
   .O(gates_586),
   .I0(InputBits[545]),
   .I1(InputBits[11]),
   .I2(InputBits[567]),
   .I3(InputBits[430]),
   .I4(InputBits[159]),
   .I5(InputBits[215])
);
LUT6 #(
   .INIT(64'b0000011111010011000000001111001011100111111110111110001010111010)  
) LUT6_587 (
   .O(gates_587),
   .I0(InputBits[261]),
   .I1(InputBits[175]),
   .I2(InputBits[222]),
   .I3(InputBits[485]),
   .I4(InputBits[366]),
   .I5(InputBits[281])
);
LUT6 #(
   .INIT(64'b0000110101011111010011110101111100000100110101010000000011000011)  
) LUT6_588 (
   .O(gates_588),
   .I0(InputBits[492]),
   .I1(InputBits[109]),
   .I2(InputBits[503]),
   .I3(InputBits[460]),
   .I4(InputBits[61]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100110001001101010001)  
) LUT6_589 (
   .O(gates_589),
   .I0(InputBits[489]),
   .I1(InputBits[76]),
   .I2(InputBits[461]),
   .I3(InputBits[288]),
   .I4(InputBits[94]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0000000001011101000000000100110010010101110111111100011100000001)  
) LUT6_590 (
   .O(gates_590),
   .I0(InputBits[299]),
   .I1(InputBits[353]),
   .I2(InputBits[126]),
   .I3(InputBits[33]),
   .I4(InputBits[261]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0000001000100000001000111101001100010010000000100011001110001011)  
) LUT6_591 (
   .O(gates_591),
   .I0(InputBits[163]),
   .I1(InputBits[567]),
   .I2(InputBits[303]),
   .I3(InputBits[36]),
   .I4(InputBits[16]),
   .I5(InputBits[164])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000011001000000000001000100111001000110010)  
) LUT6_592 (
   .O(gates_592),
   .I0(InputBits[142]),
   .I1(InputBits[52]),
   .I2(InputBits[369]),
   .I3(InputBits[112]),
   .I4(InputBits[538]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000100011100000000010001110)  
) LUT6_593 (
   .O(gates_593),
   .I0(InputBits[272]),
   .I1(InputBits[364]),
   .I2(InputBits[250]),
   .I3(InputBits[78]),
   .I4(InputBits[88]),
   .I5(InputBits[572])
);
LUT6 #(
   .INIT(64'b0000000000011101000000001010101000000000011011110000100010001110)  
) LUT6_594 (
   .O(gates_594),
   .I0(InputBits[418]),
   .I1(InputBits[444]),
   .I2(InputBits[150]),
   .I3(InputBits[18]),
   .I4(InputBits[263]),
   .I5(InputBits[487])
);
LUT6 #(
   .INIT(64'b1001101110111111100010101010101010101110111111111111101011111111)  
) LUT6_595 (
   .O(gates_595),
   .I0(InputBits[390]),
   .I1(InputBits[137]),
   .I2(InputBits[202]),
   .I3(InputBits[83]),
   .I4(InputBits[311]),
   .I5(InputBits[104])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000100000000010101010000000001000101)  
) LUT6_596 (
   .O(gates_596),
   .I0(InputBits[535]),
   .I1(InputBits[197]),
   .I2(InputBits[494]),
   .I3(InputBits[576]),
   .I4(InputBits[155]),
   .I5(InputBits[13])
);
LUT6 #(
   .INIT(64'b0001000000000001000100000001000000010001000100110000000000000000)  
) LUT6_597 (
   .O(gates_597),
   .I0(InputBits[216]),
   .I1(InputBits[507]),
   .I2(InputBits[91]),
   .I3(InputBits[137]),
   .I4(InputBits[247]),
   .I5(InputBits[45])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010101111101000101111111110110011)  
) LUT6_598 (
   .O(gates_598),
   .I0(InputBits[178]),
   .I1(InputBits[425]),
   .I2(InputBits[249]),
   .I3(InputBits[398]),
   .I4(InputBits[108]),
   .I5(InputBits[385])
);
LUT6 #(
   .INIT(64'b0000000001000100000000001100010100000000010001010000000001001111)  
) LUT6_599 (
   .O(gates_599),
   .I0(InputBits[491]),
   .I1(InputBits[40]),
   .I2(InputBits[129]),
   .I3(InputBits[530]),
   .I4(InputBits[401]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000010011000000000000001100000001000000110000000000000010)  
) LUT6_600 (
   .O(gates_600),
   .I0(InputBits[456]),
   .I1(InputBits[505]),
   .I2(InputBits[434]),
   .I3(InputBits[219]),
   .I4(InputBits[416]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b1000111100001100110111110010111100001111100011010100111101011101)  
) LUT6_601 (
   .O(gates_601),
   .I0(InputBits[158]),
   .I1(InputBits[318]),
   .I2(InputBits[253]),
   .I3(InputBits[345]),
   .I4(InputBits[489]),
   .I5(InputBits[230])
);
LUT6 #(
   .INIT(64'b0000001000111011000010101010101000000011001110111010101011111010)  
) LUT6_602 (
   .O(gates_602),
   .I0(InputBits[373]),
   .I1(InputBits[67]),
   .I2(InputBits[157]),
   .I3(InputBits[299]),
   .I4(InputBits[174]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b0000101100000100000000010000000100011110010011110001011000010111)  
) LUT6_603 (
   .O(gates_603),
   .I0(InputBits[33]),
   .I1(InputBits[36]),
   .I2(InputBits[43]),
   .I3(InputBits[85]),
   .I4(InputBits[59]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0000000000000000010101010101010100000000000000000011100100010011)  
) LUT6_604 (
   .O(gates_604),
   .I0(InputBits[266]),
   .I1(InputBits[255]),
   .I2(InputBits[163]),
   .I3(InputBits[323]),
   .I4(InputBits[575]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b0011100100000111001010101010101000000101000001010111110101001111)  
) LUT6_605 (
   .O(gates_605),
   .I0(InputBits[498]),
   .I1(InputBits[323]),
   .I2(InputBits[497]),
   .I3(InputBits[152]),
   .I4(InputBits[404]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0011001100101111001001111011111100100011001000110000000110010011)  
) LUT6_606 (
   .O(gates_606),
   .I0(InputBits[267]),
   .I1(InputBits[516]),
   .I2(InputBits[219]),
   .I3(InputBits[523]),
   .I4(InputBits[301]),
   .I5(InputBits[341])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010000000000000000)  
) LUT6_607 (
   .O(gates_607),
   .I0(InputBits[459]),
   .I1(InputBits[506]),
   .I2(InputBits[531]),
   .I3(InputBits[89]),
   .I4(InputBits[320]),
   .I5(InputBits[552])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000011100000000000000000011100000111111)  
) LUT6_608 (
   .O(gates_608),
   .I0(InputBits[138]),
   .I1(InputBits[526]),
   .I2(InputBits[144]),
   .I3(InputBits[513]),
   .I4(InputBits[553]),
   .I5(InputBits[291])
);
LUT6 #(
   .INIT(64'b0000010100000111000001010000111100000101000010000000000000000010)  
) LUT6_609 (
   .O(gates_609),
   .I0(InputBits[17]),
   .I1(InputBits[403]),
   .I2(InputBits[22]),
   .I3(InputBits[203]),
   .I4(InputBits[210]),
   .I5(InputBits[350])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000000000101)  
) LUT6_610 (
   .O(gates_610),
   .I0(InputBits[2]),
   .I1(InputBits[170]),
   .I2(InputBits[531]),
   .I3(InputBits[97]),
   .I4(InputBits[481]),
   .I5(InputBits[127])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010001001100000001000100010101)  
) LUT6_611 (
   .O(gates_611),
   .I0(InputBits[53]),
   .I1(InputBits[242]),
   .I2(InputBits[417]),
   .I3(InputBits[67]),
   .I4(InputBits[512]),
   .I5(InputBits[572])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110011001100000000000000000011000000110000)  
) LUT6_612 (
   .O(gates_612),
   .I0(InputBits[429]),
   .I1(InputBits[1]),
   .I2(InputBits[372]),
   .I3(InputBits[449]),
   .I4(InputBits[529]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000101010100000000000000010000000011111101)  
) LUT6_613 (
   .O(gates_613),
   .I0(InputBits[562]),
   .I1(InputBits[249]),
   .I2(InputBits[305]),
   .I3(InputBits[241]),
   .I4(InputBits[252]),
   .I5(InputBits[135])
);
LUT6 #(
   .INIT(64'b0111001111111011011101010000000001110011111101110011011100110000)  
) LUT6_614 (
   .O(gates_614),
   .I0(InputBits[298]),
   .I1(InputBits[509]),
   .I2(InputBits[202]),
   .I3(InputBits[349]),
   .I4(InputBits[285]),
   .I5(InputBits[206])
);
LUT6 #(
   .INIT(64'b0000000000000000001100010011000100000000000000000011000100110101)  
) LUT6_615 (
   .O(gates_615),
   .I0(InputBits[251]),
   .I1(InputBits[551]),
   .I2(InputBits[398]),
   .I3(InputBits[429]),
   .I4(InputBits[121]),
   .I5(InputBits[154])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000110000000110)  
) LUT6_616 (
   .O(gates_616),
   .I0(InputBits[477]),
   .I1(InputBits[335]),
   .I2(InputBits[560]),
   .I3(InputBits[429]),
   .I4(InputBits[97]),
   .I5(InputBits[25])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000001100000011)  
) LUT6_617 (
   .O(gates_617),
   .I0(InputBits[469]),
   .I1(InputBits[111]),
   .I2(InputBits[22]),
   .I3(InputBits[168]),
   .I4(InputBits[23]),
   .I5(InputBits[457])
);
LUT6 #(
   .INIT(64'b0000000000001011000000100001101100000000000000000001000000010011)  
) LUT6_618 (
   .O(gates_618),
   .I0(InputBits[61]),
   .I1(InputBits[508]),
   .I2(InputBits[550]),
   .I3(InputBits[377]),
   .I4(InputBits[436]),
   .I5(InputBits[153])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000101111100001010)  
) LUT6_619 (
   .O(gates_619),
   .I0(InputBits[291]),
   .I1(InputBits[164]),
   .I2(InputBits[35]),
   .I3(InputBits[259]),
   .I4(InputBits[410]),
   .I5(InputBits[410])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001101111100000000010101010000000011001110)  
) LUT6_620 (
   .O(gates_620),
   .I0(InputBits[260]),
   .I1(InputBits[342]),
   .I2(InputBits[60]),
   .I3(InputBits[52]),
   .I4(InputBits[456]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0000110100000101000011010000110100001101000011010000110100001101)  
) LUT6_621 (
   .O(gates_621),
   .I0(InputBits[254]),
   .I1(InputBits[349]),
   .I2(InputBits[27]),
   .I3(InputBits[429]),
   .I4(InputBits[134]),
   .I5(InputBits[447])
);
LUT6 #(
   .INIT(64'b1111011101110010110100010111101001010000111000001100000111001100)  
) LUT6_622 (
   .O(gates_622),
   .I0(InputBits[339]),
   .I1(InputBits[189]),
   .I2(InputBits[283]),
   .I3(InputBits[396]),
   .I4(InputBits[328]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0000000000000101000000010001111100000000000000000000000000011011)  
) LUT6_623 (
   .O(gates_623),
   .I0(InputBits[432]),
   .I1(InputBits[254]),
   .I2(InputBits[460]),
   .I3(InputBits[558]),
   .I4(InputBits[75]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0000000000110010000000110011101100000000001100110000001000000000)  
) LUT6_624 (
   .O(gates_624),
   .I0(InputBits[440]),
   .I1(InputBits[535]),
   .I2(InputBits[62]),
   .I3(InputBits[216]),
   .I4(InputBits[503]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b0010001100000000001111100000000000000000000000010000000000111110)  
) LUT6_625 (
   .O(gates_625),
   .I0(InputBits[393]),
   .I1(InputBits[335]),
   .I2(InputBits[16]),
   .I3(InputBits[322]),
   .I4(InputBits[43]),
   .I5(InputBits[322])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000011001000100001111111111011000)  
) LUT6_626 (
   .O(gates_626),
   .I0(InputBits[157]),
   .I1(InputBits[181]),
   .I2(InputBits[118]),
   .I3(InputBits[370]),
   .I4(InputBits[127]),
   .I5(InputBits[217])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000010000011000001000101011011)  
) LUT6_627 (
   .O(gates_627),
   .I0(InputBits[168]),
   .I1(InputBits[250]),
   .I2(InputBits[163]),
   .I3(InputBits[88]),
   .I4(InputBits[192]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000010100001100000101000101010100010100)  
) LUT6_628 (
   .O(gates_628),
   .I0(InputBits[557]),
   .I1(InputBits[224]),
   .I2(InputBits[14]),
   .I3(InputBits[141]),
   .I4(InputBits[211]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0000000000000000010101010000000000000000000000000001010100000000)  
) LUT6_629 (
   .O(gates_629),
   .I0(InputBits[482]),
   .I1(InputBits[88]),
   .I2(InputBits[328]),
   .I3(InputBits[294]),
   .I4(InputBits[217]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0010001000111011000000001010001100100011101011110000011010100011)  
) LUT6_630 (
   .O(gates_630),
   .I0(InputBits[270]),
   .I1(InputBits[55]),
   .I2(InputBits[105]),
   .I3(InputBits[172]),
   .I4(InputBits[340]),
   .I5(InputBits[132])
);
LUT6 #(
   .INIT(64'b0000000000000001000000010000000100010000000101000001000000010101)  
) LUT6_631 (
   .O(gates_631),
   .I0(InputBits[123]),
   .I1(InputBits[527]),
   .I2(InputBits[408]),
   .I3(InputBits[491]),
   .I4(InputBits[127]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0000000000000111000001010000010100000000000001010000000100000101)  
) LUT6_632 (
   .O(gates_632),
   .I0(InputBits[506]),
   .I1(InputBits[383]),
   .I2(InputBits[532]),
   .I3(InputBits[9]),
   .I4(InputBits[89]),
   .I5(InputBits[321])
);
LUT6 #(
   .INIT(64'b0101000001010101010001000101010100000000010101000000000000010001)  
) LUT6_633 (
   .O(gates_633),
   .I0(InputBits[337]),
   .I1(InputBits[377]),
   .I2(InputBits[162]),
   .I3(InputBits[540]),
   .I4(InputBits[380]),
   .I5(InputBits[291])
);
LUT6 #(
   .INIT(64'b0000000100000000000000110000000100000010000000000000001100000000)  
) LUT6_634 (
   .O(gates_634),
   .I0(InputBits[35]),
   .I1(InputBits[559]),
   .I2(InputBits[74]),
   .I3(InputBits[342]),
   .I4(InputBits[232]),
   .I5(InputBits[317])
);
LUT6 #(
   .INIT(64'b0000111000000000000111010010101100001000000010000001111100010011)  
) LUT6_635 (
   .O(gates_635),
   .I0(InputBits[376]),
   .I1(InputBits[425]),
   .I2(InputBits[470]),
   .I3(InputBits[467]),
   .I4(InputBits[124]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b0000000000001000000000000000000100000010000011100000000000011110)  
) LUT6_636 (
   .O(gates_636),
   .I0(InputBits[367]),
   .I1(InputBits[501]),
   .I2(InputBits[5]),
   .I3(InputBits[337]),
   .I4(InputBits[322]),
   .I5(InputBits[573])
);
LUT6 #(
   .INIT(64'b0000000000001010000000000000010000000000000000000001010100000000)  
) LUT6_637 (
   .O(gates_637),
   .I0(InputBits[209]),
   .I1(InputBits[161]),
   .I2(InputBits[542]),
   .I3(InputBits[166]),
   .I4(InputBits[209]),
   .I5(InputBits[548])
);
LUT6 #(
   .INIT(64'b0000100000011000010001010100010110011101010110110011111100100100)  
) LUT6_638 (
   .O(gates_638),
   .I0(InputBits[45]),
   .I1(InputBits[388]),
   .I2(InputBits[302]),
   .I3(InputBits[225]),
   .I4(InputBits[44]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0000010001000000011001011110010011111110110011001111111111101111)  
) LUT6_639 (
   .O(gates_639),
   .I0(InputBits[323]),
   .I1(InputBits[202]),
   .I2(InputBits[352]),
   .I3(InputBits[310]),
   .I4(InputBits[274]),
   .I5(InputBits[435])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001101010111110100111101111000)  
) LUT6_640 (
   .O(gates_640),
   .I0(InputBits[92]),
   .I1(InputBits[158]),
   .I2(InputBits[335]),
   .I3(InputBits[191]),
   .I4(InputBits[417]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0001000001010100000000000101000100000000011100000000000001010000)  
) LUT6_641 (
   .O(gates_641),
   .I0(InputBits[52]),
   .I1(InputBits[69]),
   .I2(InputBits[372]),
   .I3(InputBits[541]),
   .I4(InputBits[305]),
   .I5(InputBits[117])
);
LUT6 #(
   .INIT(64'b1011001111111111111111111111111100100000000000000011000000000011)  
) LUT6_642 (
   .O(gates_642),
   .I0(InputBits[210]),
   .I1(InputBits[490]),
   .I2(InputBits[273]),
   .I3(InputBits[297]),
   .I4(InputBits[473]),
   .I5(InputBits[342])
);
LUT6 #(
   .INIT(64'b0000000001100111000000000100110000000000010011000000000001001100)  
) LUT6_643 (
   .O(gates_643),
   .I0(InputBits[352]),
   .I1(InputBits[268]),
   .I2(InputBits[63]),
   .I3(InputBits[145]),
   .I4(InputBits[203]),
   .I5(InputBits[115])
);
LUT6 #(
   .INIT(64'b0000000000000000010000010100000100000001000000010100000111000011)  
) LUT6_644 (
   .O(gates_644),
   .I0(InputBits[81]),
   .I1(InputBits[299]),
   .I2(InputBits[299]),
   .I3(InputBits[159]),
   .I4(InputBits[108]),
   .I5(InputBits[231])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001001110101010000111111100110000)  
) LUT6_645 (
   .O(gates_645),
   .I0(InputBits[115]),
   .I1(InputBits[405]),
   .I2(InputBits[296]),
   .I3(InputBits[221]),
   .I4(InputBits[133]),
   .I5(InputBits[266])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000001111011110000000110101110)  
) LUT6_646 (
   .O(gates_646),
   .I0(InputBits[245]),
   .I1(InputBits[93]),
   .I2(InputBits[220]),
   .I3(InputBits[384]),
   .I4(InputBits[324]),
   .I5(InputBits[561])
);
LUT6 #(
   .INIT(64'b0000000101000100000001010001001100000101010101000100010101010101)  
) LUT6_647 (
   .O(gates_647),
   .I0(InputBits[567]),
   .I1(InputBits[37]),
   .I2(InputBits[437]),
   .I3(InputBits[11]),
   .I4(InputBits[108]),
   .I5(InputBits[329])
);
LUT6 #(
   .INIT(64'b0000000000100000001100111010110000000000000100000001001111110001)  
) LUT6_648 (
   .O(gates_648),
   .I0(InputBits[426]),
   .I1(InputBits[17]),
   .I2(InputBits[375]),
   .I3(InputBits[243]),
   .I4(InputBits[52]),
   .I5(InputBits[400])
);
LUT6 #(
   .INIT(64'b0010001100100010001110110011001100001010000000010011101100110011)  
) LUT6_649 (
   .O(gates_649),
   .I0(InputBits[60]),
   .I1(InputBits[9]),
   .I2(InputBits[487]),
   .I3(InputBits[423]),
   .I4(InputBits[253]),
   .I5(InputBits[478])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000010000000000000001000000000110010001)  
) LUT6_650 (
   .O(gates_650),
   .I0(InputBits[184]),
   .I1(InputBits[210]),
   .I2(InputBits[9]),
   .I3(InputBits[205]),
   .I4(InputBits[75]),
   .I5(InputBits[227])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010101010101000100010011000101000001010101)  
) LUT6_651 (
   .O(gates_651),
   .I0(InputBits[409]),
   .I1(InputBits[320]),
   .I2(InputBits[439]),
   .I3(InputBits[130]),
   .I4(InputBits[226]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010100000000111011000000000011101100)  
) LUT6_652 (
   .O(gates_652),
   .I0(InputBits[156]),
   .I1(InputBits[342]),
   .I2(InputBits[39]),
   .I3(InputBits[122]),
   .I4(InputBits[38]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0000000100000101000000010000000000000001000001010001000100010101)  
) LUT6_653 (
   .O(gates_653),
   .I0(InputBits[22]),
   .I1(InputBits[41]),
   .I2(InputBits[480]),
   .I3(InputBits[383]),
   .I4(InputBits[260]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000000001000000110000000000000001)  
) LUT6_654 (
   .O(gates_654),
   .I0(InputBits[485]),
   .I1(InputBits[104]),
   .I2(InputBits[559]),
   .I3(InputBits[558]),
   .I4(InputBits[320]),
   .I5(InputBits[150])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010011001100000000000000000011001100000001)  
) LUT6_655 (
   .O(gates_655),
   .I0(InputBits[404]),
   .I1(InputBits[19]),
   .I2(InputBits[110]),
   .I3(InputBits[479]),
   .I4(InputBits[558]),
   .I5(InputBits[41])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001110100111100001101010101010100)  
) LUT6_656 (
   .O(gates_656),
   .I0(InputBits[227]),
   .I1(InputBits[430]),
   .I2(InputBits[392]),
   .I3(InputBits[443]),
   .I4(InputBits[273]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0000000000000001111011011111101100000000000000001010000010101000)  
) LUT6_657 (
   .O(gates_657),
   .I0(InputBits[479]),
   .I1(InputBits[427]),
   .I2(InputBits[416]),
   .I3(InputBits[437]),
   .I4(InputBits[562]),
   .I5(InputBits[419])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001010101000101010001000000010111)  
) LUT6_658 (
   .O(gates_658),
   .I0(InputBits[250]),
   .I1(InputBits[402]),
   .I2(InputBits[60]),
   .I3(InputBits[110]),
   .I4(InputBits[501]),
   .I5(InputBits[122])
);
LUT6 #(
   .INIT(64'b1001111111111111110111111101111100001101000011110000111100001111)  
) LUT6_659 (
   .O(gates_659),
   .I0(InputBits[184]),
   .I1(InputBits[454]),
   .I2(InputBits[251]),
   .I3(InputBits[470]),
   .I4(InputBits[302]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000001100000000000000000000000000000011)  
) LUT6_660 (
   .O(gates_660),
   .I0(InputBits[291]),
   .I1(InputBits[24]),
   .I2(InputBits[2]),
   .I3(InputBits[483]),
   .I4(InputBits[555]),
   .I5(InputBits[363])
);
LUT6 #(
   .INIT(64'b0011001100110000001100000011100000110011001100100011100000111110)  
) LUT6_661 (
   .O(gates_661),
   .I0(InputBits[324]),
   .I1(InputBits[480]),
   .I2(InputBits[286]),
   .I3(InputBits[423]),
   .I4(InputBits[272]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b0000000000000000111011111110111000000100010001001000111110101110)  
) LUT6_662 (
   .O(gates_662),
   .I0(InputBits[286]),
   .I1(InputBits[346]),
   .I2(InputBits[255]),
   .I3(InputBits[283]),
   .I4(InputBits[31]),
   .I5(InputBits[248])
);
LUT6 #(
   .INIT(64'b0110000001100100010101000111010101100000111000100111011011111111)  
) LUT6_663 (
   .O(gates_663),
   .I0(InputBits[384]),
   .I1(InputBits[222]),
   .I2(InputBits[423]),
   .I3(InputBits[102]),
   .I4(InputBits[251]),
   .I5(InputBits[114])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000100101100000001011111111)  
) LUT6_664 (
   .O(gates_664),
   .I0(InputBits[233]),
   .I1(InputBits[137]),
   .I2(InputBits[113]),
   .I3(InputBits[256]),
   .I4(InputBits[54]),
   .I5(InputBits[529])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001010110111110000000000001011)  
) LUT6_665 (
   .O(gates_665),
   .I0(InputBits[321]),
   .I1(InputBits[257]),
   .I2(InputBits[81]),
   .I3(InputBits[123]),
   .I4(InputBits[293]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b0000000000000101000001000000010100000000000000010000010000000001)  
) LUT6_666 (
   .O(gates_666),
   .I0(InputBits[265]),
   .I1(InputBits[153]),
   .I2(InputBits[169]),
   .I3(InputBits[82]),
   .I4(InputBits[355]),
   .I5(InputBits[467])
);
LUT6 #(
   .INIT(64'b0000010000000000000001110000010100000110000001000000111100001110)  
) LUT6_667 (
   .O(gates_667),
   .I0(InputBits[544]),
   .I1(InputBits[398]),
   .I2(InputBits[241]),
   .I3(InputBits[390]),
   .I4(InputBits[149]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001010101000000000010101010000000111101111)  
) LUT6_668 (
   .O(gates_668),
   .I0(InputBits[213]),
   .I1(InputBits[415]),
   .I2(InputBits[133]),
   .I3(InputBits[5]),
   .I4(InputBits[9]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000010100000101000000010100001100000101000011110101101100001111)  
) LUT6_669 (
   .O(gates_669),
   .I0(InputBits[70]),
   .I1(InputBits[127]),
   .I2(InputBits[54]),
   .I3(InputBits[135]),
   .I4(InputBits[339]),
   .I5(InputBits[403])
);
LUT6 #(
   .INIT(64'b0000010000000101000001000000010011110111111000111111011111100011)  
) LUT6_670 (
   .O(gates_670),
   .I0(InputBits[176]),
   .I1(InputBits[58]),
   .I2(InputBits[152]),
   .I3(InputBits[430]),
   .I4(InputBits[87]),
   .I5(InputBits[9])
);
LUT6 #(
   .INIT(64'b0000111100001111000011110000111100001011000011110000001000001011)  
) LUT6_671 (
   .O(gates_671),
   .I0(InputBits[443]),
   .I1(InputBits[105]),
   .I2(InputBits[241]),
   .I3(InputBits[298]),
   .I4(InputBits[369]),
   .I5(InputBits[246])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000110000001010000110100001100)  
) LUT6_672 (
   .O(gates_672),
   .I0(InputBits[216]),
   .I1(InputBits[420]),
   .I2(InputBits[530]),
   .I3(InputBits[246]),
   .I4(InputBits[168]),
   .I5(InputBits[147])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000010000000111110000000010111111111)  
) LUT6_673 (
   .O(gates_673),
   .I0(InputBits[499]),
   .I1(InputBits[468]),
   .I2(InputBits[63]),
   .I3(InputBits[227]),
   .I4(InputBits[127]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000100010100000101010100010000000001010001)  
) LUT6_674 (
   .O(gates_674),
   .I0(InputBits[145]),
   .I1(InputBits[299]),
   .I2(InputBits[359]),
   .I3(InputBits[570]),
   .I4(InputBits[282]),
   .I5(InputBits[408])
);
LUT6 #(
   .INIT(64'b0000000000110000000000110000000000010000000000100000000100110000)  
) LUT6_675 (
   .O(gates_675),
   .I0(InputBits[445]),
   .I1(InputBits[553]),
   .I2(InputBits[320]),
   .I3(InputBits[480]),
   .I4(InputBits[174]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b0000011100000000000010110000101100001111000001010000111100000111)  
) LUT6_676 (
   .O(gates_676),
   .I0(InputBits[499]),
   .I1(InputBits[488]),
   .I2(InputBits[556]),
   .I3(InputBits[165]),
   .I4(InputBits[403]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0000000000000000000001110101000000000000000000000000010100010111)  
) LUT6_677 (
   .O(gates_677),
   .I0(InputBits[513]),
   .I1(InputBits[111]),
   .I2(InputBits[61]),
   .I3(InputBits[312]),
   .I4(InputBits[28]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0001010101010101000000000000000000010001010101010001000101000111)  
) LUT6_678 (
   .O(gates_678),
   .I0(InputBits[528]),
   .I1(InputBits[31]),
   .I2(InputBits[82]),
   .I3(InputBits[175]),
   .I4(InputBits[368]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0000001100000001011100111011100011110111001110111111001110110000)  
) LUT6_679 (
   .O(gates_679),
   .I0(InputBits[442]),
   .I1(InputBits[82]),
   .I2(InputBits[348]),
   .I3(InputBits[248]),
   .I4(InputBits[215]),
   .I5(InputBits[68])
);
LUT6 #(
   .INIT(64'b0000010101010011000000011111001100000001111100110000010100110111)  
) LUT6_680 (
   .O(gates_680),
   .I0(InputBits[56]),
   .I1(InputBits[472]),
   .I2(InputBits[432]),
   .I3(InputBits[69]),
   .I4(InputBits[182]),
   .I5(InputBits[185])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000001010000000100000101)  
) LUT6_681 (
   .O(gates_681),
   .I0(InputBits[3]),
   .I1(InputBits[13]),
   .I2(InputBits[536]),
   .I3(InputBits[479]),
   .I4(InputBits[455]),
   .I5(InputBits[169])
);
LUT6 #(
   .INIT(64'b0000001100000011000000111011101100000000000000010010011000100011)  
) LUT6_682 (
   .O(gates_682),
   .I0(InputBits[307]),
   .I1(InputBits[194]),
   .I2(InputBits[497]),
   .I3(InputBits[489]),
   .I4(InputBits[228]),
   .I5(InputBits[346])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000101000010010000101100001011)  
) LUT6_683 (
   .O(gates_683),
   .I0(InputBits[142]),
   .I1(InputBits[490]),
   .I2(InputBits[556]),
   .I3(InputBits[158]),
   .I4(InputBits[192]),
   .I5(InputBits[434])
);
LUT6 #(
   .INIT(64'b0000001100000001000000000000000000000111011001110000010101100111)  
) LUT6_684 (
   .O(gates_684),
   .I0(InputBits[564]),
   .I1(InputBits[453]),
   .I2(InputBits[277]),
   .I3(InputBits[133]),
   .I4(InputBits[211]),
   .I5(InputBits[229])
);
LUT6 #(
   .INIT(64'b0101011100010001010000100000000101011111010100110101010101010111)  
) LUT6_685 (
   .O(gates_685),
   .I0(InputBits[534]),
   .I1(InputBits[110]),
   .I2(InputBits[452]),
   .I3(InputBits[390]),
   .I4(InputBits[188]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010110001010100101111100111010)  
) LUT6_686 (
   .O(gates_686),
   .I0(InputBits[309]),
   .I1(InputBits[90]),
   .I2(InputBits[38]),
   .I3(InputBits[477]),
   .I4(InputBits[158]),
   .I5(InputBits[569])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000011110000000000110010)  
) LUT6_687 (
   .O(gates_687),
   .I0(InputBits[350]),
   .I1(InputBits[510]),
   .I2(InputBits[550]),
   .I3(InputBits[75]),
   .I4(InputBits[383]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0001000100000000000100010000000000010001100000110101000111110011)  
) LUT6_688 (
   .O(gates_688),
   .I0(InputBits[480]),
   .I1(InputBits[255]),
   .I2(InputBits[302]),
   .I3(InputBits[260]),
   .I4(InputBits[447]),
   .I5(InputBits[564])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000001110111011101110011011100110011)  
) LUT6_689 (
   .O(gates_689),
   .I0(InputBits[14]),
   .I1(InputBits[493]),
   .I2(InputBits[329]),
   .I3(InputBits[89]),
   .I4(InputBits[421]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000010000100010010100100101111001111111011)  
) LUT6_690 (
   .O(gates_690),
   .I0(InputBits[166]),
   .I1(InputBits[539]),
   .I2(InputBits[214]),
   .I3(InputBits[522]),
   .I4(InputBits[278]),
   .I5(InputBits[13])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000001000000110011000000110001)  
) LUT6_691 (
   .O(gates_691),
   .I0(InputBits[508]),
   .I1(InputBits[457]),
   .I2(InputBits[68]),
   .I3(InputBits[130]),
   .I4(InputBits[119]),
   .I5(InputBits[572])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100010111011001010001011101110)  
) LUT6_692 (
   .O(gates_692),
   .I0(InputBits[366]),
   .I1(InputBits[502]),
   .I2(InputBits[475]),
   .I3(InputBits[272]),
   .I4(InputBits[257]),
   .I5(InputBits[51])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000000000000001)  
) LUT6_693 (
   .O(gates_693),
   .I0(InputBits[452]),
   .I1(InputBits[111]),
   .I2(InputBits[557]),
   .I3(InputBits[170]),
   .I4(InputBits[195]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0000000010100011011000001111111100000000101000101001001011110011)  
) LUT6_694 (
   .O(gates_694),
   .I0(InputBits[346]),
   .I1(InputBits[302]),
   .I2(InputBits[325]),
   .I3(InputBits[338]),
   .I4(InputBits[83]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0000001111011111000010111010001000000101111111101001011111111010)  
) LUT6_695 (
   .O(gates_695),
   .I0(InputBits[345]),
   .I1(InputBits[404]),
   .I2(InputBits[406]),
   .I3(InputBits[167]),
   .I4(InputBits[388]),
   .I5(InputBits[297])
);
LUT6 #(
   .INIT(64'b0001000011011111000010000011111101010000110111110011100100011111)  
) LUT6_696 (
   .O(gates_696),
   .I0(InputBits[438]),
   .I1(InputBits[213]),
   .I2(InputBits[94]),
   .I3(InputBits[255]),
   .I4(InputBits[189]),
   .I5(InputBits[424])
);
LUT6 #(
   .INIT(64'b0000010101010101000000000000001001010101010101010000000000000000)  
) LUT6_697 (
   .O(gates_697),
   .I0(InputBits[9]),
   .I1(InputBits[57]),
   .I2(InputBits[378]),
   .I3(InputBits[101]),
   .I4(InputBits[371]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0000000000000000000011100100111000001000000000001100111000011111)  
) LUT6_698 (
   .O(gates_698),
   .I0(InputBits[389]),
   .I1(InputBits[391]),
   .I2(InputBits[75]),
   .I3(InputBits[356]),
   .I4(InputBits[21]),
   .I5(InputBits[132])
);
LUT6 #(
   .INIT(64'b0000000001010011000000001100010000000000111111110000001011111111)  
) LUT6_699 (
   .O(gates_699),
   .I0(InputBits[138]),
   .I1(InputBits[455]),
   .I2(InputBits[62]),
   .I3(InputBits[21]),
   .I4(InputBits[180]),
   .I5(InputBits[206])
);
LUT6 #(
   .INIT(64'b0000000010001111000000000000100000000001110111110000010100001100)  
) LUT6_700 (
   .O(gates_700),
   .I0(InputBits[61]),
   .I1(InputBits[198]),
   .I2(InputBits[182]),
   .I3(InputBits[70]),
   .I4(InputBits[418]),
   .I5(InputBits[173])
);
LUT6 #(
   .INIT(64'b0000001100001111000100110001111100010011001100110001110000010100)  
) LUT6_701 (
   .O(gates_701),
   .I0(InputBits[205]),
   .I1(InputBits[312]),
   .I2(InputBits[546]),
   .I3(InputBits[496]),
   .I4(InputBits[261]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0000001100000010000000110000111100000000000000000000001000000011)  
) LUT6_702 (
   .O(gates_702),
   .I0(InputBits[186]),
   .I1(InputBits[511]),
   .I2(InputBits[576]),
   .I3(InputBits[219]),
   .I4(InputBits[79]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0000000000000100000000001010001011001100111011101010001011101111)  
) LUT6_703 (
   .O(gates_703),
   .I0(InputBits[287]),
   .I1(InputBits[320]),
   .I2(InputBits[426]),
   .I3(InputBits[485]),
   .I4(InputBits[400]),
   .I5(InputBits[104])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000101010100000000000000000001010011111000)  
) LUT6_704 (
   .O(gates_704),
   .I0(InputBits[118]),
   .I1(InputBits[174]),
   .I2(InputBits[319]),
   .I3(InputBits[33]),
   .I4(InputBits[241]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000000000001110000011110000111100000000000010000000110100000000)  
) LUT6_705 (
   .O(gates_705),
   .I0(InputBits[389]),
   .I1(InputBits[188]),
   .I2(InputBits[574]),
   .I3(InputBits[39]),
   .I4(InputBits[182]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0000000000000000000011110000110100000000000000000000110100001101)  
) LUT6_706 (
   .O(gates_706),
   .I0(InputBits[126]),
   .I1(InputBits[221]),
   .I2(InputBits[362]),
   .I3(InputBits[243]),
   .I4(InputBits[385]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010011001100000000000000000000000000000011)  
) LUT6_707 (
   .O(gates_707),
   .I0(InputBits[154]),
   .I1(InputBits[553]),
   .I2(InputBits[111]),
   .I3(InputBits[54]),
   .I4(InputBits[169]),
   .I5(InputBits[408])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000010100000000000000000001011100000001)  
) LUT6_708 (
   .O(gates_708),
   .I0(InputBits[21]),
   .I1(InputBits[425]),
   .I2(InputBits[361]),
   .I3(InputBits[340]),
   .I4(InputBits[560]),
   .I5(InputBits[32])
);
LUT6 #(
   .INIT(64'b0000001100000111000000100000001100001111000011110000000000001011)  
) LUT6_709 (
   .O(gates_709),
   .I0(InputBits[65]),
   .I1(InputBits[104]),
   .I2(InputBits[576]),
   .I3(InputBits[487]),
   .I4(InputBits[414]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0000000011001100001111110000000010101100000001001011111110101010)  
) LUT6_710 (
   .O(gates_710),
   .I0(InputBits[344]),
   .I1(InputBits[498]),
   .I2(InputBits[379]),
   .I3(InputBits[373]),
   .I4(InputBits[547]),
   .I5(InputBits[301])
);
LUT6 #(
   .INIT(64'b0001000001010101000100000101111100000000000100010000000000010001)  
) LUT6_711 (
   .O(gates_711),
   .I0(InputBits[31]),
   .I1(InputBits[208]),
   .I2(InputBits[116]),
   .I3(InputBits[123]),
   .I4(InputBits[141]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0000000000000000001000100011001100000000000100010000010100100000)  
) LUT6_712 (
   .O(gates_712),
   .I0(InputBits[416]),
   .I1(InputBits[551]),
   .I2(InputBits[153]),
   .I3(InputBits[527]),
   .I4(InputBits[266]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0000001011111111000000001111111100000010000011110000001100001111)  
) LUT6_713 (
   .O(gates_713),
   .I0(InputBits[430]),
   .I1(InputBits[453]),
   .I2(InputBits[508]),
   .I3(InputBits[253]),
   .I4(InputBits[135]),
   .I5(InputBits[464])
);
LUT6 #(
   .INIT(64'b1010000011111111111010101111101001000100100001001111111111111111)  
) LUT6_714 (
   .O(gates_714),
   .I0(InputBits[326]),
   .I1(InputBits[139]),
   .I2(InputBits[501]),
   .I3(InputBits[490]),
   .I4(InputBits[353]),
   .I5(InputBits[305])
);
LUT6 #(
   .INIT(64'b1111111111011111111111111101011101010011000100111101111101000101)  
) LUT6_715 (
   .O(gates_715),
   .I0(InputBits[275]),
   .I1(InputBits[477]),
   .I2(InputBits[82]),
   .I3(InputBits[394]),
   .I4(InputBits[294]),
   .I5(InputBits[342])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011001000110000000000000010)  
) LUT6_716 (
   .O(gates_716),
   .I0(InputBits[441]),
   .I1(InputBits[458]),
   .I2(InputBits[355]),
   .I3(InputBits[468]),
   .I4(InputBits[455]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000010000000101000001010000010100000101000001110000000000000001)  
) LUT6_717 (
   .O(gates_717),
   .I0(InputBits[18]),
   .I1(InputBits[303]),
   .I2(InputBits[313]),
   .I3(InputBits[495]),
   .I4(InputBits[397]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000001000100000000000000010000000000000001)  
) LUT6_718 (
   .O(gates_718),
   .I0(InputBits[487]),
   .I1(InputBits[534]),
   .I2(InputBits[410]),
   .I3(InputBits[145]),
   .I4(InputBits[527]),
   .I5(InputBits[196])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000000000000000000001010000010000000101)  
) LUT6_719 (
   .O(gates_719),
   .I0(InputBits[170]),
   .I1(InputBits[500]),
   .I2(InputBits[146]),
   .I3(InputBits[481]),
   .I4(InputBits[37]),
   .I5(InputBits[251])
);
LUT6 #(
   .INIT(64'b0000000100010011110111110000110100000001000101111111111100001111)  
) LUT6_720 (
   .O(gates_720),
   .I0(InputBits[487]),
   .I1(InputBits[358]),
   .I2(InputBits[251]),
   .I3(InputBits[179]),
   .I4(InputBits[549]),
   .I5(InputBits[86])
);
LUT6 #(
   .INIT(64'b0100111100011101001111110011110100001111011111110101111101111101)  
) LUT6_721 (
   .O(gates_721),
   .I0(InputBits[472]),
   .I1(InputBits[316]),
   .I2(InputBits[502]),
   .I3(InputBits[223]),
   .I4(InputBits[340]),
   .I5(InputBits[210])
);
LUT6 #(
   .INIT(64'b1000000000000011001000000000000000110011001011110010001010101011)  
) LUT6_722 (
   .O(gates_722),
   .I0(InputBits[397]),
   .I1(InputBits[77]),
   .I2(InputBits[83]),
   .I3(InputBits[154]),
   .I4(InputBits[140]),
   .I5(InputBits[510])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000101000111001000000101011110101111)  
) LUT6_723 (
   .O(gates_723),
   .I0(InputBits[550]),
   .I1(InputBits[163]),
   .I2(InputBits[274]),
   .I3(InputBits[419]),
   .I4(InputBits[184]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000000000100000000000000010000000000000000)  
) LUT6_724 (
   .O(gates_724),
   .I0(InputBits[48]),
   .I1(InputBits[576]),
   .I2(InputBits[173]),
   .I3(InputBits[458]),
   .I4(InputBits[197]),
   .I5(InputBits[295])
);
LUT6 #(
   .INIT(64'b0000000001010101110010001101101000000000110111111011101011111010)  
) LUT6_725 (
   .O(gates_725),
   .I0(InputBits[372]),
   .I1(InputBits[441]),
   .I2(InputBits[236]),
   .I3(InputBits[148]),
   .I4(InputBits[263]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0100000111011101000000000101000000001011011111110000000010111100)  
) LUT6_726 (
   .O(gates_726),
   .I0(InputBits[336]),
   .I1(InputBits[181]),
   .I2(InputBits[248]),
   .I3(InputBits[56]),
   .I4(InputBits[415]),
   .I5(InputBits[164])
);
LUT6 #(
   .INIT(64'b0001111100000010000100110000000000000010000000100000001100001111)  
) LUT6_727 (
   .O(gates_727),
   .I0(InputBits[399]),
   .I1(InputBits[410]),
   .I2(InputBits[571]),
   .I3(InputBits[210]),
   .I4(InputBits[447]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000001100000000000000010000000011111001)  
) LUT6_728 (
   .O(gates_728),
   .I0(InputBits[449]),
   .I1(InputBits[451]),
   .I2(InputBits[13]),
   .I3(InputBits[489]),
   .I4(InputBits[151]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000000010000010100000001000000000001000101010101110111011111)  
) LUT6_729 (
   .O(gates_729),
   .I0(InputBits[567]),
   .I1(InputBits[306]),
   .I2(InputBits[158]),
   .I3(InputBits[189]),
   .I4(InputBits[13]),
   .I5(InputBits[229])
);
LUT6 #(
   .INIT(64'b0001010100000001000000010000000000000101000101010000000100000000)  
) LUT6_730 (
   .O(gates_730),
   .I0(InputBits[193]),
   .I1(InputBits[507]),
   .I2(InputBits[361]),
   .I3(InputBits[420]),
   .I4(InputBits[365]),
   .I5(InputBits[301])
);
LUT6 #(
   .INIT(64'b0001000100010001000100010000000100010001000101010000000000000001)  
) LUT6_731 (
   .O(gates_731),
   .I0(InputBits[575]),
   .I1(InputBits[20]),
   .I2(InputBits[82]),
   .I3(InputBits[446]),
   .I4(InputBits[198]),
   .I5(InputBits[201])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010000000000010000000000000001)  
) LUT6_732 (
   .O(gates_732),
   .I0(InputBits[111]),
   .I1(InputBits[574]),
   .I2(InputBits[426]),
   .I3(InputBits[404]),
   .I4(InputBits[160]),
   .I5(InputBits[540])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000000000000000000001000110000000000101000)  
) LUT6_733 (
   .O(gates_733),
   .I0(InputBits[428]),
   .I1(InputBits[43]),
   .I2(InputBits[32]),
   .I3(InputBits[147]),
   .I4(InputBits[284]),
   .I5(InputBits[227])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000000000000000000000000001111001110)  
) LUT6_734 (
   .O(gates_734),
   .I0(InputBits[346]),
   .I1(InputBits[45]),
   .I2(InputBits[485]),
   .I3(InputBits[243]),
   .I4(InputBits[47]),
   .I5(InputBits[195])
);
LUT6 #(
   .INIT(64'b0000000000010011000000010001001100000000000000000001001100010011)  
) LUT6_735 (
   .O(gates_735),
   .I0(InputBits[329]),
   .I1(InputBits[194]),
   .I2(InputBits[184]),
   .I3(InputBits[43]),
   .I4(InputBits[103]),
   .I5(InputBits[175])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000000100000001000101110000011000010101)  
) LUT6_736 (
   .O(gates_736),
   .I0(InputBits[492]),
   .I1(InputBits[243]),
   .I2(InputBits[33]),
   .I3(InputBits[290]),
   .I4(InputBits[247]),
   .I5(InputBits[240])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001010000010110000011000000111)  
) LUT6_737 (
   .O(gates_737),
   .I0(InputBits[502]),
   .I1(InputBits[181]),
   .I2(InputBits[337]),
   .I3(InputBits[108]),
   .I4(InputBits[450]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0100010001001101110101011101110101010101000011000101010111001100)  
) LUT6_738 (
   .O(gates_738),
   .I0(InputBits[508]),
   .I1(InputBits[395]),
   .I2(InputBits[427]),
   .I3(InputBits[479]),
   .I4(InputBits[206]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0000000000000000010000001100000000000000000000001000001000000000)  
) LUT6_739 (
   .O(gates_739),
   .I0(InputBits[42]),
   .I1(InputBits[296]),
   .I2(InputBits[296]),
   .I3(InputBits[324]),
   .I4(InputBits[551]),
   .I5(InputBits[202])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010100000000000000000000000001010101)  
) LUT6_740 (
   .O(gates_740),
   .I0(InputBits[533]),
   .I1(InputBits[139]),
   .I2(InputBits[567]),
   .I3(InputBits[552]),
   .I4(InputBits[265]),
   .I5(InputBits[455])
);
LUT6 #(
   .INIT(64'b0000000100000001000000110000000000000001000000110000011100000000)  
) LUT6_741 (
   .O(gates_741),
   .I0(InputBits[546]),
   .I1(InputBits[459]),
   .I2(InputBits[49]),
   .I3(InputBits[420]),
   .I4(InputBits[244]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b0000000000010011000000000001000000000000001000010000000000010001)  
) LUT6_742 (
   .O(gates_742),
   .I0(InputBits[487]),
   .I1(InputBits[193]),
   .I2(InputBits[64]),
   .I3(InputBits[541]),
   .I4(InputBits[408]),
   .I5(InputBits[426])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000100000000000001010)  
) LUT6_743 (
   .O(gates_743),
   .I0(InputBits[318]),
   .I1(InputBits[541]),
   .I2(InputBits[29]),
   .I3(InputBits[571]),
   .I4(InputBits[132]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b1011000000100011001100110011100111100100011000110011011000101110)  
) LUT6_744 (
   .O(gates_744),
   .I0(InputBits[199]),
   .I1(InputBits[243]),
   .I2(InputBits[380]),
   .I3(InputBits[315]),
   .I4(InputBits[428]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110000001100000011000000110000)  
) LUT6_745 (
   .O(gates_745),
   .I0(InputBits[220]),
   .I1(InputBits[3]),
   .I2(InputBits[260]),
   .I3(InputBits[363]),
   .I4(InputBits[113]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0000000000001100000000000000110011011111010011111111111100001111)  
) LUT6_746 (
   .O(gates_746),
   .I0(InputBits[155]),
   .I1(InputBits[320]),
   .I2(InputBits[275]),
   .I3(InputBits[431]),
   .I4(InputBits[162]),
   .I5(InputBits[540])
);
LUT6 #(
   .INIT(64'b0001010101000101010101010101010100000000000111110001010100000101)  
) LUT6_747 (
   .O(gates_747),
   .I0(InputBits[565]),
   .I1(InputBits[136]),
   .I2(InputBits[299]),
   .I3(InputBits[61]),
   .I4(InputBits[273]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0100010100000100000001010000010101000100010100000101010101010100)  
) LUT6_748 (
   .O(gates_748),
   .I0(InputBits[505]),
   .I1(InputBits[422]),
   .I2(InputBits[408]),
   .I3(InputBits[198]),
   .I4(InputBits[303]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000111010100000101000000000101010111110101)  
) LUT6_749 (
   .O(gates_749),
   .I0(InputBits[435]),
   .I1(InputBits[160]),
   .I2(InputBits[282]),
   .I3(InputBits[335]),
   .I4(InputBits[126]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0000100000000000000010100000111100001100000000000000101000001001)  
) LUT6_750 (
   .O(gates_750),
   .I0(InputBits[320]),
   .I1(InputBits[328]),
   .I2(InputBits[3]),
   .I3(InputBits[249]),
   .I4(InputBits[561]),
   .I5(InputBits[393])
);
LUT6 #(
   .INIT(64'b0000000011001000000000000111011100000000000000000000000000000011)  
) LUT6_751 (
   .O(gates_751),
   .I0(InputBits[475]),
   .I1(InputBits[148]),
   .I2(InputBits[231]),
   .I3(InputBits[561]),
   .I4(InputBits[75]),
   .I5(InputBits[346])
);
LUT6 #(
   .INIT(64'b0001000000000000000111110001000000000000000001010001011100010101)  
) LUT6_752 (
   .O(gates_752),
   .I0(InputBits[96]),
   .I1(InputBits[204]),
   .I2(InputBits[503]),
   .I3(InputBits[326]),
   .I4(InputBits[540]),
   .I5(InputBits[304])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000000000000010000001100110000000000110011)  
) LUT6_753 (
   .O(gates_753),
   .I0(InputBits[496]),
   .I1(InputBits[457]),
   .I2(InputBits[452]),
   .I3(InputBits[253]),
   .I4(InputBits[451]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0000000000000001010011000100010000110001010100010111110101110101)  
) LUT6_754 (
   .O(gates_754),
   .I0(InputBits[147]),
   .I1(InputBits[447]),
   .I2(InputBits[282]),
   .I3(InputBits[111]),
   .I4(InputBits[493]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000001000000000000000000000000000010010)  
) LUT6_755 (
   .O(gates_755),
   .I0(InputBits[8]),
   .I1(InputBits[555]),
   .I2(InputBits[66]),
   .I3(InputBits[48]),
   .I4(InputBits[546]),
   .I5(InputBits[257])
);
LUT6 #(
   .INIT(64'b0000000000000000010100010001000100000000000000001000101101111111)  
) LUT6_756 (
   .O(gates_756),
   .I0(InputBits[503]),
   .I1(InputBits[59]),
   .I2(InputBits[173]),
   .I3(InputBits[183]),
   .I4(InputBits[146]),
   .I5(InputBits[243])
);
LUT6 #(
   .INIT(64'b0111001111110010111101111111111101011010010110001111101111111011)  
) LUT6_757 (
   .O(gates_757),
   .I0(InputBits[140]),
   .I1(InputBits[173]),
   .I2(InputBits[422]),
   .I3(InputBits[357]),
   .I4(InputBits[81]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0000001001000001010001101100111100000010010001001100111011001111)  
) LUT6_758 (
   .O(gates_758),
   .I0(InputBits[447]),
   .I1(InputBits[417]),
   .I2(InputBits[512]),
   .I3(InputBits[544]),
   .I4(InputBits[274]),
   .I5(InputBits[197])
);
LUT6 #(
   .INIT(64'b0101000100000010100101101000000001110001011101110101010111010100)  
) LUT6_759 (
   .O(gates_759),
   .I0(InputBits[570]),
   .I1(InputBits[137]),
   .I2(InputBits[161]),
   .I3(InputBits[244]),
   .I4(InputBits[345]),
   .I5(InputBits[277])
);
LUT6 #(
   .INIT(64'b0000000000100001001000000000000101111101011101111111001111111111)  
) LUT6_760 (
   .O(gates_760),
   .I0(InputBits[113]),
   .I1(InputBits[432]),
   .I2(InputBits[453]),
   .I3(InputBits[490]),
   .I4(InputBits[257]),
   .I5(InputBits[517])
);
LUT6 #(
   .INIT(64'b1011111111101101001100110011001111110111101111011111001011111011)  
) LUT6_761 (
   .O(gates_761),
   .I0(InputBits[88]),
   .I1(InputBits[489]),
   .I2(InputBits[113]),
   .I3(InputBits[428]),
   .I4(InputBits[478]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1011101011111111111110110011001110101011101010101011001100100000)  
) LUT6_762 (
   .O(gates_762),
   .I0(InputBits[223]),
   .I1(InputBits[231]),
   .I2(InputBits[309]),
   .I3(InputBits[292]),
   .I4(InputBits[295]),
   .I5(InputBits[366])
);
LUT6 #(
   .INIT(64'b0000010001110101010001000100010100100101111111110110000001100111)  
) LUT6_763 (
   .O(gates_763),
   .I0(InputBits[526]),
   .I1(InputBits[202]),
   .I2(InputBits[110]),
   .I3(InputBits[494]),
   .I4(InputBits[326]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0000000000010011000000000000000000000000000100010000000010001011)  
) LUT6_764 (
   .O(gates_764),
   .I0(InputBits[90]),
   .I1(InputBits[452]),
   .I2(InputBits[131]),
   .I3(InputBits[362]),
   .I4(InputBits[119]),
   .I5(InputBits[534])
);
LUT6 #(
   .INIT(64'b0000000010000000000000000000001100000010001100111010001011111111)  
) LUT6_765 (
   .O(gates_765),
   .I0(InputBits[203]),
   .I1(InputBits[207]),
   .I2(InputBits[485]),
   .I3(InputBits[511]),
   .I4(InputBits[281]),
   .I5(InputBits[362])
);
LUT6 #(
   .INIT(64'b0000000001010101000000000100010000000000010000010000010001000100)  
) LUT6_766 (
   .O(gates_766),
   .I0(InputBits[552]),
   .I1(InputBits[234]),
   .I2(InputBits[57]),
   .I3(InputBits[543]),
   .I4(InputBits[324]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0000000000000000000010000100011100001111000011001100110111001111)  
) LUT6_767 (
   .O(gates_767),
   .I0(InputBits[184]),
   .I1(InputBits[345]),
   .I2(InputBits[472]),
   .I3(InputBits[282]),
   .I4(InputBits[565]),
   .I5(InputBits[216])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110000001100010011000000011101)  
) LUT6_768 (
   .O(gates_768),
   .I0(InputBits[486]),
   .I1(InputBits[534]),
   .I2(InputBits[359]),
   .I3(InputBits[108]),
   .I4(InputBits[137]),
   .I5(InputBits[457])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100110000000000000000)  
) LUT6_769 (
   .O(gates_769),
   .I0(InputBits[497]),
   .I1(InputBits[575]),
   .I2(InputBits[314]),
   .I3(InputBits[131]),
   .I4(InputBits[350]),
   .I5(InputBits[555])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000001010000011100000101000001110)  
) LUT6_770 (
   .O(gates_770),
   .I0(InputBits[342]),
   .I1(InputBits[268]),
   .I2(InputBits[146]),
   .I3(InputBits[523]),
   .I4(InputBits[197]),
   .I5(InputBits[41])
);
LUT6 #(
   .INIT(64'b0100110100001101010011100100101000000111000000110001011100000010)  
) LUT6_771 (
   .O(gates_771),
   .I0(InputBits[311]),
   .I1(InputBits[281]),
   .I2(InputBits[144]),
   .I3(InputBits[369]),
   .I4(InputBits[317]),
   .I5(InputBits[305])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000111100000000000000000000001100001100)  
) LUT6_772 (
   .O(gates_772),
   .I0(InputBits[467]),
   .I1(InputBits[311]),
   .I2(InputBits[50]),
   .I3(InputBits[526]),
   .I4(InputBits[313]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010111100000000000000000001001100100010)  
) LUT6_773 (
   .O(gates_773),
   .I0(InputBits[350]),
   .I1(InputBits[539]),
   .I2(InputBits[151]),
   .I3(InputBits[550]),
   .I4(InputBits[509]),
   .I5(InputBits[117])
);
LUT6 #(
   .INIT(64'b0101010101010101010100010101000101010100010100000000000000000000)  
) LUT6_774 (
   .O(gates_774),
   .I0(InputBits[123]),
   .I1(InputBits[115]),
   .I2(InputBits[176]),
   .I3(InputBits[307]),
   .I4(InputBits[272]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001110011001000110011011100110011)  
) LUT6_775 (
   .O(gates_775),
   .I0(InputBits[245]),
   .I1(InputBits[572]),
   .I2(InputBits[253]),
   .I3(InputBits[344]),
   .I4(InputBits[354]),
   .I5(InputBits[553])
);
LUT6 #(
   .INIT(64'b0001000000000000000101010001010000000000000001110001000000010100)  
) LUT6_776 (
   .O(gates_776),
   .I0(InputBits[172]),
   .I1(InputBits[248]),
   .I2(InputBits[12]),
   .I3(InputBits[35]),
   .I4(InputBits[412]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000010100000000)  
) LUT6_777 (
   .O(gates_777),
   .I0(InputBits[169]),
   .I1(InputBits[328]),
   .I2(InputBits[241]),
   .I3(InputBits[372]),
   .I4(InputBits[169]),
   .I5(InputBits[27])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011000000110000000100000001)  
) LUT6_778 (
   .O(gates_778),
   .I0(InputBits[378]),
   .I1(InputBits[72]),
   .I2(InputBits[82]),
   .I3(InputBits[543]),
   .I4(InputBits[202]),
   .I5(InputBits[26])
);
LUT6 #(
   .INIT(64'b0100010000000000010001000000000000000001000101010000000000000101)  
) LUT6_779 (
   .O(gates_779),
   .I0(InputBits[265]),
   .I1(InputBits[456]),
   .I2(InputBits[79]),
   .I3(InputBits[230]),
   .I4(InputBits[343]),
   .I5(InputBits[254])
);
LUT6 #(
   .INIT(64'b0000100100011111000001010000111100000000000111110000000100000101)  
) LUT6_780 (
   .O(gates_780),
   .I0(InputBits[541]),
   .I1(InputBits[153]),
   .I2(InputBits[536]),
   .I3(InputBits[314]),
   .I4(InputBits[91]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000000000110001000000000011001100100001001100000000000100000000)  
) LUT6_781 (
   .O(gates_781),
   .I0(InputBits[174]),
   .I1(InputBits[28]),
   .I2(InputBits[245]),
   .I3(InputBits[526]),
   .I4(InputBits[258]),
   .I5(InputBits[237])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001101111100000000101111100000)  
) LUT6_782 (
   .O(gates_782),
   .I0(InputBits[153]),
   .I1(InputBits[413]),
   .I2(InputBits[293]),
   .I3(InputBits[502]),
   .I4(InputBits[375]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000010000000100010101010000000001010100)  
) LUT6_783 (
   .O(gates_783),
   .I0(InputBits[26]),
   .I1(InputBits[285]),
   .I2(InputBits[239]),
   .I3(InputBits[218]),
   .I4(InputBits[421]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000000100000001000000000000000100)  
) LUT6_784 (
   .O(gates_784),
   .I0(InputBits[169]),
   .I1(InputBits[177]),
   .I2(InputBits[482]),
   .I3(InputBits[156]),
   .I4(InputBits[438]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0001010001010101000000000000000101010101010101010101010101010101)  
) LUT6_785 (
   .O(gates_785),
   .I0(InputBits[145]),
   .I1(InputBits[390]),
   .I2(InputBits[226]),
   .I3(InputBits[232]),
   .I4(InputBits[323]),
   .I5(InputBits[254])
);
LUT6 #(
   .INIT(64'b0000000001010101001100100011001000000000111101110011101000111111)  
) LUT6_786 (
   .O(gates_786),
   .I0(InputBits[364]),
   .I1(InputBits[280]),
   .I2(InputBits[438]),
   .I3(InputBits[540]),
   .I4(InputBits[479]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000000000000001000000001)  
) LUT6_787 (
   .O(gates_787),
   .I0(InputBits[461]),
   .I1(InputBits[98]),
   .I2(InputBits[108]),
   .I3(InputBits[53]),
   .I4(InputBits[97]),
   .I5(InputBits[177])
);
LUT6 #(
   .INIT(64'b0010101100110111001010100010101000100011001110110010011000101111)  
) LUT6_788 (
   .O(gates_788),
   .I0(InputBits[261]),
   .I1(InputBits[40]),
   .I2(InputBits[539]),
   .I3(InputBits[485]),
   .I4(InputBits[166]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000100000000000000000000000100001110)  
) LUT6_789 (
   .O(gates_789),
   .I0(InputBits[39]),
   .I1(InputBits[12]),
   .I2(InputBits[98]),
   .I3(InputBits[339]),
   .I4(InputBits[481]),
   .I5(InputBits[94])
);
LUT6 #(
   .INIT(64'b0001010100010101010101000001000100010101000101010001000000010001)  
) LUT6_790 (
   .O(gates_790),
   .I0(InputBits[52]),
   .I1(InputBits[128]),
   .I2(InputBits[13]),
   .I3(InputBits[59]),
   .I4(InputBits[39]),
   .I5(InputBits[161])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001010000010100001110)  
) LUT6_791 (
   .O(gates_791),
   .I0(InputBits[40]),
   .I1(InputBits[430]),
   .I2(InputBits[28]),
   .I3(InputBits[339]),
   .I4(InputBits[548]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110011000000000001000100010000)  
) LUT6_792 (
   .O(gates_792),
   .I0(InputBits[462]),
   .I1(InputBits[146]),
   .I2(InputBits[445]),
   .I3(InputBits[291]),
   .I4(InputBits[136]),
   .I5(InputBits[572])
);
LUT6 #(
   .INIT(64'b0101010000010001010101000101010111111111000000011101011100110101)  
) LUT6_793 (
   .O(gates_793),
   .I0(InputBits[517]),
   .I1(InputBits[136]),
   .I2(InputBits[61]),
   .I3(InputBits[319]),
   .I4(InputBits[138]),
   .I5(InputBits[13])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000011100000111101)  
) LUT6_794 (
   .O(gates_794),
   .I0(InputBits[87]),
   .I1(InputBits[547]),
   .I2(InputBits[64]),
   .I3(InputBits[131]),
   .I4(InputBits[289]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010001111111110000000001010111)  
) LUT6_795 (
   .O(gates_795),
   .I0(InputBits[514]),
   .I1(InputBits[446]),
   .I2(InputBits[402]),
   .I3(InputBits[147]),
   .I4(InputBits[269]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0000000000000000001001010011011100000000000001001101010111111111)  
) LUT6_796 (
   .O(gates_796),
   .I0(InputBits[208]),
   .I1(InputBits[234]),
   .I2(InputBits[159]),
   .I3(InputBits[133]),
   .I4(InputBits[51]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000001000110011111100100011)  
) LUT6_797 (
   .O(gates_797),
   .I0(InputBits[399]),
   .I1(InputBits[515]),
   .I2(InputBits[474]),
   .I3(InputBits[93]),
   .I4(InputBits[16]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0011000100100000001100010001000000110011001100000011001100010000)  
) LUT6_798 (
   .O(gates_798),
   .I0(InputBits[405]),
   .I1(InputBits[555]),
   .I2(InputBits[261]),
   .I3(InputBits[341]),
   .I4(InputBits[136]),
   .I5(InputBits[150])
);
LUT6 #(
   .INIT(64'b0000000000110101000000001101111100000000000000000000010111001101)  
) LUT6_799 (
   .O(gates_799),
   .I0(InputBits[173]),
   .I1(InputBits[188]),
   .I2(InputBits[447]),
   .I3(InputBits[572]),
   .I4(InputBits[536]),
   .I5(InputBits[142])
);
LUT6 #(
   .INIT(64'b0000100011101111100011001110111100000000010000111010101011001110)  
) LUT6_800 (
   .O(gates_800),
   .I0(InputBits[269]),
   .I1(InputBits[236]),
   .I2(InputBits[112]),
   .I3(InputBits[149]),
   .I4(InputBits[93]),
   .I5(InputBits[165])
);
LUT6 #(
   .INIT(64'b0000000001110000011101000101000000100000001100001101111111111111)  
) LUT6_801 (
   .O(gates_801),
   .I0(InputBits[308]),
   .I1(InputBits[499]),
   .I2(InputBits[454]),
   .I3(InputBits[35]),
   .I4(InputBits[172]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0000001100000000000010110000110000110000000000001011111111001100)  
) LUT6_802 (
   .O(gates_802),
   .I0(InputBits[424]),
   .I1(InputBits[244]),
   .I2(InputBits[62]),
   .I3(InputBits[420]),
   .I4(InputBits[38]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0000000000000000010100010101000100000000000000000110011001000111)  
) LUT6_803 (
   .O(gates_803),
   .I0(InputBits[432]),
   .I1(InputBits[267]),
   .I2(InputBits[496]),
   .I3(InputBits[128]),
   .I4(InputBits[562]),
   .I5(InputBits[66])
);
LUT6 #(
   .INIT(64'b1111000000000000101011100000111101000000111001111010101010101110)  
) LUT6_804 (
   .O(gates_804),
   .I0(InputBits[371]),
   .I1(InputBits[259]),
   .I2(InputBits[174]),
   .I3(InputBits[464]),
   .I4(InputBits[220]),
   .I5(InputBits[179])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001111110100000000000101000000000110110001)  
) LUT6_805 (
   .O(gates_805),
   .I0(InputBits[148]),
   .I1(InputBits[101]),
   .I2(InputBits[316]),
   .I3(InputBits[16]),
   .I4(InputBits[458]),
   .I5(InputBits[198])
);
LUT6 #(
   .INIT(64'b0011001100110011001100100001000100110011001100110011000000010000)  
) LUT6_806 (
   .O(gates_806),
   .I0(InputBits[58]),
   .I1(InputBits[48]),
   .I2(InputBits[165]),
   .I3(InputBits[197]),
   .I4(InputBits[391]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0000000001000101000000000100110100000000000000000000000000000000)  
) LUT6_807 (
   .O(gates_807),
   .I0(InputBits[124]),
   .I1(InputBits[428]),
   .I2(InputBits[489]),
   .I3(InputBits[5]),
   .I4(InputBits[412]),
   .I5(InputBits[374])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001000000100000001110)  
) LUT6_808 (
   .O(gates_808),
   .I0(InputBits[369]),
   .I1(InputBits[394]),
   .I2(InputBits[97]),
   .I3(InputBits[148]),
   .I4(InputBits[535]),
   .I5(InputBits[555])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000100110000000000000011)  
) LUT6_809 (
   .O(gates_809),
   .I0(InputBits[205]),
   .I1(InputBits[564]),
   .I2(InputBits[509]),
   .I3(InputBits[557]),
   .I4(InputBits[480]),
   .I5(InputBits[38])
);
LUT6 #(
   .INIT(64'b0000000011111111001000011111101100000000111111110001001111111011)  
) LUT6_810 (
   .O(gates_810),
   .I0(InputBits[200]),
   .I1(InputBits[449]),
   .I2(InputBits[212]),
   .I3(InputBits[71]),
   .I4(InputBits[238]),
   .I5(InputBits[139])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000101000000000110101010101)  
) LUT6_811 (
   .O(gates_811),
   .I0(InputBits[207]),
   .I1(InputBits[181]),
   .I2(InputBits[8]),
   .I3(InputBits[412]),
   .I4(InputBits[231]),
   .I5(InputBits[147])
);
LUT6 #(
   .INIT(64'b0000110100001101000011110000111100001111000011110000111100000101)  
) LUT6_812 (
   .O(gates_812),
   .I0(InputBits[378]),
   .I1(InputBits[445]),
   .I2(InputBits[74]),
   .I3(InputBits[333]),
   .I4(InputBits[268]),
   .I5(InputBits[383])
);
LUT6 #(
   .INIT(64'b0000000000010001000000100011111100000000010111110000000000111111)  
) LUT6_813 (
   .O(gates_813),
   .I0(InputBits[222]),
   .I1(InputBits[79]),
   .I2(InputBits[227]),
   .I3(InputBits[532]),
   .I4(InputBits[479]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0000101100000011000010111010111100000010000000100000001000001010)  
) LUT6_814 (
   .O(gates_814),
   .I0(InputBits[342]),
   .I1(InputBits[104]),
   .I2(InputBits[172]),
   .I3(InputBits[93]),
   .I4(InputBits[302]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0000000000001010000011111110111000000000111100100000101011101110)  
) LUT6_815 (
   .O(gates_815),
   .I0(InputBits[372]),
   .I1(InputBits[200]),
   .I2(InputBits[546]),
   .I3(InputBits[37]),
   .I4(InputBits[172]),
   .I5(InputBits[153])
);
LUT6 #(
   .INIT(64'b0001000000010000000000000001000000010001000101010011001100000010)  
) LUT6_816 (
   .O(gates_816),
   .I0(InputBits[8]),
   .I1(InputBits[457]),
   .I2(InputBits[449]),
   .I3(InputBits[395]),
   .I4(InputBits[260]),
   .I5(InputBits[569])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010001000101010100)  
) LUT6_817 (
   .O(gates_817),
   .I0(InputBits[459]),
   .I1(InputBits[291]),
   .I2(InputBits[248]),
   .I3(InputBits[95]),
   .I4(InputBits[17]),
   .I5(InputBits[97])
);
LUT6 #(
   .INIT(64'b0000000000010001000100110000000000000000000000010001001100000110)  
) LUT6_818 (
   .O(gates_818),
   .I0(InputBits[67]),
   .I1(InputBits[13]),
   .I2(InputBits[55]),
   .I3(InputBits[501]),
   .I4(InputBits[311]),
   .I5(InputBits[469])
);
LUT6 #(
   .INIT(64'b0000000100000000000000101010101000000000000000000010001011101110)  
) LUT6_819 (
   .O(gates_819),
   .I0(InputBits[371]),
   .I1(InputBits[178]),
   .I2(InputBits[462]),
   .I3(InputBits[147]),
   .I4(InputBits[574]),
   .I5(InputBits[232])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000111110111111)  
) LUT6_820 (
   .O(gates_820),
   .I0(InputBits[304]),
   .I1(InputBits[95]),
   .I2(InputBits[105]),
   .I3(InputBits[274]),
   .I4(InputBits[18]),
   .I5(InputBits[552])
);
LUT6 #(
   .INIT(64'b0100000011001100001100010011000000000000110010000011000000110000)  
) LUT6_821 (
   .O(gates_821),
   .I0(InputBits[467]),
   .I1(InputBits[384]),
   .I2(InputBits[394]),
   .I3(InputBits[203]),
   .I4(InputBits[384]),
   .I5(InputBits[323])
);
LUT6 #(
   .INIT(64'b0111111111111111100100000101010011111111111111110000000100000100)  
) LUT6_822 (
   .O(gates_822),
   .I0(InputBits[58]),
   .I1(InputBits[158]),
   .I2(InputBits[498]),
   .I3(InputBits[327]),
   .I4(InputBits[392]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b0010000000110001001000000011000100100011000000110010001000110011)  
) LUT6_823 (
   .O(gates_823),
   .I0(InputBits[157]),
   .I1(InputBits[481]),
   .I2(InputBits[249]),
   .I3(InputBits[134]),
   .I4(InputBits[466]),
   .I5(InputBits[297])
);
LUT6 #(
   .INIT(64'b0000000100010000000100000001000101111111001100001111101111111100)  
) LUT6_824 (
   .O(gates_824),
   .I0(InputBits[151]),
   .I1(InputBits[546]),
   .I2(InputBits[398]),
   .I3(InputBits[391]),
   .I4(InputBits[405]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000000000000000100110011)  
) LUT6_825 (
   .O(gates_825),
   .I0(InputBits[451]),
   .I1(InputBits[505]),
   .I2(InputBits[33]),
   .I3(InputBits[518]),
   .I4(InputBits[457]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0000000000001000000000000000100000000000000000000000000000001001)  
) LUT6_826 (
   .O(gates_826),
   .I0(InputBits[451]),
   .I1(InputBits[425]),
   .I2(InputBits[99]),
   .I3(InputBits[509]),
   .I4(InputBits[426]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010100000000000000000000001111000011011000)  
) LUT6_827 (
   .O(gates_827),
   .I0(InputBits[63]),
   .I1(InputBits[157]),
   .I2(InputBits[247]),
   .I3(InputBits[440]),
   .I4(InputBits[145]),
   .I5(InputBits[534])
);
LUT6 #(
   .INIT(64'b0001000100010001000100010001000100000000000000000000000000010001)  
) LUT6_828 (
   .O(gates_828),
   .I0(InputBits[576]),
   .I1(InputBits[49]),
   .I2(InputBits[186]),
   .I3(InputBits[486]),
   .I4(InputBits[450]),
   .I5(InputBits[366])
);
LUT6 #(
   .INIT(64'b0000000010001101111100011000100000000000100011110101001111001101)  
) LUT6_829 (
   .O(gates_829),
   .I0(InputBits[450]),
   .I1(InputBits[188]),
   .I2(InputBits[437]),
   .I3(InputBits[215]),
   .I4(InputBits[339]),
   .I5(InputBits[109])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000100010001010100000101)  
) LUT6_830 (
   .O(gates_830),
   .I0(InputBits[265]),
   .I1(InputBits[435]),
   .I2(InputBits[513]),
   .I3(InputBits[357]),
   .I4(InputBits[479]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000011110110111101100110011111111111)  
) LUT6_831 (
   .O(gates_831),
   .I0(InputBits[92]),
   .I1(InputBits[335]),
   .I2(InputBits[176]),
   .I3(InputBits[197]),
   .I4(InputBits[463]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000000000100000000000001000000000000000111)  
) LUT6_832 (
   .O(gates_832),
   .I0(InputBits[483]),
   .I1(InputBits[6]),
   .I2(InputBits[171]),
   .I3(InputBits[560]),
   .I4(InputBits[277]),
   .I5(InputBits[510])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010001010101110000000100111011)  
) LUT6_833 (
   .O(gates_833),
   .I0(InputBits[522]),
   .I1(InputBits[509]),
   .I2(InputBits[273]),
   .I3(InputBits[403]),
   .I4(InputBits[94]),
   .I5(InputBits[218])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001100000001000000000000001100000001)  
) LUT6_834 (
   .O(gates_834),
   .I0(InputBits[113]),
   .I1(InputBits[49]),
   .I2(InputBits[22]),
   .I3(InputBits[91]),
   .I4(InputBits[134]),
   .I5(InputBits[562])
);
LUT6 #(
   .INIT(64'b0000000011111111000000001111001000000000111111110000000011111011)  
) LUT6_835 (
   .O(gates_835),
   .I0(InputBits[268]),
   .I1(InputBits[468]),
   .I2(InputBits[261]),
   .I3(InputBits[313]),
   .I4(InputBits[201]),
   .I5(InputBits[473])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000111100000011001010110000001110101011)  
) LUT6_836 (
   .O(gates_836),
   .I0(InputBits[399]),
   .I1(InputBits[100]),
   .I2(InputBits[55]),
   .I3(InputBits[13]),
   .I4(InputBits[388]),
   .I5(InputBits[547])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000100010000000110000001000001111)  
) LUT6_837 (
   .O(gates_837),
   .I0(InputBits[333]),
   .I1(InputBits[571]),
   .I2(InputBits[54]),
   .I3(InputBits[107]),
   .I4(InputBits[377]),
   .I5(InputBits[1])
);
LUT6 #(
   .INIT(64'b0010000011110101010100010101000100000000011101010101000001010001)  
) LUT6_838 (
   .O(gates_838),
   .I0(InputBits[252]),
   .I1(InputBits[102]),
   .I2(InputBits[423]),
   .I3(InputBits[30]),
   .I4(InputBits[382]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010000011011001101110011011000111000000100)  
) LUT6_839 (
   .O(gates_839),
   .I0(InputBits[79]),
   .I1(InputBits[350]),
   .I2(InputBits[124]),
   .I3(InputBits[422]),
   .I4(InputBits[165]),
   .I5(InputBits[240])
);
LUT6 #(
   .INIT(64'b0000000011011011000000001111101100000001111110110000000011001100)  
) LUT6_840 (
   .O(gates_840),
   .I0(InputBits[258]),
   .I1(InputBits[234]),
   .I2(InputBits[453]),
   .I3(InputBits[99]),
   .I4(InputBits[163]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0000000000000000110011110101111100000000000000001100010011010101)  
) LUT6_841 (
   .O(gates_841),
   .I0(InputBits[279]),
   .I1(InputBits[319]),
   .I2(InputBits[214]),
   .I3(InputBits[302]),
   .I4(InputBits[74]),
   .I5(InputBits[349])
);
LUT6 #(
   .INIT(64'b0000000001010101000100000100000000000000010101010001010100010000)  
) LUT6_842 (
   .O(gates_842),
   .I0(InputBits[21]),
   .I1(InputBits[138]),
   .I2(InputBits[181]),
   .I3(InputBits[408]),
   .I4(InputBits[190]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0000000000101001000000001000111000000000001101110000000010101111)  
) LUT6_843 (
   .O(gates_843),
   .I0(InputBits[444]),
   .I1(InputBits[199]),
   .I2(InputBits[205]),
   .I3(InputBits[409]),
   .I4(InputBits[288]),
   .I5(InputBits[425])
);
LUT6 #(
   .INIT(64'b0101000011111110000101101000111001010101101111100101111111011111)  
) LUT6_844 (
   .O(gates_844),
   .I0(InputBits[429]),
   .I1(InputBits[333]),
   .I2(InputBits[476]),
   .I3(InputBits[307]),
   .I4(InputBits[449]),
   .I5(InputBits[128])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000000000101000000000000000100110011)  
) LUT6_845 (
   .O(gates_845),
   .I0(InputBits[504]),
   .I1(InputBits[75]),
   .I2(InputBits[301]),
   .I3(InputBits[235]),
   .I4(InputBits[354]),
   .I5(InputBits[574])
);
LUT6 #(
   .INIT(64'b0000000000001111000000000000101000000000000011110000000000111010)  
) LUT6_846 (
   .O(gates_846),
   .I0(InputBits[370]),
   .I1(InputBits[469]),
   .I2(InputBits[96]),
   .I3(InputBits[27]),
   .I4(InputBits[408]),
   .I5(InputBits[138])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000011001100000000001000000011001100110000)  
) LUT6_847 (
   .O(gates_847),
   .I0(InputBits[381]),
   .I1(InputBits[531]),
   .I2(InputBits[419]),
   .I3(InputBits[288]),
   .I4(InputBits[434]),
   .I5(InputBits[215])
);
LUT6 #(
   .INIT(64'b0100111101011100010011000100100001000111010111110000000001000011)  
) LUT6_848 (
   .O(gates_848),
   .I0(InputBits[197]),
   .I1(InputBits[375]),
   .I2(InputBits[44]),
   .I3(InputBits[258]),
   .I4(InputBits[344]),
   .I5(InputBits[329])
);
LUT6 #(
   .INIT(64'b0000000000000000001000110011111100000000000000000001011110111111)  
) LUT6_849 (
   .O(gates_849),
   .I0(InputBits[477]),
   .I1(InputBits[100]),
   .I2(InputBits[515]),
   .I3(InputBits[277]),
   .I4(InputBits[49]),
   .I5(InputBits[84])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000001000000000001010100000101)  
) LUT6_850 (
   .O(gates_850),
   .I0(InputBits[19]),
   .I1(InputBits[282]),
   .I2(InputBits[512]),
   .I3(InputBits[64]),
   .I4(InputBits[490]),
   .I5(InputBits[123])
);
LUT6 #(
   .INIT(64'b0000000011111111000000001111010100000000111100000000000011100000)  
) LUT6_851 (
   .O(gates_851),
   .I0(InputBits[497]),
   .I1(InputBits[333]),
   .I2(InputBits[292]),
   .I3(InputBits[26]),
   .I4(InputBits[177]),
   .I5(InputBits[294])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000011100000000010100000000000001111011)  
) LUT6_852 (
   .O(gates_852),
   .I0(InputBits[323]),
   .I1(InputBits[486]),
   .I2(InputBits[155]),
   .I3(InputBits[574]),
   .I4(InputBits[517]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011101111111111111011111110101110)  
) LUT6_853 (
   .O(gates_853),
   .I0(InputBits[189]),
   .I1(InputBits[445]),
   .I2(InputBits[424]),
   .I3(InputBits[442]),
   .I4(InputBits[238]),
   .I5(InputBits[385])
);
LUT6 #(
   .INIT(64'b0001111000001010000011110000101000101111101110100011011100111011)  
) LUT6_854 (
   .O(gates_854),
   .I0(InputBits[292]),
   .I1(InputBits[83]),
   .I2(InputBits[546]),
   .I3(InputBits[416]),
   .I4(InputBits[151]),
   .I5(InputBits[487])
);
LUT6 #(
   .INIT(64'b0000001000000000000000100000000011111111111100101111011110111010)  
) LUT6_855 (
   .O(gates_855),
   .I0(InputBits[67]),
   .I1(InputBits[249]),
   .I2(InputBits[308]),
   .I3(InputBits[422]),
   .I4(InputBits[157]),
   .I5(InputBits[482])
);
LUT6 #(
   .INIT(64'b0000010101000101000001010000000000000001000101010000010100000111)  
) LUT6_856 (
   .O(gates_856),
   .I0(InputBits[20]),
   .I1(InputBits[136]),
   .I2(InputBits[52]),
   .I3(InputBits[143]),
   .I4(InputBits[212]),
   .I5(InputBits[487])
);
LUT6 #(
   .INIT(64'b0000000000000000000100100001001001000101000000010001001100010011)  
) LUT6_857 (
   .O(gates_857),
   .I0(InputBits[13]),
   .I1(InputBits[75]),
   .I2(InputBits[42]),
   .I3(InputBits[452]),
   .I4(InputBits[196]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010001000100010000000000010010001000110011)  
) LUT6_858 (
   .O(gates_858),
   .I0(InputBits[360]),
   .I1(InputBits[555]),
   .I2(InputBits[228]),
   .I3(InputBits[251]),
   .I4(InputBits[16]),
   .I5(InputBits[479])
);
LUT6 #(
   .INIT(64'b0000000000110010000100000011001000000000001100000000000000110000)  
) LUT6_859 (
   .O(gates_859),
   .I0(InputBits[39]),
   .I1(InputBits[2]),
   .I2(InputBits[367]),
   .I3(InputBits[75]),
   .I4(InputBits[86]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0000000100100111000001010010011000001000000011100000000000001111)  
) LUT6_860 (
   .O(gates_860),
   .I0(InputBits[381]),
   .I1(InputBits[332]),
   .I2(InputBits[410]),
   .I3(InputBits[566]),
   .I4(InputBits[297]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000000000000000010100000100010000000000000000000101011101000101)  
) LUT6_861 (
   .O(gates_861),
   .I0(InputBits[124]),
   .I1(InputBits[201]),
   .I2(InputBits[130]),
   .I3(InputBits[524]),
   .I4(InputBits[47]),
   .I5(InputBits[435])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110001000100000000000000010111011100010001)  
) LUT6_862 (
   .O(gates_862),
   .I0(InputBits[489]),
   .I1(InputBits[104]),
   .I2(InputBits[135]),
   .I3(InputBits[294]),
   .I4(InputBits[18]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0101000100000000010101010101010101010101000000000101010101000111)  
) LUT6_863 (
   .O(gates_863),
   .I0(InputBits[5]),
   .I1(InputBits[220]),
   .I2(InputBits[449]),
   .I3(InputBits[394]),
   .I4(InputBits[231]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0000000100000000001000010000000100110011001111110010001100100111)  
) LUT6_864 (
   .O(gates_864),
   .I0(InputBits[57]),
   .I1(InputBits[16]),
   .I2(InputBits[128]),
   .I3(InputBits[154]),
   .I4(InputBits[439]),
   .I5(InputBits[493])
);
LUT6 #(
   .INIT(64'b0000000000111100000101010101111110001100000011010101110101001111)  
) LUT6_865 (
   .O(gates_865),
   .I0(InputBits[517]),
   .I1(InputBits[319]),
   .I2(InputBits[53]),
   .I3(InputBits[403]),
   .I4(InputBits[516]),
   .I5(InputBits[327])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000000000000000000001111110000000100111100)  
) LUT6_866 (
   .O(gates_866),
   .I0(InputBits[461]),
   .I1(InputBits[549]),
   .I2(InputBits[191]),
   .I3(InputBits[7]),
   .I4(InputBits[212]),
   .I5(InputBits[564])
);
LUT6 #(
   .INIT(64'b0000000000000000000010110000110000000000000000100000101100000010)  
) LUT6_867 (
   .O(gates_867),
   .I0(InputBits[91]),
   .I1(InputBits[209]),
   .I2(InputBits[53]),
   .I3(InputBits[44]),
   .I4(InputBits[175]),
   .I5(InputBits[45])
);
LUT6 #(
   .INIT(64'b0000111000001110000011100010111000000110010111110101111000101110)  
) LUT6_868 (
   .O(gates_868),
   .I0(InputBits[237]),
   .I1(InputBits[373]),
   .I2(InputBits[216]),
   .I3(InputBits[227]),
   .I4(InputBits[176]),
   .I5(InputBits[132])
);
LUT6 #(
   .INIT(64'b0000000000110111011100000111010100000001111101010111010001110101)  
) LUT6_869 (
   .O(gates_869),
   .I0(InputBits[254]),
   .I1(InputBits[468]),
   .I2(InputBits[222]),
   .I3(InputBits[125]),
   .I4(InputBits[363]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1000000010000010110000001100001010000000110000100000000011000011)  
) LUT6_870 (
   .O(gates_870),
   .I0(InputBits[444]),
   .I1(InputBits[430]),
   .I2(InputBits[430]),
   .I3(InputBits[509]),
   .I4(InputBits[150]),
   .I5(InputBits[488])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000010111000001110)  
) LUT6_871 (
   .O(gates_871),
   .I0(InputBits[245]),
   .I1(InputBits[407]),
   .I2(InputBits[123]),
   .I3(InputBits[220]),
   .I4(InputBits[386]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0011000100110001000100000011000100110001001100110001000100110001)  
) LUT6_872 (
   .O(gates_872),
   .I0(InputBits[275]),
   .I1(InputBits[47]),
   .I2(InputBits[341]),
   .I3(InputBits[492]),
   .I4(InputBits[294]),
   .I5(InputBits[227])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011111111111011111011111100001010)  
) LUT6_873 (
   .O(gates_873),
   .I0(InputBits[260]),
   .I1(InputBits[165]),
   .I2(InputBits[153]),
   .I3(InputBits[420]),
   .I4(InputBits[177]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1010101011101010100010101010101000101011001011100010101111111111)  
) LUT6_874 (
   .O(gates_874),
   .I0(InputBits[416]),
   .I1(InputBits[176]),
   .I2(InputBits[523]),
   .I3(InputBits[157]),
   .I4(InputBits[486]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0000000000000000010101010000000000010001000100010101010100000111)  
) LUT6_875 (
   .O(gates_875),
   .I0(InputBits[290]),
   .I1(InputBits[64]),
   .I2(InputBits[513]),
   .I3(InputBits[418]),
   .I4(InputBits[119]),
   .I5(InputBits[77])
);
LUT6 #(
   .INIT(64'b0000000000000110000000110001001100001000000001110000111100010011)  
) LUT6_876 (
   .O(gates_876),
   .I0(InputBits[521]),
   .I1(InputBits[128]),
   .I2(InputBits[8]),
   .I3(InputBits[94]),
   .I4(InputBits[243]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100000000000000011000000110000001000100010)  
) LUT6_877 (
   .O(gates_877),
   .I0(InputBits[341]),
   .I1(InputBits[551]),
   .I2(InputBits[264]),
   .I3(InputBits[235]),
   .I4(InputBits[479]),
   .I5(InputBits[563])
);
LUT6 #(
   .INIT(64'b0000000100000011000000010001011100000001000000000000000101000101)  
) LUT6_878 (
   .O(gates_878),
   .I0(InputBits[483]),
   .I1(InputBits[314]),
   .I2(InputBits[147]),
   .I3(InputBits[408]),
   .I4(InputBits[107]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0000000011011111000000001101110111010001010101010101000001010101)  
) LUT6_879 (
   .O(gates_879),
   .I0(InputBits[275]),
   .I1(InputBits[211]),
   .I2(InputBits[89]),
   .I3(InputBits[16]),
   .I4(InputBits[446]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0000000000110111000000000111010100000000000100010000000000110011)  
) LUT6_880 (
   .O(gates_880),
   .I0(InputBits[204]),
   .I1(InputBits[434]),
   .I2(InputBits[40]),
   .I3(InputBits[533]),
   .I4(InputBits[34]),
   .I5(InputBits[451])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010000000000000000000010000000100100010)  
) LUT6_881 (
   .O(gates_881),
   .I0(InputBits[569]),
   .I1(InputBits[552]),
   .I2(InputBits[568]),
   .I3(InputBits[551]),
   .I4(InputBits[90]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000010100000000000001010000000000011111)  
) LUT6_882 (
   .O(gates_882),
   .I0(InputBits[537]),
   .I1(InputBits[160]),
   .I2(InputBits[557]),
   .I3(InputBits[105]),
   .I4(InputBits[469]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0000010000000100111111110000000001000001000100010111111110100010)  
) LUT6_883 (
   .O(gates_883),
   .I0(InputBits[260]),
   .I1(InputBits[280]),
   .I2(InputBits[452]),
   .I3(InputBits[370]),
   .I4(InputBits[12]),
   .I5(InputBits[257])
);
LUT6 #(
   .INIT(64'b0000010000000000000000000000010100000000000101000011001100110111)  
) LUT6_884 (
   .O(gates_884),
   .I0(InputBits[412]),
   .I1(InputBits[240]),
   .I2(InputBits[66]),
   .I3(InputBits[437]),
   .I4(InputBits[208]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0000000000000000111100001101000000000000000000000000000000001011)  
) LUT6_885 (
   .O(gates_885),
   .I0(InputBits[87]),
   .I1(InputBits[499]),
   .I2(InputBits[376]),
   .I3(InputBits[171]),
   .I4(InputBits[22]),
   .I5(InputBits[376])
);
LUT6 #(
   .INIT(64'b0000000000110011000000010011001100110001001101110011001100110001)  
) LUT6_886 (
   .O(gates_886),
   .I0(InputBits[80]),
   .I1(InputBits[386]),
   .I2(InputBits[197]),
   .I3(InputBits[287]),
   .I4(InputBits[477]),
   .I5(InputBits[92])
);
LUT6 #(
   .INIT(64'b0001000000000000000000000010100011011101110011001111110111110100)  
) LUT6_887 (
   .O(gates_887),
   .I0(InputBits[257]),
   .I1(InputBits[421]),
   .I2(InputBits[370]),
   .I3(InputBits[333]),
   .I4(InputBits[539]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0000000001000101000000000100010000000000010101000000000001000100)  
) LUT6_888 (
   .O(gates_888),
   .I0(InputBits[554]),
   .I1(InputBits[236]),
   .I2(InputBits[116]),
   .I3(InputBits[170]),
   .I4(InputBits[93]),
   .I5(InputBits[466])
);
LUT6 #(
   .INIT(64'b0001001100000011001100010011000100000011000000110111000100111011)  
) LUT6_889 (
   .O(gates_889),
   .I0(InputBits[109]),
   .I1(InputBits[51]),
   .I2(InputBits[478]),
   .I3(InputBits[330]),
   .I4(InputBits[335]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000101100000000000000010000000000110011)  
) LUT6_890 (
   .O(gates_890),
   .I0(InputBits[380]),
   .I1(InputBits[536]),
   .I2(InputBits[570]),
   .I3(InputBits[562]),
   .I4(InputBits[77]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0101010101010001010111110101000000010101010100010101110100000000)  
) LUT6_891 (
   .O(gates_891),
   .I0(InputBits[503]),
   .I1(InputBits[448]),
   .I2(InputBits[225]),
   .I3(InputBits[373]),
   .I4(InputBits[66]),
   .I5(InputBits[161])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000000000000000000000001)  
) LUT6_892 (
   .O(gates_892),
   .I0(InputBits[535]),
   .I1(InputBits[2]),
   .I2(InputBits[433]),
   .I3(InputBits[552]),
   .I4(InputBits[513]),
   .I5(InputBits[158])
);
LUT6 #(
   .INIT(64'b0000000000010001000000000011000000000000001100010000000011010000)  
) LUT6_893 (
   .O(gates_893),
   .I0(InputBits[257]),
   .I1(InputBits[172]),
   .I2(InputBits[444]),
   .I3(InputBits[571]),
   .I4(InputBits[239]),
   .I5(InputBits[451])
);
LUT6 #(
   .INIT(64'b0000000000000000000100110000000000000000000100010000000000010010)  
) LUT6_894 (
   .O(gates_894),
   .I0(InputBits[95]),
   .I1(InputBits[51]),
   .I2(InputBits[239]),
   .I3(InputBits[199]),
   .I4(InputBits[31]),
   .I5(InputBits[199])
);
LUT6 #(
   .INIT(64'b0001000011110000000000001111000000000100000010100000000000001110)  
) LUT6_895 (
   .O(gates_895),
   .I0(InputBits[262]),
   .I1(InputBits[292]),
   .I2(InputBits[270]),
   .I3(InputBits[434]),
   .I4(InputBits[388]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000100000100000001000100010001)  
) LUT6_896 (
   .O(gates_896),
   .I0(InputBits[171]),
   .I1(InputBits[53]),
   .I2(InputBits[339]),
   .I3(InputBits[327]),
   .I4(InputBits[509]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000000100010011)  
) LUT6_897 (
   .O(gates_897),
   .I0(InputBits[573]),
   .I1(InputBits[554]),
   .I2(InputBits[96]),
   .I3(InputBits[437]),
   .I4(InputBits[60]),
   .I5(InputBits[57])
);
LUT6 #(
   .INIT(64'b0001000101010101000001010001010100010001010101010000001101000101)  
) LUT6_898 (
   .O(gates_898),
   .I0(InputBits[572]),
   .I1(InputBits[226]),
   .I2(InputBits[463]),
   .I3(InputBits[523]),
   .I4(InputBits[441]),
   .I5(InputBits[244])
);
LUT6 #(
   .INIT(64'b0000000100110001000000010011001100000000001100010011000100110011)  
) LUT6_899 (
   .O(gates_899),
   .I0(InputBits[447]),
   .I1(InputBits[19]),
   .I2(InputBits[132]),
   .I3(InputBits[300]),
   .I4(InputBits[436]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001000100000001010000001001010100)  
) LUT6_900 (
   .O(gates_900),
   .I0(InputBits[507]),
   .I1(InputBits[41]),
   .I2(InputBits[386]),
   .I3(InputBits[411]),
   .I4(InputBits[211]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0000000000000011010100011111011100000000000000010000000111111101)  
) LUT6_901 (
   .O(gates_901),
   .I0(InputBits[515]),
   .I1(InputBits[191]),
   .I2(InputBits[142]),
   .I3(InputBits[43]),
   .I4(InputBits[524]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b0000000000000001000000010001000100000100000000010000010100000100)  
) LUT6_902 (
   .O(gates_902),
   .I0(InputBits[458]),
   .I1(InputBits[117]),
   .I2(InputBits[78]),
   .I3(InputBits[309]),
   .I4(InputBits[41]),
   .I5(InputBits[431])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100110000001010001111)  
) LUT6_903 (
   .O(gates_903),
   .I0(InputBits[499]),
   .I1(InputBits[503]),
   .I2(InputBits[497]),
   .I3(InputBits[338]),
   .I4(InputBits[357]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0000000000001111000000000000011100000000000011100000000000001000)  
) LUT6_904 (
   .O(gates_904),
   .I0(InputBits[198]),
   .I1(InputBits[466]),
   .I2(InputBits[337]),
   .I3(InputBits[73]),
   .I4(InputBits[164]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0000000000100001000000000010001000110011001100110011001100000001)  
) LUT6_905 (
   .O(gates_905),
   .I0(InputBits[305]),
   .I1(InputBits[313]),
   .I2(InputBits[353]),
   .I3(InputBits[69]),
   .I4(InputBits[368]),
   .I5(InputBits[547])
);
LUT6 #(
   .INIT(64'b0001001100000011000000010001001100010011000100110000000100010011)  
) LUT6_906 (
   .O(gates_906),
   .I0(InputBits[254]),
   .I1(InputBits[23]),
   .I2(InputBits[519]),
   .I3(InputBits[354]),
   .I4(InputBits[367]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0101010111010101011101010101010100100111101111110000001000100111)  
) LUT6_907 (
   .O(gates_907),
   .I0(InputBits[547]),
   .I1(InputBits[156]),
   .I2(InputBits[105]),
   .I3(InputBits[354]),
   .I4(InputBits[211]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0000000000000100000011010000110000000000000001010000110001011100)  
) LUT6_908 (
   .O(gates_908),
   .I0(InputBits[58]),
   .I1(InputBits[369]),
   .I2(InputBits[143]),
   .I3(InputBits[430]),
   .I4(InputBits[70]),
   .I5(InputBits[87])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110000000000000000000000000011001100000000)  
) LUT6_909 (
   .O(gates_909),
   .I0(InputBits[426]),
   .I1(InputBits[21]),
   .I2(InputBits[402]),
   .I3(InputBits[395]),
   .I4(InputBits[51]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010100000000000000000000010100000100)  
) LUT6_910 (
   .O(gates_910),
   .I0(InputBits[481]),
   .I1(InputBits[189]),
   .I2(InputBits[146]),
   .I3(InputBits[287]),
   .I4(InputBits[25]),
   .I5(InputBits[223])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000000000000000000000000000100010001010101)  
) LUT6_911 (
   .O(gates_911),
   .I0(InputBits[23]),
   .I1(InputBits[167]),
   .I2(InputBits[375]),
   .I3(InputBits[85]),
   .I4(InputBits[146]),
   .I5(InputBits[6])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010000000000000000000000000111100111110)  
) LUT6_912 (
   .O(gates_912),
   .I0(InputBits[442]),
   .I1(InputBits[70]),
   .I2(InputBits[480]),
   .I3(InputBits[166]),
   .I4(InputBits[242]),
   .I5(InputBits[54])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001010000000000000100)  
) LUT6_913 (
   .O(gates_913),
   .I0(InputBits[49]),
   .I1(InputBits[418]),
   .I2(InputBits[100]),
   .I3(InputBits[568]),
   .I4(InputBits[6]),
   .I5(InputBits[507])
);
LUT6 #(
   .INIT(64'b0000010100010101000001110001010100001111000010100001101100001000)  
) LUT6_914 (
   .O(gates_914),
   .I0(InputBits[43]),
   .I1(InputBits[484]),
   .I2(InputBits[194]),
   .I3(InputBits[398]),
   .I4(InputBits[429]),
   .I5(InputBits[316])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100100011001000010011000000100001)  
) LUT6_915 (
   .O(gates_915),
   .I0(InputBits[401]),
   .I1(InputBits[433]),
   .I2(InputBits[243]),
   .I3(InputBits[452]),
   .I4(InputBits[423]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0000000000110011000000001111001100000000101101100000000011111100)  
) LUT6_916 (
   .O(gates_916),
   .I0(InputBits[348]),
   .I1(InputBits[456]),
   .I2(InputBits[396]),
   .I3(InputBits[433]),
   .I4(InputBits[114]),
   .I5(InputBits[201])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000011000000000000000000000001000001110011)  
) LUT6_917 (
   .O(gates_917),
   .I0(InputBits[503]),
   .I1(InputBits[28]),
   .I2(InputBits[476]),
   .I3(InputBits[458]),
   .I4(InputBits[265]),
   .I5(InputBits[474])
);
LUT6 #(
   .INIT(64'b0101010101000000010000000000000001010101010101000101010000000000)  
) LUT6_918 (
   .O(gates_918),
   .I0(InputBits[47]),
   .I1(InputBits[351]),
   .I2(InputBits[398]),
   .I3(InputBits[224]),
   .I4(InputBits[367]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b0000111100101111000000111000011100101011110111110000000001111110)  
) LUT6_919 (
   .O(gates_919),
   .I0(InputBits[446]),
   .I1(InputBits[323]),
   .I2(InputBits[243]),
   .I3(InputBits[492]),
   .I4(InputBits[343]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0000000100000000000001010000001100000101000000010001000100000001)  
) LUT6_920 (
   .O(gates_920),
   .I0(InputBits[409]),
   .I1(InputBits[508]),
   .I2(InputBits[28]),
   .I3(InputBits[468]),
   .I4(InputBits[239]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000000001000010000000100000001000000010)  
) LUT6_921 (
   .O(gates_921),
   .I0(InputBits[237]),
   .I1(InputBits[281]),
   .I2(InputBits[42]),
   .I3(InputBits[187]),
   .I4(InputBits[40]),
   .I5(InputBits[144])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000111100000000000000000000111111110010)  
) LUT6_922 (
   .O(gates_922),
   .I0(InputBits[422]),
   .I1(InputBits[113]),
   .I2(InputBits[526]),
   .I3(InputBits[408]),
   .I4(InputBits[535]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000000000000000000000000000010100000011)  
) LUT6_923 (
   .O(gates_923),
   .I0(InputBits[195]),
   .I1(InputBits[536]),
   .I2(InputBits[1]),
   .I3(InputBits[200]),
   .I4(InputBits[253]),
   .I5(InputBits[128])
);
LUT6 #(
   .INIT(64'b0000000100000000010100010000000100010001000000000011000100000000)  
) LUT6_924 (
   .O(gates_924),
   .I0(InputBits[559]),
   .I1(InputBits[195]),
   .I2(InputBits[354]),
   .I3(InputBits[420]),
   .I4(InputBits[298]),
   .I5(InputBits[403])
);
LUT6 #(
   .INIT(64'b0001010100000000000000000000000100010000000100010010000101110001)  
) LUT6_925 (
   .O(gates_925),
   .I0(InputBits[30]),
   .I1(InputBits[538]),
   .I2(InputBits[468]),
   .I3(InputBits[487]),
   .I4(InputBits[267]),
   .I5(InputBits[512])
);
LUT6 #(
   .INIT(64'b0000000000010001000000001111001100000000000000010000000000000000)  
) LUT6_926 (
   .O(gates_926),
   .I0(InputBits[79]),
   .I1(InputBits[507]),
   .I2(InputBits[439]),
   .I3(InputBits[289]),
   .I4(InputBits[119]),
   .I5(InputBits[370])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100010001100000000000000000100001010110011)  
) LUT6_927 (
   .O(gates_927),
   .I0(InputBits[391]),
   .I1(InputBits[572]),
   .I2(InputBits[256]),
   .I3(InputBits[276]),
   .I4(InputBits[562]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000000000001111)  
) LUT6_928 (
   .O(gates_928),
   .I0(InputBits[485]),
   .I1(InputBits[504]),
   .I2(InputBits[147]),
   .I3(InputBits[529]),
   .I4(InputBits[492]),
   .I5(InputBits[541])
);
LUT6 #(
   .INIT(64'b1101111111010101111111111111111101001101000001010111011100110011)  
) LUT6_929 (
   .O(gates_929),
   .I0(InputBits[521]),
   .I1(InputBits[83]),
   .I2(InputBits[425]),
   .I3(InputBits[199]),
   .I4(InputBits[132]),
   .I5(InputBits[177])
);
LUT6 #(
   .INIT(64'b0000111100001011000000110000000000001111000010110000101000000010)  
) LUT6_930 (
   .O(gates_930),
   .I0(InputBits[444]),
   .I1(InputBits[84]),
   .I2(InputBits[558]),
   .I3(InputBits[350]),
   .I4(InputBits[319]),
   .I5(InputBits[115])
);
LUT6 #(
   .INIT(64'b0000000000110011000000000011001100000000101110111000100010101111)  
) LUT6_931 (
   .O(gates_931),
   .I0(InputBits[439]),
   .I1(InputBits[91]),
   .I2(InputBits[135]),
   .I3(InputBits[482]),
   .I4(InputBits[35]),
   .I5(InputBits[13])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100000001000000010001)  
) LUT6_932 (
   .O(gates_932),
   .I0(InputBits[98]),
   .I1(InputBits[253]),
   .I2(InputBits[346]),
   .I3(InputBits[361]),
   .I4(InputBits[75]),
   .I5(InputBits[170])
);
LUT6 #(
   .INIT(64'b0000101100001001101110111111101100001011000010111111001101111011)  
) LUT6_933 (
   .O(gates_933),
   .I0(InputBits[234]),
   .I1(InputBits[330]),
   .I2(InputBits[67]),
   .I3(InputBits[463]),
   .I4(InputBits[56]),
   .I5(InputBits[162])
);
LUT6 #(
   .INIT(64'b1011111110111111111111111011111110111010101110001011111110111111)  
) LUT6_934 (
   .O(gates_934),
   .I0(InputBits[285]),
   .I1(InputBits[308]),
   .I2(InputBits[382]),
   .I3(InputBits[62]),
   .I4(InputBits[105]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0000010100000101000001010000010100000000000000000000000100000001)  
) LUT6_935 (
   .O(gates_935),
   .I0(InputBits[529]),
   .I1(InputBits[110]),
   .I2(InputBits[49]),
   .I3(InputBits[439]),
   .I4(InputBits[459]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000010001000100001000100010001)  
) LUT6_936 (
   .O(gates_936),
   .I0(InputBits[282]),
   .I1(InputBits[552]),
   .I2(InputBits[290]),
   .I3(InputBits[571]),
   .I4(InputBits[353]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0000000000000100000010010000111100001101000011110000110000001111)  
) LUT6_937 (
   .O(gates_937),
   .I0(InputBits[111]),
   .I1(InputBits[373]),
   .I2(InputBits[4]),
   .I3(InputBits[230]),
   .I4(InputBits[165]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0011001100110011001100000011000000110011000000000011001100100011)  
) LUT6_938 (
   .O(gates_938),
   .I0(InputBits[116]),
   .I1(InputBits[2]),
   .I2(InputBits[473]),
   .I3(InputBits[177]),
   .I4(InputBits[471]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0011111100100111001111110011011100111111001110100011111100110110)  
) LUT6_939 (
   .O(gates_939),
   .I0(InputBits[334]),
   .I1(InputBits[67]),
   .I2(InputBits[335]),
   .I3(InputBits[343]),
   .I4(InputBits[423]),
   .I5(InputBits[373])
);
LUT6 #(
   .INIT(64'b0000001100010011010000011111001100000001000000111101011101010111)  
) LUT6_940 (
   .O(gates_940),
   .I0(InputBits[195]),
   .I1(InputBits[230]),
   .I2(InputBits[180]),
   .I3(InputBits[303]),
   .I4(InputBits[81]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000010101010000000001010101)  
) LUT6_941 (
   .O(gates_941),
   .I0(InputBits[537]),
   .I1(InputBits[138]),
   .I2(InputBits[62]),
   .I3(InputBits[218]),
   .I4(InputBits[65]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011000000100011000000010011)  
) LUT6_942 (
   .O(gates_942),
   .I0(InputBits[282]),
   .I1(InputBits[559]),
   .I2(InputBits[32]),
   .I3(InputBits[111]),
   .I4(InputBits[547]),
   .I5(InputBits[27])
);
LUT6 #(
   .INIT(64'b0011001100110011001100110010001000110011001101110000001100000011)  
) LUT6_943 (
   .O(gates_943),
   .I0(InputBits[399]),
   .I1(InputBits[557]),
   .I2(InputBits[84]),
   .I3(InputBits[66]),
   .I4(InputBits[371]),
   .I5(InputBits[498])
);
LUT6 #(
   .INIT(64'b0000101010111111001100111011101100100000001010100011101110111011)  
) LUT6_944 (
   .O(gates_944),
   .I0(InputBits[397]),
   .I1(InputBits[276]),
   .I2(InputBits[282]),
   .I3(InputBits[173]),
   .I4(InputBits[229]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0100000001000101110101010101010101000100000000000101000100000001)  
) LUT6_945 (
   .O(gates_945),
   .I0(InputBits[434]),
   .I1(InputBits[427]),
   .I2(InputBits[437]),
   .I3(InputBits[91]),
   .I4(InputBits[108]),
   .I5(InputBits[211])
);
LUT6 #(
   .INIT(64'b0000000001000000000000110000001110111111000000111111001100010011)  
) LUT6_946 (
   .O(gates_946),
   .I0(InputBits[451]),
   .I1(InputBits[491]),
   .I2(InputBits[132]),
   .I3(InputBits[389]),
   .I4(InputBits[151]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010001000000000000000000000001000100010000)  
) LUT6_947 (
   .O(gates_947),
   .I0(InputBits[505]),
   .I1(InputBits[532]),
   .I2(InputBits[418]),
   .I3(InputBits[118]),
   .I4(InputBits[575]),
   .I5(InputBits[375])
);
LUT6 #(
   .INIT(64'b0011001100110011001000100011001000110011001100110011001000110010)  
) LUT6_948 (
   .O(gates_948),
   .I0(InputBits[178]),
   .I1(InputBits[3]),
   .I2(InputBits[119]),
   .I3(InputBits[465]),
   .I4(InputBits[347]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0000001100000010000000110000000000000011000000010000001100000111)  
) LUT6_949 (
   .O(gates_949),
   .I0(InputBits[32]),
   .I1(InputBits[574]),
   .I2(InputBits[576]),
   .I3(InputBits[344]),
   .I4(InputBits[88]),
   .I5(InputBits[488])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000001000000001000110110000000100101011)  
) LUT6_950 (
   .O(gates_950),
   .I0(InputBits[142]),
   .I1(InputBits[106]),
   .I2(InputBits[565]),
   .I3(InputBits[571]),
   .I4(InputBits[332]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0011001100110011001000010011001100110111001101110010010000111111)  
) LUT6_951 (
   .O(gates_951),
   .I0(InputBits[185]),
   .I1(InputBits[119]),
   .I2(InputBits[430]),
   .I3(InputBits[105]),
   .I4(InputBits[421]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001000000001000000000011001100100010)  
) LUT6_952 (
   .O(gates_952),
   .I0(InputBits[341]),
   .I1(InputBits[146]),
   .I2(InputBits[520]),
   .I3(InputBits[287]),
   .I4(InputBits[561]),
   .I5(InputBits[99])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010001000000000000000100000001000100010001)  
) LUT6_953 (
   .O(gates_953),
   .I0(InputBits[53]),
   .I1(InputBits[98]),
   .I2(InputBits[244]),
   .I3(InputBits[439]),
   .I4(InputBits[571]),
   .I5(InputBits[133])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001100010000000000000000000000000011011111)  
) LUT6_954 (
   .O(gates_954),
   .I0(InputBits[519]),
   .I1(InputBits[157]),
   .I2(InputBits[414]),
   .I3(InputBits[337]),
   .I4(InputBits[123]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000001000100001001000110011001100110011001)  
) LUT6_955 (
   .O(gates_955),
   .I0(InputBits[280]),
   .I1(InputBits[280]),
   .I2(InputBits[222]),
   .I3(InputBits[448]),
   .I4(InputBits[503]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000011001000000000000000110001000000110000)  
) LUT6_956 (
   .O(gates_956),
   .I0(InputBits[203]),
   .I1(InputBits[386]),
   .I2(InputBits[268]),
   .I3(InputBits[242]),
   .I4(InputBits[14]),
   .I5(InputBits[165])
);
LUT6 #(
   .INIT(64'b0000000001101111000000001000111100000000101010110000000010101010)  
) LUT6_957 (
   .O(gates_957),
   .I0(InputBits[199]),
   .I1(InputBits[382]),
   .I2(InputBits[448]),
   .I3(InputBits[313]),
   .I4(InputBits[258]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0000000000000000101110111111111100110011001000001011001111111010)  
) LUT6_958 (
   .O(gates_958),
   .I0(InputBits[369]),
   .I1(InputBits[149]),
   .I2(InputBits[394]),
   .I3(InputBits[320]),
   .I4(InputBits[9]),
   .I5(InputBits[214])
);
LUT6 #(
   .INIT(64'b0000000100110011000000000000011000010001000100011010101100110111)  
) LUT6_959 (
   .O(gates_959),
   .I0(InputBits[90]),
   .I1(InputBits[17]),
   .I2(InputBits[473]),
   .I3(InputBits[328]),
   .I4(InputBits[432]),
   .I5(InputBits[299])
);
LUT6 #(
   .INIT(64'b0001001101010111000100110101111100000011000001000000000100001101)  
) LUT6_960 (
   .O(gates_960),
   .I0(InputBits[127]),
   .I1(InputBits[119]),
   .I2(InputBits[228]),
   .I3(InputBits[67]),
   .I4(InputBits[164]),
   .I5(InputBits[319])
);
LUT6 #(
   .INIT(64'b0101000101010001010100010101001100010000000100000101000100010011)  
) LUT6_961 (
   .O(gates_961),
   .I0(InputBits[168]),
   .I1(InputBits[253]),
   .I2(InputBits[310]),
   .I3(InputBits[186]),
   .I4(InputBits[133]),
   .I5(InputBits[179])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000100010000000100000000000000000001001110)  
) LUT6_962 (
   .O(gates_962),
   .I0(InputBits[119]),
   .I1(InputBits[319]),
   .I2(InputBits[90]),
   .I3(InputBits[172]),
   .I4(InputBits[76]),
   .I5(InputBits[161])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000001100000001)  
) LUT6_963 (
   .O(gates_963),
   .I0(InputBits[534]),
   .I1(InputBits[561]),
   .I2(InputBits[145]),
   .I3(InputBits[413]),
   .I4(InputBits[514]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000101010100000000010101010100000011000101)  
) LUT6_964 (
   .O(gates_964),
   .I0(InputBits[51]),
   .I1(InputBits[477]),
   .I2(InputBits[402]),
   .I3(InputBits[218]),
   .I4(InputBits[432]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0000000000010011001100010011001100000000001100110000000100000001)  
) LUT6_965 (
   .O(gates_965),
   .I0(InputBits[144]),
   .I1(InputBits[55]),
   .I2(InputBits[511]),
   .I3(InputBits[96]),
   .I4(InputBits[167]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1011111100101110111111110000110100110011001100111111111100111011)  
) LUT6_966 (
   .O(gates_966),
   .I0(InputBits[136]),
   .I1(InputBits[253]),
   .I2(InputBits[250]),
   .I3(InputBits[344]),
   .I4(InputBits[134]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b1101101011111000111100000101000011111000110111111111110011111110)  
) LUT6_967 (
   .O(gates_967),
   .I0(InputBits[64]),
   .I1(InputBits[224]),
   .I2(InputBits[365]),
   .I3(InputBits[380]),
   .I4(InputBits[179]),
   .I5(InputBits[488])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000000110001000000000001)  
) LUT6_968 (
   .O(gates_968),
   .I0(InputBits[280]),
   .I1(InputBits[531]),
   .I2(InputBits[51]),
   .I3(InputBits[147]),
   .I4(InputBits[46]),
   .I5(InputBits[175])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011000100000000001000000000110011101110)  
) LUT6_969 (
   .O(gates_969),
   .I0(InputBits[390]),
   .I1(InputBits[214]),
   .I2(InputBits[186]),
   .I3(InputBits[171]),
   .I4(InputBits[573]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000111000111111000111010001000)  
) LUT6_970 (
   .O(gates_970),
   .I0(InputBits[315]),
   .I1(InputBits[153]),
   .I2(InputBits[513]),
   .I3(InputBits[267]),
   .I4(InputBits[372]),
   .I5(InputBits[21])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001010101000000010101010000000000000000)  
) LUT6_971 (
   .O(gates_971),
   .I0(InputBits[49]),
   .I1(InputBits[138]),
   .I2(InputBits[404]),
   .I3(InputBits[53]),
   .I4(InputBits[286]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0100000100000100000001010101010101110111111101110111001101111111)  
) LUT6_972 (
   .O(gates_972),
   .I0(InputBits[473]),
   .I1(InputBits[336]),
   .I2(InputBits[111]),
   .I3(InputBits[226]),
   .I4(InputBits[328]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0000000000000000000011010000111100001100000001000000110100001101)  
) LUT6_973 (
   .O(gates_973),
   .I0(InputBits[108]),
   .I1(InputBits[389]),
   .I2(InputBits[529]),
   .I3(InputBits[65]),
   .I4(InputBits[482]),
   .I5(InputBits[334])
);
LUT6 #(
   .INIT(64'b0010001011110111111111111111111100000010010001000101111111010100)  
) LUT6_974 (
   .O(gates_974),
   .I0(InputBits[305]),
   .I1(InputBits[416]),
   .I2(InputBits[157]),
   .I3(InputBits[324]),
   .I4(InputBits[543]),
   .I5(InputBits[365])
);
LUT6 #(
   .INIT(64'b1101001000000010111100111011101111110011001000111100111011101111)  
) LUT6_975 (
   .O(gates_975),
   .I0(InputBits[258]),
   .I1(InputBits[180]),
   .I2(InputBits[131]),
   .I3(InputBits[438]),
   .I4(InputBits[475]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0011000000110001001000010011001111101100111111010011111111111111)  
) LUT6_976 (
   .O(gates_976),
   .I0(InputBits[438]),
   .I1(InputBits[287]),
   .I2(InputBits[222]),
   .I3(InputBits[512]),
   .I4(InputBits[492]),
   .I5(InputBits[291])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000000000000000000000101010000000000000000)  
) LUT6_977 (
   .O(gates_977),
   .I0(InputBits[528]),
   .I1(InputBits[129]),
   .I2(InputBits[227]),
   .I3(InputBits[532]),
   .I4(InputBits[395]),
   .I5(InputBits[482])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000100000111000000010101011101)  
) LUT6_978 (
   .O(gates_978),
   .I0(InputBits[124]),
   .I1(InputBits[395]),
   .I2(InputBits[215]),
   .I3(InputBits[387]),
   .I4(InputBits[84]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0000001000100000001100111111001000010011001100010011001100110001)  
) LUT6_979 (
   .O(gates_979),
   .I0(InputBits[328]),
   .I1(InputBits[29]),
   .I2(InputBits[370]),
   .I3(InputBits[43]),
   .I4(InputBits[206]),
   .I5(InputBits[281])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100111111100000000000000010000000101110000)  
) LUT6_980 (
   .O(gates_980),
   .I0(InputBits[416]),
   .I1(InputBits[519]),
   .I2(InputBits[118]),
   .I3(InputBits[9]),
   .I4(InputBits[216]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001111010000000001000000000000000011110000)  
) LUT6_981 (
   .O(gates_981),
   .I0(InputBits[499]),
   .I1(InputBits[332]),
   .I2(InputBits[260]),
   .I3(InputBits[571]),
   .I4(InputBits[571]),
   .I5(InputBits[352])
);
LUT6 #(
   .INIT(64'b0111001100010101001110100011001000111011001100010011101001111111)  
) LUT6_982 (
   .O(gates_982),
   .I0(InputBits[359]),
   .I1(InputBits[172]),
   .I2(InputBits[287]),
   .I3(InputBits[380]),
   .I4(InputBits[308]),
   .I5(InputBits[425])
);
LUT6 #(
   .INIT(64'b0000000000010001010000000010001000000001000100010000000000100010)  
) LUT6_983 (
   .O(gates_983),
   .I0(InputBits[261]),
   .I1(InputBits[31]),
   .I2(InputBits[88]),
   .I3(InputBits[77]),
   .I4(InputBits[432]),
   .I5(InputBits[161])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000000000000000100000001)  
) LUT6_984 (
   .O(gates_984),
   .I0(InputBits[86]),
   .I1(InputBits[122]),
   .I2(InputBits[313]),
   .I3(InputBits[573]),
   .I4(InputBits[559]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0000000100000011000000110000011100000000000000000000000100000001)  
) LUT6_985 (
   .O(gates_985),
   .I0(InputBits[54]),
   .I1(InputBits[338]),
   .I2(InputBits[265]),
   .I3(InputBits[357]),
   .I4(InputBits[512]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000001011000010110000001100001100)  
) LUT6_986 (
   .O(gates_986),
   .I0(InputBits[90]),
   .I1(InputBits[356]),
   .I2(InputBits[361]),
   .I3(InputBits[282]),
   .I4(InputBits[453]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1000011100000101100011110101110110111001010101011011111100100111)  
) LUT6_987 (
   .O(gates_987),
   .I0(InputBits[230]),
   .I1(InputBits[463]),
   .I2(InputBits[255]),
   .I3(InputBits[237]),
   .I4(InputBits[256]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000001000000000000010100000000000101010101)  
) LUT6_988 (
   .O(gates_988),
   .I0(InputBits[409]),
   .I1(InputBits[7]),
   .I2(InputBits[444]),
   .I3(InputBits[482]),
   .I4(InputBits[276]),
   .I5(InputBits[77])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000111100000000000000100000000011001111)  
) LUT6_989 (
   .O(gates_989),
   .I0(InputBits[445]),
   .I1(InputBits[186]),
   .I2(InputBits[81]),
   .I3(InputBits[533]),
   .I4(InputBits[279]),
   .I5(InputBits[387])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000001000010011000110110000)  
) LUT6_990 (
   .O(gates_990),
   .I0(InputBits[376]),
   .I1(InputBits[459]),
   .I2(InputBits[319]),
   .I3(InputBits[167]),
   .I4(InputBits[290]),
   .I5(InputBits[562])
);
LUT6 #(
   .INIT(64'b0000000010101111000100011111111100000000000011100000000010101111)  
) LUT6_991 (
   .O(gates_991),
   .I0(InputBits[262]),
   .I1(InputBits[334]),
   .I2(InputBits[104]),
   .I3(InputBits[434]),
   .I4(InputBits[536]),
   .I5(InputBits[366])
);
LUT6 #(
   .INIT(64'b0000001101000101010001010101111100010000000010100101000011001111)  
) LUT6_992 (
   .O(gates_992),
   .I0(InputBits[143]),
   .I1(InputBits[379]),
   .I2(InputBits[380]),
   .I3(InputBits[449]),
   .I4(InputBits[128]),
   .I5(InputBits[283])
);
LUT6 #(
   .INIT(64'b1110101001111111110000001111000111111010111110111111101011111011)  
) LUT6_993 (
   .O(gates_993),
   .I0(InputBits[247]),
   .I1(InputBits[377]),
   .I2(InputBits[390]),
   .I3(InputBits[355]),
   .I4(InputBits[234]),
   .I5(InputBits[452])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000100000000010001)  
) LUT6_994 (
   .O(gates_994),
   .I0(InputBits[450]),
   .I1(InputBits[425]),
   .I2(InputBits[120]),
   .I3(InputBits[400]),
   .I4(InputBits[48]),
   .I5(InputBits[82])
);
LUT6 #(
   .INIT(64'b0000000000000000000011110001111100000000000000000000000000000001)  
) LUT6_995 (
   .O(gates_995),
   .I0(InputBits[461]),
   .I1(InputBits[80]),
   .I2(InputBits[266]),
   .I3(InputBits[132]),
   .I4(InputBits[555]),
   .I5(InputBits[342])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000001001100110011000100010001)  
) LUT6_996 (
   .O(gates_996),
   .I0(InputBits[275]),
   .I1(InputBits[48]),
   .I2(InputBits[234]),
   .I3(InputBits[44]),
   .I4(InputBits[285]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0000001100011111000000110001101100000111000100110000001101010000)  
) LUT6_997 (
   .O(gates_997),
   .I0(InputBits[65]),
   .I1(InputBits[509]),
   .I2(InputBits[120]),
   .I3(InputBits[407]),
   .I4(InputBits[397]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000101100001100010011111000111111)  
) LUT6_998 (
   .O(gates_998),
   .I0(InputBits[439]),
   .I1(InputBits[32]),
   .I2(InputBits[291]),
   .I3(InputBits[132]),
   .I4(InputBits[206]),
   .I5(InputBits[74])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000000000000010001000000011110111011101111)  
) LUT6_999 (
   .O(gates_999),
   .I0(InputBits[214]),
   .I1(InputBits[270]),
   .I2(InputBits[84]),
   .I3(InputBits[60]),
   .I4(InputBits[11]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0101010101010101001001000100111100010101010101010000000001011111)  
) LUT6_1000 (
   .O(gates_1000),
   .I0(InputBits[384]),
   .I1(InputBits[422]),
   .I2(InputBits[498]),
   .I3(InputBits[515]),
   .I4(InputBits[165]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000100010000000000110011)  
) LUT6_1001 (
   .O(gates_1001),
   .I0(InputBits[304]),
   .I1(InputBits[576]),
   .I2(InputBits[415]),
   .I3(InputBits[145]),
   .I4(InputBits[230]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000000000110001001100110111001100000000001101010011000100110001)  
) LUT6_1002 (
   .O(gates_1002),
   .I0(InputBits[471]),
   .I1(InputBits[560]),
   .I2(InputBits[222]),
   .I3(InputBits[65]),
   .I4(InputBits[143]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0001010100010101010101010101010100000001000100000000000100010001)  
) LUT6_1003 (
   .O(gates_1003),
   .I0(InputBits[122]),
   .I1(InputBits[101]),
   .I2(InputBits[248]),
   .I3(InputBits[476]),
   .I4(InputBits[112]),
   .I5(InputBits[244])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010100000000000001110000001000000010)  
) LUT6_1004 (
   .O(gates_1004),
   .I0(InputBits[144]),
   .I1(InputBits[63]),
   .I2(InputBits[361]),
   .I3(InputBits[301]),
   .I4(InputBits[141]),
   .I5(InputBits[455])
);
LUT6 #(
   .INIT(64'b1100010111001101100000010101111111101111101011100101110110101011)  
) LUT6_1005 (
   .O(gates_1005),
   .I0(InputBits[478]),
   .I1(InputBits[234]),
   .I2(InputBits[403]),
   .I3(InputBits[201]),
   .I4(InputBits[327]),
   .I5(InputBits[524])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000000000010000000001010101)  
) LUT6_1006 (
   .O(gates_1006),
   .I0(InputBits[483]),
   .I1(InputBits[196]),
   .I2(InputBits[545]),
   .I3(InputBits[540]),
   .I4(InputBits[29]),
   .I5(InputBits[57])
);
LUT6 #(
   .INIT(64'b0011000100000011000000000001000000110001001101010011000100111111)  
) LUT6_1007 (
   .O(gates_1007),
   .I0(InputBits[302]),
   .I1(InputBits[17]),
   .I2(InputBits[271]),
   .I3(InputBits[353]),
   .I4(InputBits[387]),
   .I5(InputBits[434])
);
LUT6 #(
   .INIT(64'b1101000111110101000100010011010100110011111101110001001111110011)  
) LUT6_1008 (
   .O(gates_1008),
   .I0(InputBits[173]),
   .I1(InputBits[83]),
   .I2(InputBits[465]),
   .I3(InputBits[273]),
   .I4(InputBits[164]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000110010001111)  
) LUT6_1009 (
   .O(gates_1009),
   .I0(InputBits[296]),
   .I1(InputBits[320]),
   .I2(InputBits[493]),
   .I3(InputBits[133]),
   .I4(InputBits[17]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0000000001010101000000001111000000000000110111110000000010110000)  
) LUT6_1010 (
   .O(gates_1010),
   .I0(InputBits[175]),
   .I1(InputBits[114]),
   .I2(InputBits[164]),
   .I3(InputBits[21]),
   .I4(InputBits[191]),
   .I5(InputBits[181])
);
LUT6 #(
   .INIT(64'b0000000100001111000000010000111100000001000000000000100000001000)  
) LUT6_1011 (
   .O(gates_1011),
   .I0(InputBits[336]),
   .I1(InputBits[107]),
   .I2(InputBits[28]),
   .I3(InputBits[517]),
   .I4(InputBits[422]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1010001011100011010000001111111101010000000100000011000011110000)  
) LUT6_1012 (
   .O(gates_1012),
   .I0(InputBits[476]),
   .I1(InputBits[332]),
   .I2(InputBits[294]),
   .I3(InputBits[171]),
   .I4(InputBits[100]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0000000000000000000101010000010000000000000000000101010101000101)  
) LUT6_1013 (
   .O(gates_1013),
   .I0(InputBits[554]),
   .I1(InputBits[44]),
   .I2(InputBits[434]),
   .I3(InputBits[391]),
   .I4(InputBits[97]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000000000000001011110011001100000000000000011111111100000001)  
) LUT6_1014 (
   .O(gates_1014),
   .I0(InputBits[112]),
   .I1(InputBits[158]),
   .I2(InputBits[486]),
   .I3(InputBits[366]),
   .I4(InputBits[561]),
   .I5(InputBits[523])
);
LUT6 #(
   .INIT(64'b0000000000000000001100110011001100110000000100100011011100111111)  
) LUT6_1015 (
   .O(gates_1015),
   .I0(InputBits[91]),
   .I1(InputBits[216]),
   .I2(InputBits[364]),
   .I3(InputBits[139]),
   .I4(InputBits[539]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110111110111001111111111001111)  
) LUT6_1016 (
   .O(gates_1016),
   .I0(InputBits[158]),
   .I1(InputBits[310]),
   .I2(InputBits[297]),
   .I3(InputBits[190]),
   .I4(InputBits[328]),
   .I5(InputBits[99])
);
LUT6 #(
   .INIT(64'b0001000101010000000100000001010100000000010001110001010100000001)  
) LUT6_1017 (
   .O(gates_1017),
   .I0(InputBits[565]),
   .I1(InputBits[380]),
   .I2(InputBits[160]),
   .I3(InputBits[480]),
   .I4(InputBits[210]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b0000000100000100000000100000001000000101000001000000100000001100)  
) LUT6_1018 (
   .O(gates_1018),
   .I0(InputBits[35]),
   .I1(InputBits[163]),
   .I2(InputBits[146]),
   .I3(InputBits[114]),
   .I4(InputBits[203]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000000001000000000000000000000000000001111)  
) LUT6_1019 (
   .O(gates_1019),
   .I0(InputBits[202]),
   .I1(InputBits[301]),
   .I2(InputBits[313]),
   .I3(InputBits[48]),
   .I4(InputBits[107]),
   .I5(InputBits[132])
);
LUT6 #(
   .INIT(64'b0011001100110011001100110011001100110011001000110000001100100000)  
) LUT6_1020 (
   .O(gates_1020),
   .I0(InputBits[418]),
   .I1(InputBits[572]),
   .I2(InputBits[325]),
   .I3(InputBits[237]),
   .I4(InputBits[344]),
   .I5(InputBits[294])
);
LUT6 #(
   .INIT(64'b0000000000000000010011100000001100000000000000001110111111111111)  
) LUT6_1021 (
   .O(gates_1021),
   .I0(InputBits[157]),
   .I1(InputBits[437]),
   .I2(InputBits[487]),
   .I3(InputBits[191]),
   .I4(InputBits[27]),
   .I5(InputBits[277])
);
LUT6 #(
   .INIT(64'b0000000000000000000100110001001100000101010001010001011101011111)  
) LUT6_1022 (
   .O(gates_1022),
   .I0(InputBits[516]),
   .I1(InputBits[428]),
   .I2(InputBits[231]),
   .I3(InputBits[249]),
   .I4(InputBits[37]),
   .I5(InputBits[119])
);
LUT6 #(
   .INIT(64'b0000000000000000001111110001001100000000001101001111101100111011)  
) LUT6_1023 (
   .O(gates_1023),
   .I0(InputBits[414]),
   .I1(InputBits[275]),
   .I2(InputBits[302]),
   .I3(InputBits[285]),
   .I4(InputBits[527]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010111000101010000010001000111)  
) LUT6_1024 (
   .O(gates_1024),
   .I0(InputBits[572]),
   .I1(InputBits[166]),
   .I2(InputBits[80]),
   .I3(InputBits[299]),
   .I4(InputBits[364]),
   .I5(InputBits[19])
);
LUT6 #(
   .INIT(64'b0100110000001010010011110000111100001011000010110000111100000011)  
) LUT6_1025 (
   .O(gates_1025),
   .I0(InputBits[63]),
   .I1(InputBits[330]),
   .I2(InputBits[99]),
   .I3(InputBits[165]),
   .I4(InputBits[430]),
   .I5(InputBits[308])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000111000000000000000110000000000001111)  
) LUT6_1026 (
   .O(gates_1026),
   .I0(InputBits[318]),
   .I1(InputBits[30]),
   .I2(InputBits[253]),
   .I3(InputBits[552]),
   .I4(InputBits[264]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0001000100010001010101010101000100010001000100010001000000010000)  
) LUT6_1027 (
   .O(gates_1027),
   .I0(InputBits[22]),
   .I1(InputBits[386]),
   .I2(InputBits[340]),
   .I3(InputBits[141]),
   .I4(InputBits[221]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b0000000000001110000000000000111100000000000010100000010100001111)  
) LUT6_1028 (
   .O(gates_1028),
   .I0(InputBits[310]),
   .I1(InputBits[165]),
   .I2(InputBits[433]),
   .I3(InputBits[571]),
   .I4(InputBits[83]),
   .I5(InputBits[375])
);
LUT6 #(
   .INIT(64'b0000010000000000000001010000010100000000000000000000000100000101)  
) LUT6_1029 (
   .O(gates_1029),
   .I0(InputBits[97]),
   .I1(InputBits[358]),
   .I2(InputBits[576]),
   .I3(InputBits[300]),
   .I4(InputBits[276]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0000100000000010111110101111111000100000000010001111101011111010)  
) LUT6_1030 (
   .O(gates_1030),
   .I0(InputBits[396]),
   .I1(InputBits[419]),
   .I2(InputBits[260]),
   .I3(InputBits[425]),
   .I4(InputBits[75]),
   .I5(InputBits[184])
);
LUT6 #(
   .INIT(64'b0101000101110101011100110111011101010001010101010100010001010101)  
) LUT6_1031 (
   .O(gates_1031),
   .I0(InputBits[509]),
   .I1(InputBits[34]),
   .I2(InputBits[466]),
   .I3(InputBits[127]),
   .I4(InputBits[234]),
   .I5(InputBits[365])
);
LUT6 #(
   .INIT(64'b0000001000000010000100100001011100010010000101100001000000010101)  
) LUT6_1032 (
   .O(gates_1032),
   .I0(InputBits[34]),
   .I1(InputBits[168]),
   .I2(InputBits[263]),
   .I3(InputBits[83]),
   .I4(InputBits[475]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0001001100000011001100110011001100000011000000110000001100000011)  
) LUT6_1033 (
   .O(gates_1033),
   .I0(InputBits[140]),
   .I1(InputBits[19]),
   .I2(InputBits[253]),
   .I3(InputBits[204]),
   .I4(InputBits[221]),
   .I5(InputBits[349])
);
LUT6 #(
   .INIT(64'b0000010100000000011101010000000011101111101011101111111110101111)  
) LUT6_1034 (
   .O(gates_1034),
   .I0(InputBits[317]),
   .I1(InputBits[444]),
   .I2(InputBits[485]),
   .I3(InputBits[260]),
   .I4(InputBits[109]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000100000000000000110000000000000010)  
) LUT6_1035 (
   .O(gates_1035),
   .I0(InputBits[527]),
   .I1(InputBits[558]),
   .I2(InputBits[52]),
   .I3(InputBits[1]),
   .I4(InputBits[294]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000000011000000101000001110)  
) LUT6_1036 (
   .O(gates_1036),
   .I0(InputBits[65]),
   .I1(InputBits[248]),
   .I2(InputBits[553]),
   .I3(InputBits[60]),
   .I4(InputBits[184]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0001000100010001000000000001000101010001110101010000000000110001)  
) LUT6_1037 (
   .O(gates_1037),
   .I0(InputBits[124]),
   .I1(InputBits[79]),
   .I2(InputBits[114]),
   .I3(InputBits[508]),
   .I4(InputBits[439]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b0000000000000010010000110001011100000000001100010000110101001111)  
) LUT6_1038 (
   .O(gates_1038),
   .I0(InputBits[330]),
   .I1(InputBits[226]),
   .I2(InputBits[516]),
   .I3(InputBits[387]),
   .I4(InputBits[550]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000111001000000000000000000101110011111111)  
) LUT6_1039 (
   .O(gates_1039),
   .I0(InputBits[267]),
   .I1(InputBits[158]),
   .I2(InputBits[326]),
   .I3(InputBits[228]),
   .I4(InputBits[74]),
   .I5(InputBits[100])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101000000010000000000000101)  
) LUT6_1040 (
   .O(gates_1040),
   .I0(InputBits[194]),
   .I1(InputBits[412]),
   .I2(InputBits[553]),
   .I3(InputBits[231]),
   .I4(InputBits[243]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b0000000000010001000000100001000110111111111101110000000000010001)  
) LUT6_1041 (
   .O(gates_1041),
   .I0(InputBits[425]),
   .I1(InputBits[536]),
   .I2(InputBits[273]),
   .I3(InputBits[426]),
   .I4(InputBits[317]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b0000001000001111000000100000111100000010000000000000001100001100)  
) LUT6_1042 (
   .O(gates_1042),
   .I0(InputBits[441]),
   .I1(InputBits[308]),
   .I2(InputBits[559]),
   .I3(InputBits[15]),
   .I4(InputBits[234]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b0001000100010001000001010000010000010001000100010101011101010100)  
) LUT6_1043 (
   .O(gates_1043),
   .I0(InputBits[99]),
   .I1(InputBits[339]),
   .I2(InputBits[88]),
   .I3(InputBits[421]),
   .I4(InputBits[525]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000001011100000000000001000000000001001111)  
) LUT6_1044 (
   .O(gates_1044),
   .I0(InputBits[267]),
   .I1(InputBits[437]),
   .I2(InputBits[564]),
   .I3(InputBits[553]),
   .I4(InputBits[507]),
   .I5(InputBits[375])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000011111111111111111011001111111111)  
) LUT6_1045 (
   .O(gates_1045),
   .I0(InputBits[365]),
   .I1(InputBits[108]),
   .I2(InputBits[390]),
   .I3(InputBits[513]),
   .I4(InputBits[236]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000110011001111110011001000000000)  
) LUT6_1046 (
   .O(gates_1046),
   .I0(InputBits[423]),
   .I1(InputBits[539]),
   .I2(InputBits[62]),
   .I3(InputBits[501]),
   .I4(InputBits[342]),
   .I5(InputBits[26])
);
LUT6 #(
   .INIT(64'b0000000000000000010000101110111100011011000011011011101111111111)  
) LUT6_1047 (
   .O(gates_1047),
   .I0(InputBits[160]),
   .I1(InputBits[428]),
   .I2(InputBits[303]),
   .I3(InputBits[226]),
   .I4(InputBits[493]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0000000000000000000011100101111100000000000000000000111100000001)  
) LUT6_1048 (
   .O(gates_1048),
   .I0(InputBits[450]),
   .I1(InputBits[424]),
   .I2(InputBits[565]),
   .I3(InputBits[431]),
   .I4(InputBits[337]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1111110111111110111111001111111101010100011100000101110001110000)  
) LUT6_1049 (
   .O(gates_1049),
   .I0(InputBits[496]),
   .I1(InputBits[224]),
   .I2(InputBits[238]),
   .I3(InputBits[295]),
   .I4(InputBits[165]),
   .I5(InputBits[294])
);
LUT6 #(
   .INIT(64'b0000000000000000111100111111101100000000000000001110001011110000)  
) LUT6_1050 (
   .O(gates_1050),
   .I0(InputBits[423]),
   .I1(InputBits[327]),
   .I2(InputBits[369]),
   .I3(InputBits[357]),
   .I4(InputBits[563]),
   .I5(InputBits[199])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100000001100001110101010110000111110111111)  
) LUT6_1051 (
   .O(gates_1051),
   .I0(InputBits[417]),
   .I1(InputBits[106]),
   .I2(InputBits[512]),
   .I3(InputBits[36]),
   .I4(InputBits[279]),
   .I5(InputBits[362])
);
LUT6 #(
   .INIT(64'b0000000010100010101000111011101100000010000011110010011100101111)  
) LUT6_1052 (
   .O(gates_1052),
   .I0(InputBits[444]),
   .I1(InputBits[510]),
   .I2(InputBits[83]),
   .I3(InputBits[256]),
   .I4(InputBits[513]),
   .I5(InputBits[152])
);
LUT6 #(
   .INIT(64'b0000000000001100000000111110111100000000100011000000010111001111)  
) LUT6_1053 (
   .O(gates_1053),
   .I0(InputBits[59]),
   .I1(InputBits[348]),
   .I2(InputBits[78]),
   .I3(InputBits[314]),
   .I4(InputBits[275]),
   .I5(InputBits[467])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000010001000000000000000000001000000010001)  
) LUT6_1054 (
   .O(gates_1054),
   .I0(InputBits[34]),
   .I1(InputBits[48]),
   .I2(InputBits[394]),
   .I3(InputBits[279]),
   .I4(InputBits[555]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0000000100000000000000010011001100000011000000100000001100110011)  
) LUT6_1055 (
   .O(gates_1055),
   .I0(InputBits[292]),
   .I1(InputBits[72]),
   .I2(InputBits[279]),
   .I3(InputBits[438]),
   .I4(InputBits[512]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010001000100110001010100000001)  
) LUT6_1056 (
   .O(gates_1056),
   .I0(InputBits[566]),
   .I1(InputBits[534]),
   .I2(InputBits[82]),
   .I3(InputBits[359]),
   .I4(InputBits[320]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0000000000001000101111110100110000001100000011001111111101011100)  
) LUT6_1057 (
   .O(gates_1057),
   .I0(InputBits[282]),
   .I1(InputBits[246]),
   .I2(InputBits[406]),
   .I3(InputBits[373]),
   .I4(InputBits[567]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000111111100000000000000010000000000000011)  
) LUT6_1058 (
   .O(gates_1058),
   .I0(InputBits[387]),
   .I1(InputBits[106]),
   .I2(InputBits[488]),
   .I3(InputBits[558]),
   .I4(InputBits[528]),
   .I5(InputBits[419])
);
LUT6 #(
   .INIT(64'b0011001100110011000100110001001100100011001100110000001100000011)  
) LUT6_1059 (
   .O(gates_1059),
   .I0(InputBits[322]),
   .I1(InputBits[481]),
   .I2(InputBits[494]),
   .I3(InputBits[468]),
   .I4(InputBits[142]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010100000000000000000101010100000000)  
) LUT6_1060 (
   .O(gates_1060),
   .I0(InputBits[50]),
   .I1(InputBits[127]),
   .I2(InputBits[148]),
   .I3(InputBits[397]),
   .I4(InputBits[193]),
   .I5(InputBits[69])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000001010000000000000000)  
) LUT6_1061 (
   .O(gates_1061),
   .I0(InputBits[194]),
   .I1(InputBits[89]),
   .I2(InputBits[554]),
   .I3(InputBits[196]),
   .I4(InputBits[263]),
   .I5(InputBits[119])
);
LUT6 #(
   .INIT(64'b0000000000000000001100111111111100000000000100001011001010111011)  
) LUT6_1062 (
   .O(gates_1062),
   .I0(InputBits[270]),
   .I1(InputBits[276]),
   .I2(InputBits[163]),
   .I3(InputBits[496]),
   .I4(InputBits[28]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000000111100001111)  
) LUT6_1063 (
   .O(gates_1063),
   .I0(InputBits[351]),
   .I1(InputBits[519]),
   .I2(InputBits[47]),
   .I3(InputBits[138]),
   .I4(InputBits[251]),
   .I5(InputBits[553])
);
LUT6 #(
   .INIT(64'b0100000001000100000000000110010100000000010001000000000001101010)  
) LUT6_1064 (
   .O(gates_1064),
   .I0(InputBits[549]),
   .I1(InputBits[284]),
   .I2(InputBits[187]),
   .I3(InputBits[386]),
   .I4(InputBits[400]),
   .I5(InputBits[90])
);
LUT6 #(
   .INIT(64'b0000010100000000000000000000000000000000000000111101010101010011)  
) LUT6_1065 (
   .O(gates_1065),
   .I0(InputBits[112]),
   .I1(InputBits[299]),
   .I2(InputBits[144]),
   .I3(InputBits[281]),
   .I4(InputBits[451]),
   .I5(InputBits[218])
);
LUT6 #(
   .INIT(64'b0010000101100100000001110011001101100110011001000110011101110111)  
) LUT6_1066 (
   .O(gates_1066),
   .I0(InputBits[165]),
   .I1(InputBits[384]),
   .I2(InputBits[158]),
   .I3(InputBits[352]),
   .I4(InputBits[251]),
   .I5(InputBits[197])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001001100000000000001010000000000000011)  
) LUT6_1067 (
   .O(gates_1067),
   .I0(InputBits[105]),
   .I1(InputBits[275]),
   .I2(InputBits[564]),
   .I3(InputBits[575]),
   .I4(InputBits[571]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0000000100000101000001010000010100000001000000010000000000000001)  
) LUT6_1068 (
   .O(gates_1068),
   .I0(InputBits[75]),
   .I1(InputBits[127]),
   .I2(InputBits[552]),
   .I3(InputBits[489]),
   .I4(InputBits[202]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0101010100010101010001010100010000010101010001110101010001000110)  
) LUT6_1069 (
   .O(gates_1069),
   .I0(InputBits[10]),
   .I1(InputBits[334]),
   .I2(InputBits[544]),
   .I3(InputBits[225]),
   .I4(InputBits[397]),
   .I5(InputBits[179])
);
LUT6 #(
   .INIT(64'b0000000000001111000000000000010100000000000011100000000001011110)  
) LUT6_1070 (
   .O(gates_1070),
   .I0(InputBits[201]),
   .I1(InputBits[431]),
   .I2(InputBits[16]),
   .I3(InputBits[409]),
   .I4(InputBits[177]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010100000000000000000111011101001110)  
) LUT6_1071 (
   .O(gates_1071),
   .I0(InputBits[479]),
   .I1(InputBits[284]),
   .I2(InputBits[38]),
   .I3(InputBits[396]),
   .I4(InputBits[26]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0000000000000000111100001100000000001011000011111111110011111100)  
) LUT6_1072 (
   .O(gates_1072),
   .I0(InputBits[209]),
   .I1(InputBits[319]),
   .I2(InputBits[244]),
   .I3(InputBits[466]),
   .I4(InputBits[13]),
   .I5(InputBits[128])
);
LUT6 #(
   .INIT(64'b0101011101000100010001010100011001000111000001100100011100000110)  
) LUT6_1073 (
   .O(gates_1073),
   .I0(InputBits[14]),
   .I1(InputBits[223]),
   .I2(InputBits[498]),
   .I3(InputBits[319]),
   .I4(InputBits[234]),
   .I5(InputBits[115])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000111110000000000000100010000000000101010)  
) LUT6_1074 (
   .O(gates_1074),
   .I0(InputBits[92]),
   .I1(InputBits[249]),
   .I2(InputBits[452]),
   .I3(InputBits[21]),
   .I4(InputBits[527]),
   .I5(InputBits[164])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000011001000000000000000010011001100110000)  
) LUT6_1075 (
   .O(gates_1075),
   .I0(InputBits[157]),
   .I1(InputBits[362]),
   .I2(InputBits[421]),
   .I3(InputBits[432]),
   .I4(InputBits[551]),
   .I5(InputBits[7])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000000001000001010000000100000001)  
) LUT6_1076 (
   .O(gates_1076),
   .I0(InputBits[385]),
   .I1(InputBits[483]),
   .I2(InputBits[74]),
   .I3(InputBits[71]),
   .I4(InputBits[180]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0100000000000000010101010100010000000100000000000001000100000001)  
) LUT6_1077 (
   .O(gates_1077),
   .I0(InputBits[146]),
   .I1(InputBits[59]),
   .I2(InputBits[426]),
   .I3(InputBits[140]),
   .I4(InputBits[362]),
   .I5(InputBits[152])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010100000000000000000000000000000101)  
) LUT6_1078 (
   .O(gates_1078),
   .I0(InputBits[253]),
   .I1(InputBits[322]),
   .I2(InputBits[97]),
   .I3(InputBits[2]),
   .I4(InputBits[217]),
   .I5(InputBits[438])
);
LUT6 #(
   .INIT(64'b0001000101110111000100000011001100000001000000100000000001110111)  
) LUT6_1079 (
   .O(gates_1079),
   .I0(InputBits[287]),
   .I1(InputBits[411]),
   .I2(InputBits[164]),
   .I3(InputBits[570]),
   .I4(InputBits[305]),
   .I5(InputBits[258])
);
LUT6 #(
   .INIT(64'b0000000000000000000101010001010100000000000000000001001100011111)  
) LUT6_1080 (
   .O(gates_1080),
   .I0(InputBits[94]),
   .I1(InputBits[250]),
   .I2(InputBits[124]),
   .I3(InputBits[79]),
   .I4(InputBits[241]),
   .I5(InputBits[478])
);
LUT6 #(
   .INIT(64'b0000000000000000001100010011000100000000000000000011000100010000)  
) LUT6_1081 (
   .O(gates_1081),
   .I0(InputBits[299]),
   .I1(InputBits[409]),
   .I2(InputBits[344]),
   .I3(InputBits[247]),
   .I4(InputBits[532]),
   .I5(InputBits[359])
);
LUT6 #(
   .INIT(64'b0000010010101110000001101010111110110101101010101111111110101110)  
) LUT6_1082 (
   .O(gates_1082),
   .I0(InputBits[373]),
   .I1(InputBits[389]),
   .I2(InputBits[329]),
   .I3(InputBits[335]),
   .I4(InputBits[490]),
   .I5(InputBits[139])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000000000000000000010100010000)  
) LUT6_1083 (
   .O(gates_1083),
   .I0(InputBits[122]),
   .I1(InputBits[568]),
   .I2(InputBits[290]),
   .I3(InputBits[270]),
   .I4(InputBits[229]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010000000000001011)  
) LUT6_1084 (
   .O(gates_1084),
   .I0(InputBits[227]),
   .I1(InputBits[558]),
   .I2(InputBits[52]),
   .I3(InputBits[402]),
   .I4(InputBits[175]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000000000000000000000110001001100110011)  
) LUT6_1085 (
   .O(gates_1085),
   .I0(InputBits[163]),
   .I1(InputBits[217]),
   .I2(InputBits[88]),
   .I3(InputBits[360]),
   .I4(InputBits[95]),
   .I5(InputBits[534])
);
LUT6 #(
   .INIT(64'b0000000011111111000000011011111100001011101011111100111110101111)  
) LUT6_1086 (
   .O(gates_1086),
   .I0(InputBits[371]),
   .I1(InputBits[333]),
   .I2(InputBits[254]),
   .I3(InputBits[143]),
   .I4(InputBits[181]),
   .I5(InputBits[383])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000100000001000101010000000000)  
) LUT6_1087 (
   .O(gates_1087),
   .I0(InputBits[529]),
   .I1(InputBits[350]),
   .I2(InputBits[173]),
   .I3(InputBits[398]),
   .I4(InputBits[41]),
   .I5(InputBits[74])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000100001110110011110000111001101110)  
) LUT6_1088 (
   .O(gates_1088),
   .I0(InputBits[359]),
   .I1(InputBits[222]),
   .I2(InputBits[100]),
   .I3(InputBits[60]),
   .I4(InputBits[271]),
   .I5(InputBits[504])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010100000101000101010100010100)  
) LUT6_1089 (
   .O(gates_1089),
   .I0(InputBits[4]),
   .I1(InputBits[213]),
   .I2(InputBits[70]),
   .I3(InputBits[422]),
   .I4(InputBits[491]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0000000000110011000000000011101100000000000000000000000000100011)  
) LUT6_1090 (
   .O(gates_1090),
   .I0(InputBits[211]),
   .I1(InputBits[508]),
   .I2(InputBits[447]),
   .I3(InputBits[48]),
   .I4(InputBits[103]),
   .I5(InputBits[335])
);
LUT6 #(
   .INIT(64'b0000000011111111000000000100000100000000110111110000000001000101)  
) LUT6_1091 (
   .O(gates_1091),
   .I0(InputBits[130]),
   .I1(InputBits[249]),
   .I2(InputBits[377]),
   .I3(InputBits[72]),
   .I4(InputBits[199]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0001000000001000010101110101111110000000010111010100000011101111)  
) LUT6_1092 (
   .O(gates_1092),
   .I0(InputBits[463]),
   .I1(InputBits[163]),
   .I2(InputBits[547]),
   .I3(InputBits[279]),
   .I4(InputBits[82]),
   .I5(InputBits[326])
);
LUT6 #(
   .INIT(64'b1001110000001000000011010000000011111111010010101010101110001010)  
) LUT6_1093 (
   .O(gates_1093),
   .I0(InputBits[523]),
   .I1(InputBits[114]),
   .I2(InputBits[427]),
   .I3(InputBits[345]),
   .I4(InputBits[415]),
   .I5(InputBits[520])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001111111100000000100100110000000011011111)  
) LUT6_1094 (
   .O(gates_1094),
   .I0(InputBits[134]),
   .I1(InputBits[204]),
   .I2(InputBits[298]),
   .I3(InputBits[146]),
   .I4(InputBits[526]),
   .I5(InputBits[68])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000110000000000000100010000000000110011)  
) LUT6_1095 (
   .O(gates_1095),
   .I0(InputBits[466]),
   .I1(InputBits[331]),
   .I2(InputBits[380]),
   .I3(InputBits[481]),
   .I4(InputBits[338]),
   .I5(InputBits[331])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000000001100000000000000110000000000010011)  
) LUT6_1096 (
   .O(gates_1096),
   .I0(InputBits[480]),
   .I1(InputBits[555]),
   .I2(InputBits[28]),
   .I3(InputBits[534]),
   .I4(InputBits[474]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0000000100000011000000000001010000000001000000110000000000000100)  
) LUT6_1097 (
   .O(gates_1097),
   .I0(InputBits[404]),
   .I1(InputBits[44]),
   .I2(InputBits[46]),
   .I3(InputBits[569]),
   .I4(InputBits[222]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0000000000010000000000110011101100000000000000000000001100010010)  
) LUT6_1098 (
   .O(gates_1098),
   .I0(InputBits[271]),
   .I1(InputBits[550]),
   .I2(InputBits[454]),
   .I3(InputBits[70]),
   .I4(InputBits[253]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0000000011011101000000000101110000000000010111010000010001011100)  
) LUT6_1099 (
   .O(gates_1099),
   .I0(InputBits[458]),
   .I1(InputBits[369]),
   .I2(InputBits[222]),
   .I3(InputBits[409]),
   .I4(InputBits[259]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0000000100010101011111111111111100000000000000001010111100001111)  
) LUT6_1100 (
   .O(gates_1100),
   .I0(InputBits[93]),
   .I1(InputBits[67]),
   .I2(InputBits[275]),
   .I3(InputBits[330]),
   .I4(InputBits[78]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0001000001010101000000000000000000000001010101010001010100010001)  
) LUT6_1101 (
   .O(gates_1101),
   .I0(InputBits[409]),
   .I1(InputBits[305]),
   .I2(InputBits[137]),
   .I3(InputBits[173]),
   .I4(InputBits[176]),
   .I5(InputBits[497])
);
LUT6 #(
   .INIT(64'b0000000000000000010000000001000000000000000000011111110111111111)  
) LUT6_1102 (
   .O(gates_1102),
   .I0(InputBits[86]),
   .I1(InputBits[466]),
   .I2(InputBits[413]),
   .I3(InputBits[137]),
   .I4(InputBits[551]),
   .I5(InputBits[100])
);
LUT6 #(
   .INIT(64'b0000001001000000010011000100000011111111011111111111111111110101)  
) LUT6_1103 (
   .O(gates_1103),
   .I0(InputBits[306]),
   .I1(InputBits[356]),
   .I2(InputBits[156]),
   .I3(InputBits[245]),
   .I4(InputBits[326]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0000010000000000000111110000101000001100000001000111111100101111)  
) LUT6_1104 (
   .O(gates_1104),
   .I0(InputBits[440]),
   .I1(InputBits[204]),
   .I2(InputBits[96]),
   .I3(InputBits[443]),
   .I4(InputBits[251]),
   .I5(InputBits[515])
);
LUT6 #(
   .INIT(64'b0011011100111111000101010000000100110111001011110001011100010011)  
) LUT6_1105 (
   .O(gates_1105),
   .I0(InputBits[255]),
   .I1(InputBits[228]),
   .I2(InputBits[101]),
   .I3(InputBits[446]),
   .I4(InputBits[419]),
   .I5(InputBits[513])
);
LUT6 #(
   .INIT(64'b0000111100001111000011110000111100001110000011110001111000001110)  
) LUT6_1106 (
   .O(gates_1106),
   .I0(InputBits[285]),
   .I1(InputBits[345]),
   .I2(InputBits[572]),
   .I3(InputBits[353]),
   .I4(InputBits[444]),
   .I5(InputBits[269])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000111100000000000001010000000000001110)  
) LUT6_1107 (
   .O(gates_1107),
   .I0(InputBits[93]),
   .I1(InputBits[190]),
   .I2(InputBits[576]),
   .I3(InputBits[576]),
   .I4(InputBits[525]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0000000000000000001101110001010001110000001100100111011100110111)  
) LUT6_1108 (
   .O(gates_1108),
   .I0(InputBits[68]),
   .I1(InputBits[548]),
   .I2(InputBits[225]),
   .I3(InputBits[247]),
   .I4(InputBits[250]),
   .I5(InputBits[495])
);
LUT6 #(
   .INIT(64'b0000101100100111000000010000010100001011000011110000000100000001)  
) LUT6_1109 (
   .O(gates_1109),
   .I0(InputBits[305]),
   .I1(InputBits[338]),
   .I2(InputBits[123]),
   .I3(InputBits[87]),
   .I4(InputBits[350]),
   .I5(InputBits[500])
);
LUT6 #(
   .INIT(64'b0000010000000100000000000000000011001100010011000001000000110010)  
) LUT6_1110 (
   .O(gates_1110),
   .I0(InputBits[92]),
   .I1(InputBits[421]),
   .I2(InputBits[524]),
   .I3(InputBits[422]),
   .I4(InputBits[421]),
   .I5(InputBits[36])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000001101000000000000000000001000100001110)  
) LUT6_1111 (
   .O(gates_1111),
   .I0(InputBits[13]),
   .I1(InputBits[12]),
   .I2(InputBits[222]),
   .I3(InputBits[188]),
   .I4(InputBits[573]),
   .I5(InputBits[210])
);
LUT6 #(
   .INIT(64'b0000000100001111000000000011111100000000000000110000000000000010)  
) LUT6_1112 (
   .O(gates_1112),
   .I0(InputBits[321]),
   .I1(InputBits[87]),
   .I2(InputBits[562]),
   .I3(InputBits[483]),
   .I4(InputBits[89]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b1000000000110000000000000011101000110110011100101111101011111111)  
) LUT6_1113 (
   .O(gates_1113),
   .I0(InputBits[222]),
   .I1(InputBits[546]),
   .I2(InputBits[202]),
   .I3(InputBits[129]),
   .I4(InputBits[487]),
   .I5(InputBits[251])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001000000000000001100110000000011111100)  
) LUT6_1114 (
   .O(gates_1114),
   .I0(InputBits[176]),
   .I1(InputBits[239]),
   .I2(InputBits[397]),
   .I3(InputBits[194]),
   .I4(InputBits[360]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0001010100010000000001010101000000000000000000000101010101010001)  
) LUT6_1115 (
   .O(gates_1115),
   .I0(InputBits[529]),
   .I1(InputBits[331]),
   .I2(InputBits[220]),
   .I3(InputBits[347]),
   .I4(InputBits[486]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000000000000111000111111101111100001010)  
) LUT6_1116 (
   .O(gates_1116),
   .I0(InputBits[335]),
   .I1(InputBits[303]),
   .I2(InputBits[37]),
   .I3(InputBits[418]),
   .I4(InputBits[245]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1101011101011101010100010101000011111101010101110010000000010101)  
) LUT6_1117 (
   .O(gates_1117),
   .I0(InputBits[53]),
   .I1(InputBits[255]),
   .I2(InputBits[424]),
   .I3(InputBits[57]),
   .I4(InputBits[393]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0010000011110010010000001111111110111010001110101111111111111111)  
) LUT6_1118 (
   .O(gates_1118),
   .I0(InputBits[325]),
   .I1(InputBits[111]),
   .I2(InputBits[223]),
   .I3(InputBits[476]),
   .I4(InputBits[277]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000000000000000011000000110000001000000010)  
) LUT6_1119 (
   .O(gates_1119),
   .I0(InputBits[65]),
   .I1(InputBits[482]),
   .I2(InputBits[565]),
   .I3(InputBits[322]),
   .I4(InputBits[115]),
   .I5(InputBits[232])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001111100000000000000000001000000010110)  
) LUT6_1120 (
   .O(gates_1120),
   .I0(InputBits[39]),
   .I1(InputBits[316]),
   .I2(InputBits[7]),
   .I3(InputBits[5]),
   .I4(InputBits[557]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100010000000100000011110110111111)  
) LUT6_1121 (
   .O(gates_1121),
   .I0(InputBits[513]),
   .I1(InputBits[549]),
   .I2(InputBits[226]),
   .I3(InputBits[515]),
   .I4(InputBits[564]),
   .I5(InputBits[266])
);
LUT6 #(
   .INIT(64'b0000000000000111000000000000000100000000000000110000000000000001)  
) LUT6_1122 (
   .O(gates_1122),
   .I0(InputBits[302]),
   .I1(InputBits[123]),
   .I2(InputBits[313]),
   .I3(InputBits[121]),
   .I4(InputBits[68]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000000000001000001000000011111101000000011101110010000000110101)  
) LUT6_1123 (
   .O(gates_1123),
   .I0(InputBits[451]),
   .I1(InputBits[280]),
   .I2(InputBits[465]),
   .I3(InputBits[55]),
   .I4(InputBits[239]),
   .I5(InputBits[220])
);
LUT6 #(
   .INIT(64'b0000000001010101000000000100000001111111111111010011110111111100)  
) LUT6_1124 (
   .O(gates_1124),
   .I0(InputBits[252]),
   .I1(InputBits[237]),
   .I2(InputBits[371]),
   .I3(InputBits[383]),
   .I4(InputBits[343]),
   .I5(InputBits[195])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000010100000000001101110100000100001111)  
) LUT6_1125 (
   .O(gates_1125),
   .I0(InputBits[78]),
   .I1(InputBits[522]),
   .I2(InputBits[509]),
   .I3(InputBits[252]),
   .I4(InputBits[428]),
   .I5(InputBits[253])
);
LUT6 #(
   .INIT(64'b1011001110111011000000111111101110000010111100000000001001010011)  
) LUT6_1126 (
   .O(gates_1126),
   .I0(InputBits[161]),
   .I1(InputBits[136]),
   .I2(InputBits[88]),
   .I3(InputBits[279]),
   .I4(InputBits[500]),
   .I5(InputBits[210])
);
LUT6 #(
   .INIT(64'b0000000001000101011100000101000100000000000001010111000001110001)  
) LUT6_1127 (
   .O(gates_1127),
   .I0(InputBits[149]),
   .I1(InputBits[280]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[45]),
   .I5(InputBits[185])
);
LUT6 #(
   .INIT(64'b0000000000000000000000111000001000010010001100110011001111111011)  
) LUT6_1128 (
   .O(gates_1128),
   .I0(InputBits[282]),
   .I1(InputBits[171]),
   .I2(InputBits[449]),
   .I3(InputBits[167]),
   .I4(InputBits[381]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0010000100110011001000000011001000110010001100100010000000110010)  
) LUT6_1129 (
   .O(gates_1129),
   .I0(InputBits[248]),
   .I1(InputBits[72]),
   .I2(InputBits[284]),
   .I3(InputBits[250]),
   .I4(InputBits[346]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b0000000000000011000000000000010000000000000010100000000001111111)  
) LUT6_1130 (
   .O(gates_1130),
   .I0(InputBits[40]),
   .I1(InputBits[301]),
   .I2(InputBits[150]),
   .I3(InputBits[538]),
   .I4(InputBits[299]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0000100100000011000011100000001100001101000000000100110100001101)  
) LUT6_1131 (
   .O(gates_1131),
   .I0(InputBits[489]),
   .I1(InputBits[245]),
   .I2(InputBits[75]),
   .I3(InputBits[198]),
   .I4(InputBits[81]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0101000101010100010101010100010001010001010101010100010001000100)  
) LUT6_1132 (
   .O(gates_1132),
   .I0(InputBits[51]),
   .I1(InputBits[268]),
   .I2(InputBits[180]),
   .I3(InputBits[296]),
   .I4(InputBits[393]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000100000000000000010101)  
) LUT6_1133 (
   .O(gates_1133),
   .I0(InputBits[102]),
   .I1(InputBits[88]),
   .I2(InputBits[71]),
   .I3(InputBits[529]),
   .I4(InputBits[470]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011000000000000001100010011001100110000)  
) LUT6_1134 (
   .O(gates_1134),
   .I0(InputBits[489]),
   .I1(InputBits[575]),
   .I2(InputBits[349]),
   .I3(InputBits[549]),
   .I4(InputBits[40]),
   .I5(InputBits[504])
);
LUT6 #(
   .INIT(64'b0101010101010101010011001100110001010101010100011111111011111111)  
) LUT6_1135 (
   .O(gates_1135),
   .I0(InputBits[191]),
   .I1(InputBits[246]),
   .I2(InputBits[157]),
   .I3(InputBits[404]),
   .I4(InputBits[407]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0000001000000111000000000000011100000010000000110000001000010011)  
) LUT6_1136 (
   .O(gates_1136),
   .I0(InputBits[245]),
   .I1(InputBits[483]),
   .I2(InputBits[572]),
   .I3(InputBits[230]),
   .I4(InputBits[203]),
   .I5(InputBits[438])
);
LUT6 #(
   .INIT(64'b0000000001110100000000000011000011101111111101110010111101110000)  
) LUT6_1137 (
   .O(gates_1137),
   .I0(InputBits[131]),
   .I1(InputBits[80]),
   .I2(InputBits[420]),
   .I3(InputBits[526]),
   .I4(InputBits[394]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0000000000000000000011110101111100010000000000000001010100010101)  
) LUT6_1138 (
   .O(gates_1138),
   .I0(InputBits[536]),
   .I1(InputBits[491]),
   .I2(InputBits[59]),
   .I3(InputBits[162]),
   .I4(InputBits[481]),
   .I5(InputBits[142])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000010100000101000000010000000100000101)  
) LUT6_1139 (
   .O(gates_1139),
   .I0(InputBits[575]),
   .I1(InputBits[474]),
   .I2(InputBits[124]),
   .I3(InputBits[545]),
   .I4(InputBits[306]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0000000000000101110111011101111100000000000001011101110101001101)  
) LUT6_1140 (
   .O(gates_1140),
   .I0(InputBits[494]),
   .I1(InputBits[416]),
   .I2(InputBits[127]),
   .I3(InputBits[477]),
   .I4(InputBits[14]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000000000100000000000000010001000010011001111110000000000101111)  
) LUT6_1141 (
   .O(gates_1141),
   .I0(InputBits[234]),
   .I1(InputBits[232]),
   .I2(InputBits[131]),
   .I3(InputBits[508]),
   .I4(InputBits[180]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0000000100000001000100010001000100010000000101010001000100010001)  
) LUT6_1142 (
   .O(gates_1142),
   .I0(InputBits[27]),
   .I1(InputBits[459]),
   .I2(InputBits[239]),
   .I3(InputBits[110]),
   .I4(InputBits[536]),
   .I5(InputBits[143])
);
LUT6 #(
   .INIT(64'b0001000000000000110001001000000001010000111011001111111111111101)  
) LUT6_1143 (
   .O(gates_1143),
   .I0(InputBits[523]),
   .I1(InputBits[414]),
   .I2(InputBits[161]),
   .I3(InputBits[221]),
   .I4(InputBits[459]),
   .I5(InputBits[493])
);
LUT6 #(
   .INIT(64'b0011001000110010001100100011001000100010001000100011001000111010)  
) LUT6_1144 (
   .O(gates_1144),
   .I0(InputBits[293]),
   .I1(InputBits[574]),
   .I2(InputBits[374]),
   .I3(InputBits[435]),
   .I4(InputBits[486]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101000001110000000101000101)  
) LUT6_1145 (
   .O(gates_1145),
   .I0(InputBits[434]),
   .I1(InputBits[178]),
   .I2(InputBits[536]),
   .I3(InputBits[568]),
   .I4(InputBits[321]),
   .I5(InputBits[145])
);
LUT6 #(
   .INIT(64'b0000000000000001001100010011001100000001000000010011000101110001)  
) LUT6_1146 (
   .O(gates_1146),
   .I0(InputBits[107]),
   .I1(InputBits[508]),
   .I2(InputBits[334]),
   .I3(InputBits[108]),
   .I4(InputBits[6]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0000000000010000000011100000011100000000000000100000101000001111)  
) LUT6_1147 (
   .O(gates_1147),
   .I0(InputBits[198]),
   .I1(InputBits[155]),
   .I2(InputBits[170]),
   .I3(InputBits[471]),
   .I4(InputBits[171]),
   .I5(InputBits[66])
);
LUT6 #(
   .INIT(64'b0000001100000011000000110000001100000011000000110000001100000010)  
) LUT6_1148 (
   .O(gates_1148),
   .I0(InputBits[367]),
   .I1(InputBits[529]),
   .I2(InputBits[73]),
   .I3(InputBits[442]),
   .I4(InputBits[202]),
   .I5(InputBits[335])
);
LUT6 #(
   .INIT(64'b0000000000000000111110110001001000000000000000000111111000000010)  
) LUT6_1149 (
   .O(gates_1149),
   .I0(InputBits[315]),
   .I1(InputBits[387]),
   .I2(InputBits[415]),
   .I3(InputBits[178]),
   .I4(InputBits[573]),
   .I5(InputBits[211])
);
LUT6 #(
   .INIT(64'b0000111100001111000011110001111100001111000000010000111100000101)  
) LUT6_1150 (
   .O(gates_1150),
   .I0(InputBits[495]),
   .I1(InputBits[132]),
   .I2(InputBits[170]),
   .I3(InputBits[286]),
   .I4(InputBits[208]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0000000000000101000100000000110000000100000111010001010100001101)  
) LUT6_1151 (
   .O(gates_1151),
   .I0(InputBits[508]),
   .I1(InputBits[428]),
   .I2(InputBits[473]),
   .I3(InputBits[549]),
   .I4(InputBits[406]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b0000000000000010000000000000001100000000000100000000000000010011)  
) LUT6_1152 (
   .O(gates_1152),
   .I0(InputBits[9]),
   .I1(InputBits[481]),
   .I2(InputBits[363]),
   .I3(InputBits[72]),
   .I4(InputBits[205]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b0000000000000010000010001000101000000000000000110000101000011011)  
) LUT6_1153 (
   .O(gates_1153),
   .I0(InputBits[368]),
   .I1(InputBits[254]),
   .I2(InputBits[562]),
   .I3(InputBits[482]),
   .I4(InputBits[543]),
   .I5(InputBits[206])
);
LUT6 #(
   .INIT(64'b0000000000000000000001000000000000000000000000000100010000000001)  
) LUT6_1154 (
   .O(gates_1154),
   .I0(InputBits[289]),
   .I1(InputBits[221]),
   .I2(InputBits[512]),
   .I3(InputBits[221]),
   .I4(InputBits[27]),
   .I5(InputBits[507])
);
LUT6 #(
   .INIT(64'b0000000100110011001100110011001100000000000100110001000000000001)  
) LUT6_1155 (
   .O(gates_1155),
   .I0(InputBits[452]),
   .I1(InputBits[552]),
   .I2(InputBits[112]),
   .I3(InputBits[10]),
   .I4(InputBits[383]),
   .I5(InputBits[415])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000010111000001010001010101010100)  
) LUT6_1156 (
   .O(gates_1156),
   .I0(InputBits[532]),
   .I1(InputBits[287]),
   .I2(InputBits[478]),
   .I3(InputBits[365]),
   .I4(InputBits[202]),
   .I5(InputBits[218])
);
LUT6 #(
   .INIT(64'b0000000000000000010000000000010100000000000000000001000000000111)  
) LUT6_1157 (
   .O(gates_1157),
   .I0(InputBits[134]),
   .I1(InputBits[329]),
   .I2(InputBits[208]),
   .I3(InputBits[208]),
   .I4(InputBits[555]),
   .I5(InputBits[520])
);
LUT6 #(
   .INIT(64'b0000111100001100000011110000110000000100000011000000110000001100)  
) LUT6_1158 (
   .O(gates_1158),
   .I0(InputBits[452]),
   .I1(InputBits[237]),
   .I2(InputBits[566]),
   .I3(InputBits[315]),
   .I4(InputBits[356]),
   .I5(InputBits[198])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000111000100011001011111010)  
) LUT6_1159 (
   .O(gates_1159),
   .I0(InputBits[200]),
   .I1(InputBits[111]),
   .I2(InputBits[350]),
   .I3(InputBits[168]),
   .I4(InputBits[569]),
   .I5(InputBits[505])
);
LUT6 #(
   .INIT(64'b1111111111111111000100001111101011101110011111111111001011111010)  
) LUT6_1160 (
   .O(gates_1160),
   .I0(InputBits[139]),
   .I1(InputBits[327]),
   .I2(InputBits[444]),
   .I3(InputBits[87]),
   .I4(InputBits[364]),
   .I5(InputBits[162])
);
LUT6 #(
   .INIT(64'b0000000000010000000000000000000000000000000100110101000101000110)  
) LUT6_1161 (
   .O(gates_1161),
   .I0(InputBits[96]),
   .I1(InputBits[7]),
   .I2(InputBits[428]),
   .I3(InputBits[10]),
   .I4(InputBits[222]),
   .I5(InputBits[170])
);
LUT6 #(
   .INIT(64'b0000100000010001000001100000001010101010101111111011101000111011)  
) LUT6_1162 (
   .O(gates_1162),
   .I0(InputBits[391]),
   .I1(InputBits[125]),
   .I2(InputBits[388]),
   .I3(InputBits[105]),
   .I4(InputBits[258]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1101010111010001001100010001010110110011101110110010001010100000)  
) LUT6_1163 (
   .O(gates_1163),
   .I0(InputBits[215]),
   .I1(InputBits[250]),
   .I2(InputBits[135]),
   .I3(InputBits[153]),
   .I4(InputBits[248]),
   .I5(InputBits[393])
);
LUT6 #(
   .INIT(64'b0000001000000011000000100100111100000010000000000000000001000000)  
) LUT6_1164 (
   .O(gates_1164),
   .I0(InputBits[204]),
   .I1(InputBits[327]),
   .I2(InputBits[570]),
   .I3(InputBits[133]),
   .I4(InputBits[88]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001001111100000000000000000000110010001100)  
) LUT6_1165 (
   .O(gates_1165),
   .I0(InputBits[467]),
   .I1(InputBits[248]),
   .I2(InputBits[459]),
   .I3(InputBits[565]),
   .I4(InputBits[230]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b0000010100000011000001110001001101001101010001110000010000000000)  
) LUT6_1166 (
   .O(gates_1166),
   .I0(InputBits[488]),
   .I1(InputBits[305]),
   .I2(InputBits[266]),
   .I3(InputBits[399]),
   .I4(InputBits[348]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000001011000000110000101100000010)  
) LUT6_1167 (
   .O(gates_1167),
   .I0(InputBits[317]),
   .I1(InputBits[255]),
   .I2(InputBits[99]),
   .I3(InputBits[200]),
   .I4(InputBits[391]),
   .I5(InputBits[507])
);
LUT6 #(
   .INIT(64'b0000000001000100000011000000110000000101000001000100111000001110)  
) LUT6_1168 (
   .O(gates_1168),
   .I0(InputBits[15]),
   .I1(InputBits[366]),
   .I2(InputBits[54]),
   .I3(InputBits[139]),
   .I4(InputBits[157]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b0010101100000011000011110000001100001111000001010000111100000101)  
) LUT6_1169 (
   .O(gates_1169),
   .I0(InputBits[495]),
   .I1(InputBits[151]),
   .I2(InputBits[361]),
   .I3(InputBits[294]),
   .I4(InputBits[90]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000011001100000000000000000000000011001101)  
) LUT6_1170 (
   .O(gates_1170),
   .I0(InputBits[424]),
   .I1(InputBits[94]),
   .I2(InputBits[435]),
   .I3(InputBits[2]),
   .I4(InputBits[555]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0101010101010001010001010100000100000101000001000000000000000110)  
) LUT6_1171 (
   .O(gates_1171),
   .I0(InputBits[96]),
   .I1(InputBits[67]),
   .I2(InputBits[435]),
   .I3(InputBits[66]),
   .I4(InputBits[113]),
   .I5(InputBits[213])
);
LUT6 #(
   .INIT(64'b0000001000010111000000000001011100000000000001110000000000000001)  
) LUT6_1172 (
   .O(gates_1172),
   .I0(InputBits[461]),
   .I1(InputBits[434]),
   .I2(InputBits[75]),
   .I3(InputBits[511]),
   .I4(InputBits[163]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b0000000000001011000000010000000000001100000011110000010011111111)  
) LUT6_1173 (
   .O(gates_1173),
   .I0(InputBits[357]),
   .I1(InputBits[452]),
   .I2(InputBits[12]),
   .I3(InputBits[266]),
   .I4(InputBits[188]),
   .I5(InputBits[495])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000110000000111110001)  
) LUT6_1174 (
   .O(gates_1174),
   .I0(InputBits[110]),
   .I1(InputBits[499]),
   .I2(InputBits[214]),
   .I3(InputBits[46]),
   .I4(InputBits[9]),
   .I5(InputBits[558])
);
LUT6 #(
   .INIT(64'b0000000000000000000000110000001100000010000000110011001100111000)  
) LUT6_1175 (
   .O(gates_1175),
   .I0(InputBits[164]),
   .I1(InputBits[565]),
   .I2(InputBits[359]),
   .I3(InputBits[416]),
   .I4(InputBits[143]),
   .I5(InputBits[243])
);
LUT6 #(
   .INIT(64'b0000000101011111000100000111111100000000010101010000000011011100)  
) LUT6_1176 (
   .O(gates_1176),
   .I0(InputBits[493]),
   .I1(InputBits[198]),
   .I2(InputBits[441]),
   .I3(InputBits[482]),
   .I4(InputBits[324]),
   .I5(InputBits[93])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000000000000100000101)  
) LUT6_1177 (
   .O(gates_1177),
   .I0(InputBits[128]),
   .I1(InputBits[6]),
   .I2(InputBits[409]),
   .I3(InputBits[296]),
   .I4(InputBits[461]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0011001100010011001100110000001100010011000000000011101100010011)  
) LUT6_1178 (
   .O(gates_1178),
   .I0(InputBits[280]),
   .I1(InputBits[242]),
   .I2(InputBits[469]),
   .I3(InputBits[344]),
   .I4(InputBits[82]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0000000000000000001110110011001000000000000000000011001100010000)  
) LUT6_1179 (
   .O(gates_1179),
   .I0(InputBits[281]),
   .I1(InputBits[559]),
   .I2(InputBits[445]),
   .I3(InputBits[311]),
   .I4(InputBits[51]),
   .I5(InputBits[323])
);
LUT6 #(
   .INIT(64'b0000000000000000000000101111110000000000000000000000100011110001)  
) LUT6_1180 (
   .O(gates_1180),
   .I0(InputBits[425]),
   .I1(InputBits[58]),
   .I2(InputBits[335]),
   .I3(InputBits[314]),
   .I4(InputBits[25]),
   .I5(InputBits[151])
);
LUT6 #(
   .INIT(64'b0000111100101111000001000001111100010111110011010001011101111111)  
) LUT6_1181 (
   .O(gates_1181),
   .I0(InputBits[520]),
   .I1(InputBits[524]),
   .I2(InputBits[205]),
   .I3(InputBits[243]),
   .I4(InputBits[450]),
   .I5(InputBits[547])
);
LUT6 #(
   .INIT(64'b0100010001010000000000000111000001010101010111010001000101010101)  
) LUT6_1182 (
   .O(gates_1182),
   .I0(InputBits[536]),
   .I1(InputBits[112]),
   .I2(InputBits[326]),
   .I3(InputBits[486]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000111010101000000001110110000000001110111110100010111101111)  
) LUT6_1183 (
   .O(gates_1183),
   .I0(InputBits[358]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[216]),
   .I4(InputBits[118]),
   .I5(InputBits[473])
);
LUT6 #(
   .INIT(64'b0000000000111101000000000111110100000000001111000000000010111110)  
) LUT6_1184 (
   .O(gates_1184),
   .I0(InputBits[296]),
   .I1(InputBits[384]),
   .I2(InputBits[212]),
   .I3(InputBits[24]),
   .I4(InputBits[463]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b0000000000000001000011111011001100000011000011110000111111010001)  
) LUT6_1185 (
   .O(gates_1185),
   .I0(InputBits[207]),
   .I1(InputBits[232]),
   .I2(InputBits[360]),
   .I3(InputBits[431]),
   .I4(InputBits[13]),
   .I5(InputBits[157])
);
LUT6 #(
   .INIT(64'b0000000000000000000000001000001000000000111000000000000111101111)  
) LUT6_1186 (
   .O(gates_1186),
   .I0(InputBits[187]),
   .I1(InputBits[156]),
   .I2(InputBits[203]),
   .I3(InputBits[9]),
   .I4(InputBits[484]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010000000000110001001100000011001100000000)  
) LUT6_1187 (
   .O(gates_1187),
   .I0(InputBits[196]),
   .I1(InputBits[529]),
   .I2(InputBits[165]),
   .I3(InputBits[420]),
   .I4(InputBits[180]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1110110011111110001011100101111000001100110010001110111111001100)  
) LUT6_1188 (
   .O(gates_1188),
   .I0(InputBits[334]),
   .I1(InputBits[269]),
   .I2(InputBits[64]),
   .I3(InputBits[209]),
   .I4(InputBits[112]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0000110000000100000000000000010000000101000001010000110000000101)  
) LUT6_1189 (
   .O(gates_1189),
   .I0(InputBits[508]),
   .I1(InputBits[69]),
   .I2(InputBits[3]),
   .I3(InputBits[462]),
   .I4(InputBits[153]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010011001100000000000000000001010110100010)  
) LUT6_1190 (
   .O(gates_1190),
   .I0(InputBits[176]),
   .I1(InputBits[132]),
   .I2(InputBits[139]),
   .I3(InputBits[15]),
   .I4(InputBits[409]),
   .I5(InputBits[323])
);
LUT6 #(
   .INIT(64'b0111001111110111001000011111111110110111110111010001011101010101)  
) LUT6_1191 (
   .O(gates_1191),
   .I0(InputBits[492]),
   .I1(InputBits[429]),
   .I2(InputBits[467]),
   .I3(InputBits[118]),
   .I4(InputBits[165]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000010000000011011111)  
) LUT6_1192 (
   .O(gates_1192),
   .I0(InputBits[253]),
   .I1(InputBits[360]),
   .I2(InputBits[130]),
   .I3(InputBits[1]),
   .I4(InputBits[559]),
   .I5(InputBits[265])
);
LUT6 #(
   .INIT(64'b0001000111010000000111111111010000001111010111000001111101010111)  
) LUT6_1193 (
   .O(gates_1193),
   .I0(InputBits[490]),
   .I1(InputBits[162]),
   .I2(InputBits[58]),
   .I3(InputBits[118]),
   .I4(InputBits[473]),
   .I5(InputBits[150])
);
LUT6 #(
   .INIT(64'b0001000101010001010100000101010100010101010101010100010001000101)  
) LUT6_1194 (
   .O(gates_1194),
   .I0(InputBits[530]),
   .I1(InputBits[37]),
   .I2(InputBits[425]),
   .I3(InputBits[150]),
   .I4(InputBits[246]),
   .I5(InputBits[364])
);
LUT6 #(
   .INIT(64'b0101000011011011010100000101000001111101011111010101110011110100)  
) LUT6_1195 (
   .O(gates_1195),
   .I0(InputBits[196]),
   .I1(InputBits[283]),
   .I2(InputBits[286]),
   .I3(InputBits[140]),
   .I4(InputBits[340]),
   .I5(InputBits[207])
);
LUT6 #(
   .INIT(64'b0011000000110111000000000000000000110001001101110011010100000001)  
) LUT6_1196 (
   .O(gates_1196),
   .I0(InputBits[511]),
   .I1(InputBits[148]),
   .I2(InputBits[227]),
   .I3(InputBits[143]),
   .I4(InputBits[366]),
   .I5(InputBits[436])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000101000000110000000100001010)  
) LUT6_1197 (
   .O(gates_1197),
   .I0(InputBits[502]),
   .I1(InputBits[483]),
   .I2(InputBits[27]),
   .I3(InputBits[68]),
   .I4(InputBits[189]),
   .I5(InputBits[530])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100010000000000000100110100000010011111111)  
) LUT6_1198 (
   .O(gates_1198),
   .I0(InputBits[424]),
   .I1(InputBits[130]),
   .I2(InputBits[524]),
   .I3(InputBits[338]),
   .I4(InputBits[77]),
   .I5(InputBits[251])
);
LUT6 #(
   .INIT(64'b0000000000000000000000100001001100000000000000000000000000100010)  
) LUT6_1199 (
   .O(gates_1199),
   .I0(InputBits[268]),
   .I1(InputBits[193]),
   .I2(InputBits[484]),
   .I3(InputBits[255]),
   .I4(InputBits[145]),
   .I5(InputBits[367])
);
LUT6 #(
   .INIT(64'b0000000000010010000000000010000000000000000100100000000000010000)  
) LUT6_1200 (
   .O(gates_1200),
   .I0(InputBits[41]),
   .I1(InputBits[50]),
   .I2(InputBits[213]),
   .I3(InputBits[52]),
   .I4(InputBits[499]),
   .I5(InputBits[305])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000001000000010000010000000111)  
) LUT6_1201 (
   .O(gates_1201),
   .I0(InputBits[551]),
   .I1(InputBits[407]),
   .I2(InputBits[123]),
   .I3(InputBits[279]),
   .I4(InputBits[166]),
   .I5(InputBits[566])
);
LUT6 #(
   .INIT(64'b0000000000001111010000001111001000000000001100111110001111111111)  
) LUT6_1202 (
   .O(gates_1202),
   .I0(InputBits[351]),
   .I1(InputBits[469]),
   .I2(InputBits[332]),
   .I3(InputBits[513]),
   .I4(InputBits[12]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010001000000010000001110000001000000011)  
) LUT6_1203 (
   .O(gates_1203),
   .I0(InputBits[309]),
   .I1(InputBits[28]),
   .I2(InputBits[194]),
   .I3(InputBits[471]),
   .I4(InputBits[86]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0011001100110011001100110011011100110011000000010011101110011101)  
) LUT6_1204 (
   .O(gates_1204),
   .I0(InputBits[106]),
   .I1(InputBits[550]),
   .I2(InputBits[155]),
   .I3(InputBits[358]),
   .I4(InputBits[164]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0000000000000000100000001111111100000000010101011000110111001100)  
) LUT6_1205 (
   .O(gates_1205),
   .I0(InputBits[140]),
   .I1(InputBits[395]),
   .I2(InputBits[207]),
   .I3(InputBits[120]),
   .I4(InputBits[408]),
   .I5(InputBits[261])
);
LUT6 #(
   .INIT(64'b0000000010001000000000001101100000000000101100110000000011111011)  
) LUT6_1206 (
   .O(gates_1206),
   .I0(InputBits[90]),
   .I1(InputBits[451]),
   .I2(InputBits[163]),
   .I3(InputBits[560]),
   .I4(InputBits[323]),
   .I5(InputBits[447])
);
LUT6 #(
   .INIT(64'b0000000000000000000100000000000000000000000000000001000100010001)  
) LUT6_1207 (
   .O(gates_1207),
   .I0(InputBits[82]),
   .I1(InputBits[409]),
   .I2(InputBits[331]),
   .I3(InputBits[403]),
   .I4(InputBits[361]),
   .I5(InputBits[266])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000000010000000000000001111)  
) LUT6_1208 (
   .O(gates_1208),
   .I0(InputBits[450]),
   .I1(InputBits[405]),
   .I2(InputBits[313]),
   .I3(InputBits[27]),
   .I4(InputBits[539]),
   .I5(InputBits[255])
);
LUT6 #(
   .INIT(64'b0000000000000101000000010000010100000000000001000000000001000111)  
) LUT6_1209 (
   .O(gates_1209),
   .I0(InputBits[17]),
   .I1(InputBits[68]),
   .I2(InputBits[277]),
   .I3(InputBits[7]),
   .I4(InputBits[158]),
   .I5(InputBits[135])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010000001100000011000010110000)  
) LUT6_1210 (
   .O(gates_1210),
   .I0(InputBits[181]),
   .I1(InputBits[561]),
   .I2(InputBits[372]),
   .I3(InputBits[487]),
   .I4(InputBits[120]),
   .I5(InputBits[563])
);
LUT6 #(
   .INIT(64'b0000010100000101000000010111011100000001000001010000000000010001)  
) LUT6_1211 (
   .O(gates_1211),
   .I0(InputBits[410]),
   .I1(InputBits[537]),
   .I2(InputBits[543]),
   .I3(InputBits[230]),
   .I4(InputBits[239]),
   .I5(InputBits[341])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000011001011110000111100101010)  
) LUT6_1212 (
   .O(gates_1212),
   .I0(InputBits[347]),
   .I1(InputBits[297]),
   .I2(InputBits[53]),
   .I3(InputBits[267]),
   .I4(InputBits[388]),
   .I5(InputBits[1])
);
LUT6 #(
   .INIT(64'b0110110001111100000100000101110000000100000111010001000011111111)  
) LUT6_1213 (
   .O(gates_1213),
   .I0(InputBits[305]),
   .I1(InputBits[369]),
   .I2(InputBits[262]),
   .I3(InputBits[533]),
   .I4(InputBits[229]),
   .I5(InputBits[251])
);
LUT6 #(
   .INIT(64'b0000000000000101000000000000010101000100000011000110011101001101)  
) LUT6_1214 (
   .O(gates_1214),
   .I0(InputBits[53]),
   .I1(InputBits[421]),
   .I2(InputBits[516]),
   .I3(InputBits[197]),
   .I4(InputBits[436]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001100000000000001000000000000001100)  
) LUT6_1215 (
   .O(gates_1215),
   .I0(InputBits[89]),
   .I1(InputBits[549]),
   .I2(InputBits[482]),
   .I3(InputBits[53]),
   .I4(InputBits[273]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b0010001100110000001111110001100000110011000100100111011100010100)  
) LUT6_1216 (
   .O(gates_1216),
   .I0(InputBits[428]),
   .I1(InputBits[480]),
   .I2(InputBits[381]),
   .I3(InputBits[394]),
   .I4(InputBits[91]),
   .I5(InputBits[427])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000010000000000110111000000000001000100)  
) LUT6_1217 (
   .O(gates_1217),
   .I0(InputBits[562]),
   .I1(InputBits[349]),
   .I2(InputBits[227]),
   .I3(InputBits[265]),
   .I4(InputBits[141]),
   .I5(InputBits[196])
);
LUT6 #(
   .INIT(64'b0000111100001111011111110000001100001011000011110000011100000011)  
) LUT6_1218 (
   .O(gates_1218),
   .I0(InputBits[163]),
   .I1(InputBits[133]),
   .I2(InputBits[557]),
   .I3(InputBits[211]),
   .I4(InputBits[501]),
   .I5(InputBits[466])
);
LUT6 #(
   .INIT(64'b0011001100010010001000110000001100100010001000100000001000000010)  
) LUT6_1219 (
   .O(gates_1219),
   .I0(InputBits[263]),
   .I1(InputBits[505]),
   .I2(InputBits[498]),
   .I3(InputBits[152]),
   .I4(InputBits[438]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000001100000000000000000000000000000011)  
) LUT6_1220 (
   .O(gates_1220),
   .I0(InputBits[525]),
   .I1(InputBits[72]),
   .I2(InputBits[533]),
   .I3(InputBits[560]),
   .I4(InputBits[4]),
   .I5(InputBits[173])
);
LUT6 #(
   .INIT(64'b0000000000000000010011101110100000000001000000000111111111111111)  
) LUT6_1221 (
   .O(gates_1221),
   .I0(InputBits[465]),
   .I1(InputBits[199]),
   .I2(InputBits[431]),
   .I3(InputBits[320]),
   .I4(InputBits[51]),
   .I5(InputBits[495])
);
LUT6 #(
   .INIT(64'b0000000000000010010101010101010100000000010001101111010111110111)  
) LUT6_1222 (
   .O(gates_1222),
   .I0(InputBits[277]),
   .I1(InputBits[462]),
   .I2(InputBits[405]),
   .I3(InputBits[108]),
   .I4(InputBits[229]),
   .I5(InputBits[517])
);
LUT6 #(
   .INIT(64'b0000000011101111000000011110111100000000101111110000000110101110)  
) LUT6_1223 (
   .O(gates_1223),
   .I0(InputBits[393]),
   .I1(InputBits[413]),
   .I2(InputBits[488]),
   .I3(InputBits[571]),
   .I4(InputBits[347]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000010011111100110011010101010101)  
) LUT6_1224 (
   .O(gates_1224),
   .I0(InputBits[518]),
   .I1(InputBits[384]),
   .I2(InputBits[162]),
   .I3(InputBits[90]),
   .I4(InputBits[163]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b1100001101001100001111110100010011110111111111111111110111110101)  
) LUT6_1225 (
   .O(gates_1225),
   .I0(InputBits[488]),
   .I1(InputBits[244]),
   .I2(InputBits[357]),
   .I3(InputBits[422]),
   .I4(InputBits[308]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0000000000000000111111111001111000000001000000011111111100111111)  
) LUT6_1226 (
   .O(gates_1226),
   .I0(InputBits[407]),
   .I1(InputBits[282]),
   .I2(InputBits[332]),
   .I3(InputBits[366]),
   .I4(InputBits[504]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0000000000010001000100010001001100000000000100000000000000010000)  
) LUT6_1227 (
   .O(gates_1227),
   .I0(InputBits[482]),
   .I1(InputBits[1]),
   .I2(InputBits[430]),
   .I3(InputBits[306]),
   .I4(InputBits[465]),
   .I5(InputBits[388])
);
LUT6 #(
   .INIT(64'b0000001100000011000000110000101100010111000000110000110100000011)  
) LUT6_1228 (
   .O(gates_1228),
   .I0(InputBits[330]),
   .I1(InputBits[527]),
   .I2(InputBits[481]),
   .I3(InputBits[255]),
   .I4(InputBits[346]),
   .I5(InputBits[317])
);
LUT6 #(
   .INIT(64'b0000111000001110001010100101111110001110000001100000110001001111)  
) LUT6_1229 (
   .O(gates_1229),
   .I0(InputBits[523]),
   .I1(InputBits[325]),
   .I2(InputBits[518]),
   .I3(InputBits[108]),
   .I4(InputBits[56]),
   .I5(InputBits[424])
);
LUT6 #(
   .INIT(64'b0000000011001101000000000100010000000000110011000000000011001101)  
) LUT6_1230 (
   .O(gates_1230),
   .I0(InputBits[110]),
   .I1(InputBits[318]),
   .I2(InputBits[427]),
   .I3(InputBits[289]),
   .I4(InputBits[413]),
   .I5(InputBits[173])
);
LUT6 #(
   .INIT(64'b0011001100000000001100100001000000110011000100110011000100110000)  
) LUT6_1231 (
   .O(gates_1231),
   .I0(InputBits[389]),
   .I1(InputBits[561]),
   .I2(InputBits[407]),
   .I3(InputBits[366]),
   .I4(InputBits[319]),
   .I5(InputBits[450])
);
LUT6 #(
   .INIT(64'b0010111100001111001011110010011100100011000111110011011100111100)  
) LUT6_1232 (
   .O(gates_1232),
   .I0(InputBits[358]),
   .I1(InputBits[291]),
   .I2(InputBits[360]),
   .I3(InputBits[397]),
   .I4(InputBits[365]),
   .I5(InputBits[201])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000000000000001000000110001000000011111)  
) LUT6_1233 (
   .O(gates_1233),
   .I0(InputBits[43]),
   .I1(InputBits[16]),
   .I2(InputBits[570]),
   .I3(InputBits[148]),
   .I4(InputBits[286]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000001010100010101000101010001010001011111)  
) LUT6_1234 (
   .O(gates_1234),
   .I0(InputBits[495]),
   .I1(InputBits[475]),
   .I2(InputBits[229]),
   .I3(InputBits[100]),
   .I4(InputBits[77]),
   .I5(InputBits[45])
);
LUT6 #(
   .INIT(64'b0000000000000000000011110100101100000010000000000001110001011010)  
) LUT6_1235 (
   .O(gates_1235),
   .I0(InputBits[270]),
   .I1(InputBits[389]),
   .I2(InputBits[14]),
   .I3(InputBits[157]),
   .I4(InputBits[557]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0001000011111111110100001111111101000100010001000110010011101110)  
) LUT6_1236 (
   .O(gates_1236),
   .I0(InputBits[340]),
   .I1(InputBits[396]),
   .I2(InputBits[401]),
   .I3(InputBits[100]),
   .I4(InputBits[86]),
   .I5(InputBits[342])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000010111110000000000010101)  
) LUT6_1237 (
   .O(gates_1237),
   .I0(InputBits[194]),
   .I1(InputBits[110]),
   .I2(InputBits[298]),
   .I3(InputBits[289]),
   .I4(InputBits[370]),
   .I5(InputBits[193])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000100110011101110)  
) LUT6_1238 (
   .O(gates_1238),
   .I0(InputBits[191]),
   .I1(InputBits[318]),
   .I2(InputBits[187]),
   .I3(InputBits[65]),
   .I4(InputBits[507]),
   .I5(InputBits[552])
);
LUT6 #(
   .INIT(64'b0000001100000010000001010000011100000010010101100000001100000011)  
) LUT6_1239 (
   .O(gates_1239),
   .I0(InputBits[34]),
   .I1(InputBits[521]),
   .I2(InputBits[242]),
   .I3(InputBits[158]),
   .I4(InputBits[377]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000010000000000000000010000010100010101)  
) LUT6_1240 (
   .O(gates_1240),
   .I0(InputBits[72]),
   .I1(InputBits[339]),
   .I2(InputBits[264]),
   .I3(InputBits[438]),
   .I4(InputBits[551]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0000000100000010000000000000001000000000001000100000000000100010)  
) LUT6_1241 (
   .O(gates_1241),
   .I0(InputBits[367]),
   .I1(InputBits[386]),
   .I2(InputBits[195]),
   .I3(InputBits[314]),
   .I4(InputBits[249]),
   .I5(InputBits[164])
);
LUT6 #(
   .INIT(64'b0000000100110000000000110011000100000000001101010000000100110101)  
) LUT6_1242 (
   .O(gates_1242),
   .I0(InputBits[79]),
   .I1(InputBits[144]),
   .I2(InputBits[525]),
   .I3(InputBits[53]),
   .I4(InputBits[281]),
   .I5(InputBits[86])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000010000100110010001110100000000011111010)  
) LUT6_1243 (
   .O(gates_1243),
   .I0(InputBits[345]),
   .I1(InputBits[471]),
   .I2(InputBits[324]),
   .I3(InputBits[562]),
   .I4(InputBits[492]),
   .I5(InputBits[45])
);
LUT6 #(
   .INIT(64'b0000000000000111000000000000000000000000000001110000000100000100)  
) LUT6_1244 (
   .O(gates_1244),
   .I0(InputBits[172]),
   .I1(InputBits[272]),
   .I2(InputBits[97]),
   .I3(InputBits[528]),
   .I4(InputBits[190]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0000000011111111001000101110101000000000111011100000000110101110)  
) LUT6_1245 (
   .O(gates_1245),
   .I0(InputBits[236]),
   .I1(InputBits[199]),
   .I2(InputBits[113]),
   .I3(InputBits[43]),
   .I4(InputBits[333]),
   .I5(InputBits[66])
);
LUT6 #(
   .INIT(64'b0000000000110110000000000111111100000000000000100000000010111010)  
) LUT6_1246 (
   .O(gates_1246),
   .I0(InputBits[247]),
   .I1(InputBits[499]),
   .I2(InputBits[118]),
   .I3(InputBits[409]),
   .I4(InputBits[459]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b0011000001110010001000110101000100100010011100110001001100010000)  
) LUT6_1247 (
   .O(gates_1247),
   .I0(InputBits[175]),
   .I1(InputBits[561]),
   .I2(InputBits[202]),
   .I3(InputBits[454]),
   .I4(InputBits[270]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0001110100001100000001010100111111101100110011000000110011111110)  
) LUT6_1248 (
   .O(gates_1248),
   .I0(InputBits[382]),
   .I1(InputBits[372]),
   .I2(InputBits[38]),
   .I3(InputBits[330]),
   .I4(InputBits[329]),
   .I5(InputBits[117])
);
LUT6 #(
   .INIT(64'b0000000000010000101000100001100100110010000100001111111110011101)  
) LUT6_1249 (
   .O(gates_1249),
   .I0(InputBits[135]),
   .I1(InputBits[183]),
   .I2(InputBits[258]),
   .I3(InputBits[202]),
   .I4(InputBits[128]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0000010100110011000011010011111100000000000000100000100000111111)  
) LUT6_1250 (
   .O(gates_1250),
   .I0(InputBits[356]),
   .I1(InputBits[131]),
   .I2(InputBits[299]),
   .I3(InputBits[81]),
   .I4(InputBits[125]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0001000100110000001100110011000100100000000000000011001100110110)  
) LUT6_1251 (
   .O(gates_1251),
   .I0(InputBits[296]),
   .I1(InputBits[18]),
   .I2(InputBits[349]),
   .I3(InputBits[175]),
   .I4(InputBits[126]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b0000111100001111000011110000111100001111000111100000111100001111)  
) LUT6_1252 (
   .O(gates_1252),
   .I0(InputBits[443]),
   .I1(InputBits[388]),
   .I2(InputBits[361]),
   .I3(InputBits[430]),
   .I4(InputBits[134]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000000000000100000000000000000000000100010101000000000001010100)  
) LUT6_1253 (
   .O(gates_1253),
   .I0(InputBits[553]),
   .I1(InputBits[373]),
   .I2(InputBits[334]),
   .I3(InputBits[75]),
   .I4(InputBits[233]),
   .I5(InputBits[242])
);
LUT6 #(
   .INIT(64'b0000000100000101000010100000111100000101000001010000001100001111)  
) LUT6_1254 (
   .O(gates_1254),
   .I0(InputBits[243]),
   .I1(InputBits[306]),
   .I2(InputBits[25]),
   .I3(InputBits[472]),
   .I4(InputBits[263]),
   .I5(InputBits[401])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000110010001100000011)  
) LUT6_1255 (
   .O(gates_1255),
   .I0(InputBits[297]),
   .I1(InputBits[217]),
   .I2(InputBits[573]),
   .I3(InputBits[300]),
   .I4(InputBits[108]),
   .I5(InputBits[56])
);
LUT6 #(
   .INIT(64'b0000000000000111000010000000000000000100000011110000111000001111)  
) LUT6_1256 (
   .O(gates_1256),
   .I0(InputBits[399]),
   .I1(InputBits[260]),
   .I2(InputBits[73]),
   .I3(InputBits[519]),
   .I4(InputBits[476]),
   .I5(InputBits[255])
);
LUT6 #(
   .INIT(64'b0000000100000101000000010000010100000000000000010000000000010001)  
) LUT6_1257 (
   .O(gates_1257),
   .I0(InputBits[289]),
   .I1(InputBits[124]),
   .I2(InputBits[551]),
   .I3(InputBits[276]),
   .I4(InputBits[382]),
   .I5(InputBits[349])
);
LUT6 #(
   .INIT(64'b0000111100001000000011110000110100001111000011000000111100001101)  
) LUT6_1258 (
   .O(gates_1258),
   .I0(InputBits[158]),
   .I1(InputBits[235]),
   .I2(InputBits[4]),
   .I3(InputBits[396]),
   .I4(InputBits[111]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0000000000000001000000010100111100000000000001000000010000000111)  
) LUT6_1259 (
   .O(gates_1259),
   .I0(InputBits[250]),
   .I1(InputBits[450]),
   .I2(InputBits[266]),
   .I3(InputBits[99]),
   .I4(InputBits[504]),
   .I5(InputBits[186])
);
LUT6 #(
   .INIT(64'b0001111100001111010011110000100001001111010011110100111100001010)  
) LUT6_1260 (
   .O(gates_1260),
   .I0(InputBits[455]),
   .I1(InputBits[426]),
   .I2(InputBits[362]),
   .I3(InputBits[396]),
   .I4(InputBits[392]),
   .I5(InputBits[403])
);
LUT6 #(
   .INIT(64'b0000000000000000000100010000000100010011001100111111111100011111)  
) LUT6_1261 (
   .O(gates_1261),
   .I0(InputBits[517]),
   .I1(InputBits[119]),
   .I2(InputBits[127]),
   .I3(InputBits[245]),
   .I4(InputBits[67]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0000000000001111000000000000110100000000111110110100000111110001)  
) LUT6_1262 (
   .O(gates_1262),
   .I0(InputBits[82]),
   .I1(InputBits[304]),
   .I2(InputBits[200]),
   .I3(InputBits[314]),
   .I4(InputBits[36]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b0000000000000000001000000011001100110010001100110011000100110011)  
) LUT6_1263 (
   .O(gates_1263),
   .I0(InputBits[424]),
   .I1(InputBits[73]),
   .I2(InputBits[235]),
   .I3(InputBits[229]),
   .I4(InputBits[309]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000001101111000001110101111100000000)  
) LUT6_1264 (
   .O(gates_1264),
   .I0(InputBits[324]),
   .I1(InputBits[158]),
   .I2(InputBits[559]),
   .I3(InputBits[419]),
   .I4(InputBits[179]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000011010000011100001111)  
) LUT6_1265 (
   .O(gates_1265),
   .I0(InputBits[149]),
   .I1(InputBits[465]),
   .I2(InputBits[433]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1100101001011111011111110111111101111010010010100101101101011011)  
) LUT6_1266 (
   .O(gates_1266),
   .I0(InputBits[454]),
   .I1(InputBits[449]),
   .I2(InputBits[291]),
   .I3(InputBits[174]),
   .I4(InputBits[131]),
   .I5(InputBits[319])
);
LUT6 #(
   .INIT(64'b0000000000000001000000000000001100000000000000010000000000000010)  
) LUT6_1267 (
   .O(gates_1267),
   .I0(InputBits[550]),
   .I1(InputBits[481]),
   .I2(InputBits[99]),
   .I3(InputBits[242]),
   .I4(InputBits[14]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000010000000000000001010000010001000100)  
) LUT6_1268 (
   .O(gates_1268),
   .I0(InputBits[145]),
   .I1(InputBits[246]),
   .I2(InputBits[566]),
   .I3(InputBits[63]),
   .I4(InputBits[168]),
   .I5(InputBits[523])
);
LUT6 #(
   .INIT(64'b0000000000000000000000010000000000000000000000000001000100101011)  
) LUT6_1269 (
   .O(gates_1269),
   .I0(InputBits[42]),
   .I1(InputBits[148]),
   .I2(InputBits[81]),
   .I3(InputBits[70]),
   .I4(InputBits[410]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0000010100000101000100010000000000000001000001000000000100000100)  
) LUT6_1270 (
   .O(gates_1270),
   .I0(InputBits[481]),
   .I1(InputBits[67]),
   .I2(InputBits[469]),
   .I3(InputBits[36]),
   .I4(InputBits[412]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b0000000000010011000000110011001100000000000000110000000000011001)  
) LUT6_1271 (
   .O(gates_1271),
   .I0(InputBits[303]),
   .I1(InputBits[571]),
   .I2(InputBits[62]),
   .I3(InputBits[102]),
   .I4(InputBits[215]),
   .I5(InputBits[286])
);
LUT6 #(
   .INIT(64'b0000000000000000110100010111011100100101000000001111000111010000)  
) LUT6_1272 (
   .O(gates_1272),
   .I0(InputBits[232]),
   .I1(InputBits[174]),
   .I2(InputBits[389]),
   .I3(InputBits[324]),
   .I4(InputBits[338]),
   .I5(InputBits[190])
);
LUT6 #(
   .INIT(64'b0000000000110011001100110001001100000000001100110000011100000111)  
) LUT6_1273 (
   .O(gates_1273),
   .I0(InputBits[130]),
   .I1(InputBits[171]),
   .I2(InputBits[515]),
   .I3(InputBits[523]),
   .I4(InputBits[263]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b0000001000101010000000100011101000000000001010100010001000101011)  
) LUT6_1274 (
   .O(gates_1274),
   .I0(InputBits[397]),
   .I1(InputBits[518]),
   .I2(InputBits[36]),
   .I3(InputBits[386]),
   .I4(InputBits[446]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0000000000000000010000001101110100000000000000001000000011010000)  
) LUT6_1275 (
   .O(gates_1275),
   .I0(InputBits[135]),
   .I1(InputBits[34]),
   .I2(InputBits[422]),
   .I3(InputBits[53]),
   .I4(InputBits[507]),
   .I5(InputBits[234])
);
LUT6 #(
   .INIT(64'b0111000111111010111101111011001100111011101110101111011100111010)  
) LUT6_1276 (
   .O(gates_1276),
   .I0(InputBits[421]),
   .I1(InputBits[125]),
   .I2(InputBits[212]),
   .I3(InputBits[222]),
   .I4(InputBits[60]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0000000000000000000001010000000000000000000000000000010100000100)  
) LUT6_1277 (
   .O(gates_1277),
   .I0(InputBits[535]),
   .I1(InputBits[346]),
   .I2(InputBits[47]),
   .I3(InputBits[397]),
   .I4(InputBits[50]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0000010000000100000100010001011100000100000000100001000000000111)  
) LUT6_1278 (
   .O(gates_1278),
   .I0(InputBits[12]),
   .I1(InputBits[570]),
   .I2(InputBits[52]),
   .I3(InputBits[148]),
   .I4(InputBits[231]),
   .I5(InputBits[235])
);
LUT6 #(
   .INIT(64'b0000010101010101000000000101000000000101010101010001000001010001)  
) LUT6_1279 (
   .O(gates_1279),
   .I0(InputBits[194]),
   .I1(InputBits[541]),
   .I2(InputBits[186]),
   .I3(InputBits[127]),
   .I4(InputBits[165]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000111100001111000001110000011100000001000000110000001000000011)  
) LUT6_1280 (
   .O(gates_1280),
   .I0(InputBits[257]),
   .I1(InputBits[514]),
   .I2(InputBits[575]),
   .I3(InputBits[355]),
   .I4(InputBits[315]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0000000001010101010100000101010100000001101010100101000000110000)  
) LUT6_1281 (
   .O(gates_1281),
   .I0(InputBits[32]),
   .I1(InputBits[273]),
   .I2(InputBits[325]),
   .I3(InputBits[95]),
   .I4(InputBits[400]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0011001000010010001100110010001000110011000100010011001110100110)  
) LUT6_1282 (
   .O(gates_1282),
   .I0(InputBits[213]),
   .I1(InputBits[360]),
   .I2(InputBits[497]),
   .I3(InputBits[259]),
   .I4(InputBits[501]),
   .I5(InputBits[165])
);
LUT6 #(
   .INIT(64'b0000000101110101000000000010010100010001111111110000000000000001)  
) LUT6_1283 (
   .O(gates_1283),
   .I0(InputBits[520]),
   .I1(InputBits[54]),
   .I2(InputBits[448]),
   .I3(InputBits[535]),
   .I4(InputBits[393]),
   .I5(InputBits[376])
);
LUT6 #(
   .INIT(64'b0000000000001101000000000000111100000000000000010000000011111111)  
) LUT6_1284 (
   .O(gates_1284),
   .I0(InputBits[298]),
   .I1(InputBits[328]),
   .I2(InputBits[35]),
   .I3(InputBits[23]),
   .I4(InputBits[515]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000001010000000000000100)  
) LUT6_1285 (
   .O(gates_1285),
   .I0(InputBits[146]),
   .I1(InputBits[43]),
   .I2(InputBits[99]),
   .I3(InputBits[73]),
   .I4(InputBits[188]),
   .I5(InputBits[386])
);
LUT6 #(
   .INIT(64'b0000010100000101000001010000111100001111000011110000000101001111)  
) LUT6_1286 (
   .O(gates_1286),
   .I0(InputBits[58]),
   .I1(InputBits[428]),
   .I2(InputBits[528]),
   .I3(InputBits[226]),
   .I4(InputBits[177]),
   .I5(InputBits[67])
);
LUT6 #(
   .INIT(64'b0000000000000000000010110000111100000011000000000000111100000000)  
) LUT6_1287 (
   .O(gates_1287),
   .I0(InputBits[257]),
   .I1(InputBits[55]),
   .I2(InputBits[97]),
   .I3(InputBits[366]),
   .I4(InputBits[482]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000000000000000010001000111011100000000000000000101011001010111)  
) LUT6_1288 (
   .O(gates_1288),
   .I0(InputBits[120]),
   .I1(InputBits[454]),
   .I2(InputBits[186]),
   .I3(InputBits[426]),
   .I4(InputBits[27]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0001000000110011000000000000000000010011001100110000001000100010)  
) LUT6_1289 (
   .O(gates_1289),
   .I0(InputBits[333]),
   .I1(InputBits[25]),
   .I2(InputBits[428]),
   .I3(InputBits[206]),
   .I4(InputBits[393]),
   .I5(InputBits[54])
);
LUT6 #(
   .INIT(64'b0000111010001110000011110000111110001010100011110000111010101110)  
) LUT6_1290 (
   .O(gates_1290),
   .I0(InputBits[392]),
   .I1(InputBits[418]),
   .I2(InputBits[507]),
   .I3(InputBits[473]),
   .I4(InputBits[157]),
   .I5(InputBits[199])
);
LUT6 #(
   .INIT(64'b0000000100110111001100000011001000100010001101110011000000110011)  
) LUT6_1291 (
   .O(gates_1291),
   .I0(InputBits[284]),
   .I1(InputBits[557]),
   .I2(InputBits[316]),
   .I3(InputBits[231]),
   .I4(InputBits[443]),
   .I5(InputBits[278])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000000000000000000000101000111110001)  
) LUT6_1292 (
   .O(gates_1292),
   .I0(InputBits[460]),
   .I1(InputBits[107]),
   .I2(InputBits[335]),
   .I3(InputBits[264]),
   .I4(InputBits[97]),
   .I5(InputBits[97])
);
LUT6 #(
   .INIT(64'b0101010100000000011101010000000000110001000000000111110100010001)  
) LUT6_1293 (
   .O(gates_1293),
   .I0(InputBits[410]),
   .I1(InputBits[207]),
   .I2(InputBits[90]),
   .I3(InputBits[294]),
   .I4(InputBits[299]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000000001111000000000100011100000000000000000100000101000101)  
) LUT6_1294 (
   .O(gates_1294),
   .I0(InputBits[124]),
   .I1(InputBits[323]),
   .I2(InputBits[227]),
   .I3(InputBits[566]),
   .I4(InputBits[148]),
   .I5(InputBits[478])
);
LUT6 #(
   .INIT(64'b0000010100000001000001000000000101011111010111110001111101011011)  
) LUT6_1295 (
   .O(gates_1295),
   .I0(InputBits[214]),
   .I1(InputBits[128]),
   .I2(InputBits[70]),
   .I3(InputBits[176]),
   .I4(InputBits[341]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0000000000000000000000000000000100000000000010000000000000100011)  
) LUT6_1296 (
   .O(gates_1296),
   .I0(InputBits[320]),
   .I1(InputBits[75]),
   .I2(InputBits[490]),
   .I3(InputBits[289]),
   .I4(InputBits[99]),
   .I5(InputBits[28])
);
LUT6 #(
   .INIT(64'b1111111011000000111110101000000010100000111000001010100000000000)  
) LUT6_1297 (
   .O(gates_1297),
   .I0(gates_6),
   .I1(gates_5),
   .I2(gates_4),
   .I3(gates_3),
   .I4(gates_2),
   .I5(gates_1)
);
LUT6 #(
   .INIT(64'b1101110111111110111111001111110011011101111011001000000011110000)  
) LUT6_1298 (
   .O(gates_1298),
   .I0(gates_12),
   .I1(gates_11),
   .I2(gates_10),
   .I3(gates_9),
   .I4(gates_8),
   .I5(gates_7)
);
LUT6 #(
   .INIT(64'b1111111111111110111111111110111011110000100000001100100000001000)  
) LUT6_1299 (
   .O(gates_1299),
   .I0(gates_18),
   .I1(gates_17),
   .I2(gates_16),
   .I3(gates_15),
   .I4(gates_14),
   .I5(gates_13)
);
LUT6 #(
   .INIT(64'b1111111111111010110010001000000011101111110011001100110000000000)  
) LUT6_1300 (
   .O(gates_1300),
   .I0(gates_24),
   .I1(gates_23),
   .I2(gates_22),
   .I3(gates_21),
   .I4(gates_20),
   .I5(gates_19)
);
LUT6 #(
   .INIT(64'b1111100111101110111111111100100011111000111010001110000000000000)  
) LUT6_1301 (
   .O(gates_1301),
   .I0(gates_30),
   .I1(gates_29),
   .I2(gates_28),
   .I3(gates_27),
   .I4(gates_26),
   .I5(gates_25)
);
LUT6 #(
   .INIT(64'b1111100011111010111010001100000011111011111110101000100010000000)  
) LUT6_1302 (
   .O(gates_1302),
   .I0(gates_36),
   .I1(gates_35),
   .I2(gates_34),
   .I3(gates_33),
   .I4(gates_32),
   .I5(gates_31)
);
LUT6 #(
   .INIT(64'b1111101111111010101111111010101011111111100000001111111100000000)  
) LUT6_1303 (
   .O(gates_1303),
   .I0(gates_42),
   .I1(gates_41),
   .I2(gates_40),
   .I3(gates_39),
   .I4(gates_38),
   .I5(gates_37)
);
LUT6 #(
   .INIT(64'b1111101011111000111000001010000010100000101000000000000000000000)  
) LUT6_1304 (
   .O(gates_1304),
   .I0(gates_48),
   .I1(gates_47),
   .I2(gates_46),
   .I3(gates_45),
   .I4(gates_44),
   .I5(gates_43)
);
LUT6 #(
   .INIT(64'b1110111010000000101010001000000011101010100000000000000000000000)  
) LUT6_1305 (
   .O(gates_1305),
   .I0(gates_54),
   .I1(gates_53),
   .I2(gates_52),
   .I3(gates_51),
   .I4(gates_50),
   .I5(gates_49)
);
LUT6 #(
   .INIT(64'b1110111011111010100010001100100011101100100000001000100010000000)  
) LUT6_1306 (
   .O(gates_1306),
   .I0(gates_60),
   .I1(gates_59),
   .I2(gates_58),
   .I3(gates_57),
   .I4(gates_56),
   .I5(gates_55)
);
LUT6 #(
   .INIT(64'b1111111111111110111111111110111011111111111000001111111100000000)  
) LUT6_1307 (
   .O(gates_1307),
   .I0(gates_66),
   .I1(gates_65),
   .I2(gates_64),
   .I3(gates_63),
   .I4(gates_62),
   .I5(gates_61)
);
LUT6 #(
   .INIT(64'b1111111111111010111110101111100011111000101010001100100010000000)  
) LUT6_1308 (
   .O(gates_1308),
   .I0(gates_72),
   .I1(gates_71),
   .I2(gates_70),
   .I3(gates_69),
   .I4(gates_68),
   .I5(gates_67)
);
LUT6 #(
   .INIT(64'b1111111011101010110011101000100011001000100010000000000000000000)  
) LUT6_1309 (
   .O(gates_1309),
   .I0(gates_78),
   .I1(gates_77),
   .I2(gates_76),
   .I3(gates_75),
   .I4(gates_74),
   .I5(gates_73)
);
LUT6 #(
   .INIT(64'b1111111111111110111111111010101011111111110000001000100000000000)  
) LUT6_1310 (
   .O(gates_1310),
   .I0(gates_84),
   .I1(gates_83),
   .I2(gates_82),
   .I3(gates_81),
   .I4(gates_80),
   .I5(gates_79)
);
LUT6 #(
   .INIT(64'b1111111111111111111011001010101011111111101010101101110010000000)  
) LUT6_1311 (
   .O(gates_1311),
   .I0(gates_90),
   .I1(gates_89),
   .I2(gates_88),
   .I3(gates_87),
   .I4(gates_86),
   .I5(gates_85)
);
LUT6 #(
   .INIT(64'b1111111111111100111011101110110011101110101011001010100010001000)  
) LUT6_1312 (
   .O(gates_1312),
   .I0(gates_96),
   .I1(gates_95),
   .I2(gates_94),
   .I3(gates_93),
   .I4(gates_92),
   .I5(gates_91)
);
LUT6 #(
   .INIT(64'b1111111111111100111110101010000011111111111111101010111010001000)  
) LUT6_1313 (
   .O(gates_1313),
   .I0(gates_102),
   .I1(gates_101),
   .I2(gates_100),
   .I3(gates_99),
   .I4(gates_98),
   .I5(gates_97)
);
LUT6 #(
   .INIT(64'b1111111110001100110011100000000011101110101000001000100010000000)  
) LUT6_1314 (
   .O(gates_1314),
   .I0(gates_108),
   .I1(gates_107),
   .I2(gates_106),
   .I3(gates_105),
   .I4(gates_104),
   .I5(gates_103)
);
LUT6 #(
   .INIT(64'b1110101010101000100010000000000010101000100000000000100000000000)  
) LUT6_1315 (
   .O(gates_1315),
   .I0(gates_114),
   .I1(gates_113),
   .I2(gates_112),
   .I3(gates_111),
   .I4(gates_110),
   .I5(gates_109)
);
LUT6 #(
   .INIT(64'b1111111111111111111111101111111011111111010000101110000011000000)  
) LUT6_1316 (
   .O(gates_1316),
   .I0(gates_120),
   .I1(gates_119),
   .I2(gates_118),
   .I3(gates_117),
   .I4(gates_116),
   .I5(gates_115)
);
LUT6 #(
   .INIT(64'b1110111011111010111010001110100011101000111010001110100010001000)  
) LUT6_1317 (
   .O(gates_1317),
   .I0(gates_126),
   .I1(gates_125),
   .I2(gates_124),
   .I3(gates_123),
   .I4(gates_122),
   .I5(gates_121)
);
LUT6 #(
   .INIT(64'b1111111111101010111011100000000010111110101000101010101000000000)  
) LUT6_1318 (
   .O(gates_1318),
   .I0(gates_132),
   .I1(gates_131),
   .I2(gates_130),
   .I3(gates_129),
   .I4(gates_128),
   .I5(gates_127)
);
LUT6 #(
   .INIT(64'b1111111111111110111111111110111011111010111110101111110011101000)  
) LUT6_1319 (
   .O(gates_1319),
   .I0(gates_138),
   .I1(gates_137),
   .I2(gates_136),
   .I3(gates_135),
   .I4(gates_134),
   .I5(gates_133)
);
LUT6 #(
   .INIT(64'b1111111011111100101010001010000011101110111010001010000010100000)  
) LUT6_1320 (
   .O(gates_1320),
   .I0(gates_144),
   .I1(gates_143),
   .I2(gates_142),
   .I3(gates_141),
   .I4(gates_140),
   .I5(gates_139)
);
LUT6 #(
   .INIT(64'b1111101011101010111111111110101011111010111110001111000010000000)  
) LUT6_1321 (
   .O(gates_1321),
   .I0(gates_150),
   .I1(gates_149),
   .I2(gates_148),
   .I3(gates_147),
   .I4(gates_146),
   .I5(gates_145)
);
LUT6 #(
   .INIT(64'b1111111011111011111010001100000011111100100010001100100011001000)  
) LUT6_1322 (
   .O(gates_1322),
   .I0(gates_156),
   .I1(gates_155),
   .I2(gates_154),
   .I3(gates_153),
   .I4(gates_152),
   .I5(gates_151)
);
LUT6 #(
   .INIT(64'b1111111111111110111111110111011111111111111011001110111010000000)  
) LUT6_1323 (
   .O(gates_1323),
   .I0(gates_162),
   .I1(gates_161),
   .I2(gates_160),
   .I3(gates_159),
   .I4(gates_158),
   .I5(gates_157)
);
LUT6 #(
   .INIT(64'b1111111111111111111111001110100011101110111010000100100000000000)  
) LUT6_1324 (
   .O(gates_1324),
   .I0(gates_168),
   .I1(gates_167),
   .I2(gates_166),
   .I3(gates_165),
   .I4(gates_164),
   .I5(gates_163)
);
LUT6 #(
   .INIT(64'b1111111011111100111110101000100011111010100000001111001010000000)  
) LUT6_1325 (
   .O(gates_1325),
   .I0(gates_174),
   .I1(gates_173),
   .I2(gates_172),
   .I3(gates_171),
   .I4(gates_170),
   .I5(gates_169)
);
LUT6 #(
   .INIT(64'b1111111011111110111111101110100011011110110111001110000011001000)  
) LUT6_1326 (
   .O(gates_1326),
   .I0(gates_180),
   .I1(gates_179),
   .I2(gates_178),
   .I3(gates_177),
   .I4(gates_176),
   .I5(gates_175)
);
LUT6 #(
   .INIT(64'b1111111111111000111011001100000011110000111010001000000000001000)  
) LUT6_1327 (
   .O(gates_1327),
   .I0(gates_186),
   .I1(gates_185),
   .I2(gates_184),
   .I3(gates_183),
   .I4(gates_182),
   .I5(gates_181)
);
LUT6 #(
   .INIT(64'b1111111111111111111110101111101011111010111010101010100010000000)  
) LUT6_1328 (
   .O(gates_1328),
   .I0(gates_192),
   .I1(gates_191),
   .I2(gates_190),
   .I3(gates_189),
   .I4(gates_188),
   .I5(gates_187)
);
LUT6 #(
   .INIT(64'b1111111011111111111111101110111011111110111111101110111011101000)  
) LUT6_1329 (
   .O(gates_1329),
   .I0(gates_198),
   .I1(gates_197),
   .I2(gates_196),
   .I3(gates_195),
   .I4(gates_194),
   .I5(gates_193)
);
LUT6 #(
   .INIT(64'b1110111110011000111011101100100011001100100010001100100000000000)  
) LUT6_1330 (
   .O(gates_1330),
   .I0(gates_204),
   .I1(gates_203),
   .I2(gates_202),
   .I3(gates_201),
   .I4(gates_200),
   .I5(gates_199)
);
LUT6 #(
   .INIT(64'b1111111111111011111101111111101111110111111100100111010011100010)  
) LUT6_1331 (
   .O(gates_1331),
   .I0(gates_210),
   .I1(gates_209),
   .I2(gates_208),
   .I3(gates_207),
   .I4(gates_206),
   .I5(gates_205)
);
LUT6 #(
   .INIT(64'b1111111111110010111111101110100011101010111010101110101011001000)  
) LUT6_1332 (
   .O(gates_1332),
   .I0(gates_216),
   .I1(gates_215),
   .I2(gates_214),
   .I3(gates_213),
   .I4(gates_212),
   .I5(gates_211)
);
LUT6 #(
   .INIT(64'b1011111111111111111111111111110010111110001110000001110000000000)  
) LUT6_1333 (
   .O(gates_1333),
   .I0(gates_222),
   .I1(gates_221),
   .I2(gates_220),
   .I3(gates_219),
   .I4(gates_218),
   .I5(gates_217)
);
LUT6 #(
   .INIT(64'b1111111111111110111111111110100011111111111011001111011111001000)  
) LUT6_1334 (
   .O(gates_1334),
   .I0(gates_228),
   .I1(gates_227),
   .I2(gates_226),
   .I3(gates_225),
   .I4(gates_224),
   .I5(gates_223)
);
LUT6 #(
   .INIT(64'b1111111111111010111111001110100011101011101011101000000000000000)  
) LUT6_1335 (
   .O(gates_1335),
   .I0(gates_234),
   .I1(gates_233),
   .I2(gates_232),
   .I3(gates_231),
   .I4(gates_230),
   .I5(gates_229)
);
LUT6 #(
   .INIT(64'b1011111111111011111111111010101011111010111011101010000010000000)  
) LUT6_1336 (
   .O(gates_1336),
   .I0(gates_240),
   .I1(gates_239),
   .I2(gates_238),
   .I3(gates_237),
   .I4(gates_236),
   .I5(gates_235)
);
LUT6 #(
   .INIT(64'b1111111111101101111110100000100011111110111010001110100010000000)  
) LUT6_1337 (
   .O(gates_1337),
   .I0(gates_246),
   .I1(gates_245),
   .I2(gates_244),
   .I3(gates_243),
   .I4(gates_242),
   .I5(gates_241)
);
LUT6 #(
   .INIT(64'b1111111011100010111110101010001011111010101010101010001010100010)  
) LUT6_1338 (
   .O(gates_1338),
   .I0(gates_252),
   .I1(gates_251),
   .I2(gates_250),
   .I3(gates_249),
   .I4(gates_248),
   .I5(gates_247)
);
LUT6 #(
   .INIT(64'b1111111111111000111110001110100011111011111010001010100010001000)  
) LUT6_1339 (
   .O(gates_1339),
   .I0(gates_258),
   .I1(gates_257),
   .I2(gates_256),
   .I3(gates_255),
   .I4(gates_254),
   .I5(gates_253)
);
LUT6 #(
   .INIT(64'b1111111011101110111111101010000011111111111011101111111010100000)  
) LUT6_1340 (
   .O(gates_1340),
   .I0(gates_264),
   .I1(gates_263),
   .I2(gates_262),
   .I3(gates_261),
   .I4(gates_260),
   .I5(gates_259)
);
LUT6 #(
   .INIT(64'b1111101011100100111111111111100011111111111111111111111011001000)  
) LUT6_1341 (
   .O(gates_1341),
   .I0(gates_270),
   .I1(gates_269),
   .I2(gates_268),
   .I3(gates_267),
   .I4(gates_266),
   .I5(gates_265)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111101011111100111100001111100010101000)  
) LUT6_1342 (
   .O(gates_1342),
   .I0(gates_276),
   .I1(gates_275),
   .I2(gates_274),
   .I3(gates_273),
   .I4(gates_272),
   .I5(gates_271)
);
LUT6 #(
   .INIT(64'b1111111111111110111111011110110011001100010000001110100000000000)  
) LUT6_1343 (
   .O(gates_1343),
   .I0(gates_282),
   .I1(gates_281),
   .I2(gates_280),
   .I3(gates_279),
   .I4(gates_278),
   .I5(gates_277)
);
LUT6 #(
   .INIT(64'b1110111011101010101000000000000011101010100010001010100010000000)  
) LUT6_1344 (
   .O(gates_1344),
   .I0(gates_288),
   .I1(gates_287),
   .I2(gates_286),
   .I3(gates_285),
   .I4(gates_284),
   .I5(gates_283)
);
LUT6 #(
   .INIT(64'b1111111011101010111111101110101011111010110010001110101010101000)  
) LUT6_1345 (
   .O(gates_1345),
   .I0(gates_294),
   .I1(gates_293),
   .I2(gates_292),
   .I3(gates_291),
   .I4(gates_290),
   .I5(gates_289)
);
LUT6 #(
   .INIT(64'b1110111011111000101010101010100010101010111010001000111110000000)  
) LUT6_1346 (
   .O(gates_1346),
   .I0(gates_300),
   .I1(gates_299),
   .I2(gates_298),
   .I3(gates_297),
   .I4(gates_296),
   .I5(gates_295)
);
LUT6 #(
   .INIT(64'b1111111011101111111010001011100011101100110010001010000010100000)  
) LUT6_1347 (
   .O(gates_1347),
   .I0(gates_306),
   .I1(gates_305),
   .I2(gates_304),
   .I3(gates_303),
   .I4(gates_302),
   .I5(gates_301)
);
LUT6 #(
   .INIT(64'b1111011111110110111111111111110011110111101000001011110000000000)  
) LUT6_1348 (
   .O(gates_1348),
   .I0(gates_312),
   .I1(gates_311),
   .I2(gates_310),
   .I3(gates_309),
   .I4(gates_308),
   .I5(gates_307)
);
LUT6 #(
   .INIT(64'b1111111111111111111110011100100011111100100111001100000000000000)  
) LUT6_1349 (
   .O(gates_1349),
   .I0(gates_318),
   .I1(gates_317),
   .I2(gates_316),
   .I3(gates_315),
   .I4(gates_314),
   .I5(gates_313)
);
LUT6 #(
   .INIT(64'b1111111111111111111111101010100011101111111010001010101010001000)  
) LUT6_1350 (
   .O(gates_1350),
   .I0(gates_324),
   .I1(gates_323),
   .I2(gates_322),
   .I3(gates_321),
   .I4(gates_320),
   .I5(gates_319)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111110101011111101111000101111100000000000)  
) LUT6_1351 (
   .O(gates_1351),
   .I0(gates_330),
   .I1(gates_329),
   .I2(gates_328),
   .I3(gates_327),
   .I4(gates_326),
   .I5(gates_325)
);
LUT6 #(
   .INIT(64'b1111111011111111111011001010100011101000100000000000000000000000)  
) LUT6_1352 (
   .O(gates_1352),
   .I0(gates_336),
   .I1(gates_335),
   .I2(gates_334),
   .I3(gates_333),
   .I4(gates_332),
   .I5(gates_331)
);
LUT6 #(
   .INIT(64'b1110111011101100111111001100100011101110100011001010100010000000)  
) LUT6_1353 (
   .O(gates_1353),
   .I0(gates_342),
   .I1(gates_341),
   .I2(gates_340),
   .I3(gates_339),
   .I4(gates_338),
   .I5(gates_337)
);
LUT6 #(
   .INIT(64'b1110111011001010111010001000100011101010100010001010101010000000)  
) LUT6_1354 (
   .O(gates_1354),
   .I0(gates_348),
   .I1(gates_347),
   .I2(gates_346),
   .I3(gates_345),
   .I4(gates_344),
   .I5(gates_343)
);
LUT6 #(
   .INIT(64'b1111110111101000110111001000000011111100110000001100000000000000)  
) LUT6_1355 (
   .O(gates_1355),
   .I0(gates_354),
   .I1(gates_353),
   .I2(gates_352),
   .I3(gates_351),
   .I4(gates_350),
   .I5(gates_349)
);
LUT6 #(
   .INIT(64'b1111111011010000111110001100000011111010010110001010000000000000)  
) LUT6_1356 (
   .O(gates_1356),
   .I0(gates_360),
   .I1(gates_359),
   .I2(gates_358),
   .I3(gates_357),
   .I4(gates_356),
   .I5(gates_355)
);
LUT6 #(
   .INIT(64'b1110111010001100111010001000000011001000100000001000000000000000)  
) LUT6_1357 (
   .O(gates_1357),
   .I0(gates_366),
   .I1(gates_365),
   .I2(gates_364),
   .I3(gates_363),
   .I4(gates_362),
   .I5(gates_361)
);
LUT6 #(
   .INIT(64'b1111111111111110110101001101100011111110010110000111101001000000)  
) LUT6_1358 (
   .O(gates_1358),
   .I0(gates_372),
   .I1(gates_371),
   .I2(gates_370),
   .I3(gates_369),
   .I4(gates_368),
   .I5(gates_367)
);
LUT6 #(
   .INIT(64'b1110111011101010111111101110100011101000100000001111100010000000)  
) LUT6_1359 (
   .O(gates_1359),
   .I0(gates_378),
   .I1(gates_377),
   .I2(gates_376),
   .I3(gates_375),
   .I4(gates_374),
   .I5(gates_373)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111100011011111111111010101111111011000000)  
) LUT6_1360 (
   .O(gates_1360),
   .I0(gates_384),
   .I1(gates_383),
   .I2(gates_382),
   .I3(gates_381),
   .I4(gates_380),
   .I5(gates_379)
);
LUT6 #(
   .INIT(64'b1111111011101010111010101010101011100000000000001010000000000000)  
) LUT6_1361 (
   .O(gates_1361),
   .I0(gates_390),
   .I1(gates_389),
   .I2(gates_388),
   .I3(gates_387),
   .I4(gates_386),
   .I5(gates_385)
);
LUT6 #(
   .INIT(64'b1110101010111010100010000000100011101100100000001000000000000000)  
) LUT6_1362 (
   .O(gates_1362),
   .I0(gates_396),
   .I1(gates_395),
   .I2(gates_394),
   .I3(gates_393),
   .I4(gates_392),
   .I5(gates_391)
);
LUT6 #(
   .INIT(64'b1111111111101111111011111110100011101110111010001010101010001000)  
) LUT6_1363 (
   .O(gates_1363),
   .I0(gates_402),
   .I1(gates_401),
   .I2(gates_400),
   .I3(gates_399),
   .I4(gates_398),
   .I5(gates_397)
);
LUT6 #(
   .INIT(64'b1111110010110000111111000001000011110000001000001111000000000000)  
) LUT6_1364 (
   .O(gates_1364),
   .I0(gates_408),
   .I1(gates_407),
   .I2(gates_406),
   .I3(gates_405),
   .I4(gates_404),
   .I5(gates_403)
);
LUT6 #(
   .INIT(64'b1111111011101010111111001010111011101110101010001010110000000000)  
) LUT6_1365 (
   .O(gates_1365),
   .I0(gates_414),
   .I1(gates_413),
   .I2(gates_412),
   .I3(gates_411),
   .I4(gates_410),
   .I5(gates_409)
);
LUT6 #(
   .INIT(64'b1111111111101110111111101100110011100100010011001110101010000000)  
) LUT6_1366 (
   .O(gates_1366),
   .I0(gates_420),
   .I1(gates_419),
   .I2(gates_418),
   .I3(gates_417),
   .I4(gates_416),
   .I5(gates_415)
);
LUT6 #(
   .INIT(64'b1110111011101100111010101000101011111110111010001000100000000000)  
) LUT6_1367 (
   .O(gates_1367),
   .I0(gates_426),
   .I1(gates_425),
   .I2(gates_424),
   .I3(gates_423),
   .I4(gates_422),
   .I5(gates_421)
);
LUT6 #(
   .INIT(64'b1111101111100000111110111111000011111110111000001110100010000000)  
) LUT6_1368 (
   .O(gates_1368),
   .I0(gates_432),
   .I1(gates_431),
   .I2(gates_430),
   .I3(gates_429),
   .I4(gates_428),
   .I5(gates_427)
);
LUT6 #(
   .INIT(64'b1111111011111110111011101000000011101110000011000100000000000000)  
) LUT6_1369 (
   .O(gates_1369),
   .I0(gates_438),
   .I1(gates_437),
   .I2(gates_436),
   .I3(gates_435),
   .I4(gates_434),
   .I5(gates_433)
);
LUT6 #(
   .INIT(64'b1111111111100100111111001100010011111100110010001111010010000000)  
) LUT6_1370 (
   .O(gates_1370),
   .I0(gates_444),
   .I1(gates_443),
   .I2(gates_442),
   .I3(gates_441),
   .I4(gates_440),
   .I5(gates_439)
);
LUT6 #(
   .INIT(64'b1111111101011101111111101110000011111111010100001110100010000000)  
) LUT6_1371 (
   .O(gates_1371),
   .I0(gates_450),
   .I1(gates_449),
   .I2(gates_448),
   .I3(gates_447),
   .I4(gates_446),
   .I5(gates_445)
);
LUT6 #(
   .INIT(64'b1111111011101110111110101000101011101110110011001000100010001000)  
) LUT6_1372 (
   .O(gates_1372),
   .I0(gates_456),
   .I1(gates_455),
   .I2(gates_454),
   .I3(gates_453),
   .I4(gates_452),
   .I5(gates_451)
);
LUT6 #(
   .INIT(64'b1110100011000100111010001000000011111101101011001010100010001000)  
) LUT6_1373 (
   .O(gates_1373),
   .I0(gates_462),
   .I1(gates_461),
   .I2(gates_460),
   .I3(gates_459),
   .I4(gates_458),
   .I5(gates_457)
);
LUT6 #(
   .INIT(64'b1111111111100000111111101111100011111100111100001110100011000000)  
) LUT6_1374 (
   .O(gates_1374),
   .I0(gates_468),
   .I1(gates_467),
   .I2(gates_466),
   .I3(gates_465),
   .I4(gates_464),
   .I5(gates_463)
);
LUT6 #(
   .INIT(64'b1111110011110000111111101110111011111101110000011110111010101000)  
) LUT6_1375 (
   .O(gates_1375),
   .I0(gates_474),
   .I1(gates_473),
   .I2(gates_472),
   .I3(gates_471),
   .I4(gates_470),
   .I5(gates_469)
);
LUT6 #(
   .INIT(64'b1111111011101100111010000000000011101100111011000000100010000000)  
) LUT6_1376 (
   .O(gates_1376),
   .I0(gates_480),
   .I1(gates_479),
   .I2(gates_478),
   .I3(gates_477),
   .I4(gates_476),
   .I5(gates_475)
);
LUT6 #(
   .INIT(64'b1111111111111111111110101010101011111111111111111000100010001000)  
) LUT6_1377 (
   .O(gates_1377),
   .I0(gates_486),
   .I1(gates_485),
   .I2(gates_484),
   .I3(gates_483),
   .I4(gates_482),
   .I5(gates_481)
);
LUT6 #(
   .INIT(64'b1111111111111100111111001000100010000000100011001010100010000000)  
) LUT6_1378 (
   .O(gates_1378),
   .I0(gates_492),
   .I1(gates_491),
   .I2(gates_490),
   .I3(gates_489),
   .I4(gates_488),
   .I5(gates_487)
);
LUT6 #(
   .INIT(64'b1111111011101100111111110101111011101100101010001010110010101000)  
) LUT6_1379 (
   .O(gates_1379),
   .I0(gates_498),
   .I1(gates_497),
   .I2(gates_496),
   .I3(gates_495),
   .I4(gates_494),
   .I5(gates_493)
);
LUT6 #(
   .INIT(64'b1111111111001111111111111100110011101100101010101110000010000000)  
) LUT6_1380 (
   .O(gates_1380),
   .I0(gates_504),
   .I1(gates_503),
   .I2(gates_502),
   .I3(gates_501),
   .I4(gates_500),
   .I5(gates_499)
);
LUT6 #(
   .INIT(64'b1110100010000000101011100000000011000000000000000000000000000000)  
) LUT6_1381 (
   .O(gates_1381),
   .I0(gates_510),
   .I1(gates_509),
   .I2(gates_508),
   .I3(gates_507),
   .I4(gates_506),
   .I5(gates_505)
);
LUT6 #(
   .INIT(64'b1111111011101100111111101110100011100100000000001100100000000000)  
) LUT6_1382 (
   .O(gates_1382),
   .I0(gates_516),
   .I1(gates_515),
   .I2(gates_514),
   .I3(gates_513),
   .I4(gates_512),
   .I5(gates_511)
);
LUT6 #(
   .INIT(64'b1110111011101010110011101000101010001000111010101110100010000000)  
) LUT6_1383 (
   .O(gates_1383),
   .I0(gates_522),
   .I1(gates_521),
   .I2(gates_520),
   .I3(gates_519),
   .I4(gates_518),
   .I5(gates_517)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111100011111111101010101010101010001000)  
) LUT6_1384 (
   .O(gates_1384),
   .I0(gates_528),
   .I1(gates_527),
   .I2(gates_526),
   .I3(gates_525),
   .I4(gates_524),
   .I5(gates_523)
);
LUT6 #(
   .INIT(64'b1111111111111111111011001100100011111110110000001110100000000000)  
) LUT6_1385 (
   .O(gates_1385),
   .I0(gates_534),
   .I1(gates_533),
   .I2(gates_532),
   .I3(gates_531),
   .I4(gates_530),
   .I5(gates_529)
);
LUT6 #(
   .INIT(64'b1111110111101100111001001110010011100100100000001110000010100000)  
) LUT6_1386 (
   .O(gates_1386),
   .I0(gates_540),
   .I1(gates_539),
   .I2(gates_538),
   .I3(gates_537),
   .I4(gates_536),
   .I5(gates_535)
);
LUT6 #(
   .INIT(64'b1111111111111100111010101000000011111110101110101010101010100000)  
) LUT6_1387 (
   .O(gates_1387),
   .I0(gates_546),
   .I1(gates_545),
   .I2(gates_544),
   .I3(gates_543),
   .I4(gates_542),
   .I5(gates_541)
);
LUT6 #(
   .INIT(64'b1110111011101000111010001010100011001000110000001000000000000000)  
) LUT6_1388 (
   .O(gates_1388),
   .I0(gates_552),
   .I1(gates_551),
   .I2(gates_550),
   .I3(gates_549),
   .I4(gates_548),
   .I5(gates_547)
);
LUT6 #(
   .INIT(64'b1111111111111100111111101111100011111110110011001010100000000000)  
) LUT6_1389 (
   .O(gates_1389),
   .I0(gates_558),
   .I1(gates_557),
   .I2(gates_556),
   .I3(gates_555),
   .I4(gates_554),
   .I5(gates_553)
);
LUT6 #(
   .INIT(64'b1111111111111100110010101100100011111111111111100000101010001000)  
) LUT6_1390 (
   .O(gates_1390),
   .I0(gates_564),
   .I1(gates_563),
   .I2(gates_562),
   .I3(gates_561),
   .I4(gates_560),
   .I5(gates_559)
);
LUT6 #(
   .INIT(64'b1111111110101010111111111000100011011010100010001000100000000000)  
) LUT6_1391 (
   .O(gates_1391),
   .I0(gates_570),
   .I1(gates_569),
   .I2(gates_568),
   .I3(gates_567),
   .I4(gates_566),
   .I5(gates_565)
);
LUT6 #(
   .INIT(64'b1111111111111111111000000010000011111110111110001110000000000000)  
) LUT6_1392 (
   .O(gates_1392),
   .I0(gates_576),
   .I1(gates_575),
   .I2(gates_574),
   .I3(gates_573),
   .I4(gates_572),
   .I5(gates_571)
);
LUT6 #(
   .INIT(64'b1110111011101010111010100010000011001110100010100000000000000000)  
) LUT6_1393 (
   .O(gates_1393),
   .I0(gates_582),
   .I1(gates_581),
   .I2(gates_580),
   .I3(gates_579),
   .I4(gates_578),
   .I5(gates_577)
);
LUT6 #(
   .INIT(64'b1111111111101110111111111010111010101111111010001010110010000000)  
) LUT6_1394 (
   .O(gates_1394),
   .I0(gates_588),
   .I1(gates_587),
   .I2(gates_586),
   .I3(gates_585),
   .I4(gates_584),
   .I5(gates_583)
);
LUT6 #(
   .INIT(64'b1111111111111110111111101111111011111110111110101111010010100000)  
) LUT6_1395 (
   .O(gates_1395),
   .I0(gates_594),
   .I1(gates_593),
   .I2(gates_592),
   .I3(gates_591),
   .I4(gates_590),
   .I5(gates_589)
);
LUT6 #(
   .INIT(64'b1111111111111000111110111110100011101010101010001111000010000000)  
) LUT6_1396 (
   .O(gates_1396),
   .I0(gates_600),
   .I1(gates_599),
   .I2(gates_598),
   .I3(gates_597),
   .I4(gates_596),
   .I5(gates_595)
);
LUT6 #(
   .INIT(64'b1111111011111110111010001111000011111000111000001000000000000000)  
) LUT6_1397 (
   .O(gates_1397),
   .I0(gates_606),
   .I1(gates_605),
   .I2(gates_604),
   .I3(gates_603),
   .I4(gates_602),
   .I5(gates_601)
);
LUT6 #(
   .INIT(64'b1111111111001000111100001010000011101010101010001000100010100000)  
) LUT6_1398 (
   .O(gates_1398),
   .I0(gates_612),
   .I1(gates_611),
   .I2(gates_610),
   .I3(gates_609),
   .I4(gates_608),
   .I5(gates_607)
);
LUT6 #(
   .INIT(64'b1111111111111111111111101000000010111110011100000111000000100000)  
) LUT6_1399 (
   .O(gates_1399),
   .I0(gates_618),
   .I1(gates_617),
   .I2(gates_616),
   .I3(gates_615),
   .I4(gates_614),
   .I5(gates_613)
);
LUT6 #(
   .INIT(64'b1111111010101010111010000000000011111111111110001111100011000000)  
) LUT6_1400 (
   .O(gates_1400),
   .I0(gates_624),
   .I1(gates_623),
   .I2(gates_622),
   .I3(gates_621),
   .I4(gates_620),
   .I5(gates_619)
);
LUT6 #(
   .INIT(64'b1111111111111010111111111010001011111110101010101111100010000000)  
) LUT6_1401 (
   .O(gates_1401),
   .I0(gates_630),
   .I1(gates_629),
   .I2(gates_628),
   .I3(gates_627),
   .I4(gates_626),
   .I5(gates_625)
);
LUT6 #(
   .INIT(64'b1111111111111110000011000010100011111110111110100000000000000000)  
) LUT6_1402 (
   .O(gates_1402),
   .I0(gates_636),
   .I1(gates_635),
   .I2(gates_634),
   .I3(gates_633),
   .I4(gates_632),
   .I5(gates_631)
);
LUT6 #(
   .INIT(64'b1111111110111010111111111100111011111110111011101111111011001000)  
) LUT6_1403 (
   .O(gates_1403),
   .I0(gates_642),
   .I1(gates_641),
   .I2(gates_640),
   .I3(gates_639),
   .I4(gates_638),
   .I5(gates_637)
);
LUT6 #(
   .INIT(64'b1111111111011110111001100000000011111111101010101010000010000000)  
) LUT6_1404 (
   .O(gates_1404),
   .I0(gates_648),
   .I1(gates_647),
   .I2(gates_646),
   .I3(gates_645),
   .I4(gates_644),
   .I5(gates_643)
);
LUT6 #(
   .INIT(64'b1111111011111000111111101110100010001000010000001000000011000000)  
) LUT6_1405 (
   .O(gates_1405),
   .I0(gates_654),
   .I1(gates_653),
   .I2(gates_652),
   .I3(gates_651),
   .I4(gates_650),
   .I5(gates_649)
);
LUT6 #(
   .INIT(64'b1010111011001000101110001000000011101000100010001000100000000000)  
) LUT6_1406 (
   .O(gates_1406),
   .I0(gates_660),
   .I1(gates_659),
   .I2(gates_658),
   .I3(gates_657),
   .I4(gates_656),
   .I5(gates_655)
);
LUT6 #(
   .INIT(64'b1111111110101000111111101000000011111111100010001010000000000000)  
) LUT6_1407 (
   .O(gates_1407),
   .I0(gates_666),
   .I1(gates_665),
   .I2(gates_664),
   .I3(gates_663),
   .I4(gates_662),
   .I5(gates_661)
);
LUT6 #(
   .INIT(64'b1111111111101110111000001000100011101000110010001000000010000000)  
) LUT6_1408 (
   .O(gates_1408),
   .I0(gates_672),
   .I1(gates_671),
   .I2(gates_670),
   .I3(gates_669),
   .I4(gates_668),
   .I5(gates_667)
);
LUT6 #(
   .INIT(64'b1111111111101010111011001000100011111010100010001100100010000000)  
) LUT6_1409 (
   .O(gates_1409),
   .I0(gates_678),
   .I1(gates_677),
   .I2(gates_676),
   .I3(gates_675),
   .I4(gates_674),
   .I5(gates_673)
);
LUT6 #(
   .INIT(64'b1111111110101111111011101000101011101010001010101010101000000000)  
) LUT6_1410 (
   .O(gates_1410),
   .I0(gates_684),
   .I1(gates_683),
   .I2(gates_682),
   .I3(gates_681),
   .I4(gates_680),
   .I5(gates_679)
);
LUT6 #(
   .INIT(64'b1110111111111100111011101110000011111110111000001100110010100000)  
) LUT6_1411 (
   .O(gates_1411),
   .I0(gates_690),
   .I1(gates_689),
   .I2(gates_688),
   .I3(gates_687),
   .I4(gates_686),
   .I5(gates_685)
);
LUT6 #(
   .INIT(64'b1111111011111010111010001010000011101010111110101000000010000000)  
) LUT6_1412 (
   .O(gates_1412),
   .I0(gates_696),
   .I1(gates_695),
   .I2(gates_694),
   .I3(gates_693),
   .I4(gates_692),
   .I5(gates_691)
);
LUT6 #(
   .INIT(64'b1111111111111110111110001101100011111110100010001100100000000000)  
) LUT6_1413 (
   .O(gates_1413),
   .I0(gates_702),
   .I1(gates_701),
   .I2(gates_700),
   .I3(gates_699),
   .I4(gates_698),
   .I5(gates_697)
);
LUT6 #(
   .INIT(64'b1111111011110110111101011110000011110100110000001111010000000000)  
) LUT6_1414 (
   .O(gates_1414),
   .I0(gates_708),
   .I1(gates_707),
   .I2(gates_706),
   .I3(gates_705),
   .I4(gates_704),
   .I5(gates_703)
);
LUT6 #(
   .INIT(64'b1111111111101111111010001100100011101100110010001010000010000000)  
) LUT6_1415 (
   .O(gates_1415),
   .I0(gates_714),
   .I1(gates_713),
   .I2(gates_712),
   .I3(gates_711),
   .I4(gates_710),
   .I5(gates_709)
);
LUT6 #(
   .INIT(64'b1111111110111101111111111010111010011101000000001010001000000000)  
) LUT6_1416 (
   .O(gates_1416),
   .I0(gates_720),
   .I1(gates_719),
   .I2(gates_718),
   .I3(gates_717),
   .I4(gates_716),
   .I5(gates_715)
);
LUT6 #(
   .INIT(64'b1111111011111110111111001110100011111100111010001110110010000000)  
) LUT6_1417 (
   .O(gates_1417),
   .I0(gates_726),
   .I1(gates_725),
   .I2(gates_724),
   .I3(gates_723),
   .I4(gates_722),
   .I5(gates_721)
);
LUT6 #(
   .INIT(64'b1111111011101010111110001000100011111010101000101111100000000000)  
) LUT6_1418 (
   .O(gates_1418),
   .I0(gates_732),
   .I1(gates_731),
   .I2(gates_730),
   .I3(gates_729),
   .I4(gates_728),
   .I5(gates_727)
);
LUT6 #(
   .INIT(64'b1111111111111011111111111111111011111110111010101110101010101010)  
) LUT6_1419 (
   .O(gates_1419),
   .I0(gates_738),
   .I1(gates_737),
   .I2(gates_736),
   .I3(gates_735),
   .I4(gates_734),
   .I5(gates_733)
);
LUT6 #(
   .INIT(64'b1111111111111111000000111000100011111111111010000000000000001000)  
) LUT6_1420 (
   .O(gates_1420),
   .I0(gates_744),
   .I1(gates_743),
   .I2(gates_742),
   .I3(gates_741),
   .I4(gates_740),
   .I5(gates_739)
);
LUT6 #(
   .INIT(64'b1111111011111110111010001100000011111010101010001000000000000000)  
) LUT6_1421 (
   .O(gates_1421),
   .I0(gates_750),
   .I1(gates_749),
   .I2(gates_748),
   .I3(gates_747),
   .I4(gates_746),
   .I5(gates_745)
);
LUT6 #(
   .INIT(64'b1111111111111010101110110000000011111010111000000110000000000000)  
) LUT6_1422 (
   .O(gates_1422),
   .I0(gates_756),
   .I1(gates_755),
   .I2(gates_754),
   .I3(gates_753),
   .I4(gates_752),
   .I5(gates_751)
);
LUT6 #(
   .INIT(64'b1111111111111010111110111010100011111011101010101000101010000000)  
) LUT6_1423 (
   .O(gates_1423),
   .I0(gates_762),
   .I1(gates_761),
   .I2(gates_760),
   .I3(gates_759),
   .I4(gates_758),
   .I5(gates_757)
);
LUT6 #(
   .INIT(64'b1111111011111000111111011100100011101000100000001010101000000000)  
) LUT6_1424 (
   .O(gates_1424),
   .I0(gates_768),
   .I1(gates_767),
   .I2(gates_766),
   .I3(gates_765),
   .I4(gates_764),
   .I5(gates_763)
);
LUT6 #(
   .INIT(64'b1111111111101101111011111111111011111111111111111111111101001000)  
) LUT6_1425 (
   .O(gates_1425),
   .I0(gates_774),
   .I1(gates_773),
   .I2(gates_772),
   .I3(gates_771),
   .I4(gates_770),
   .I5(gates_769)
);
LUT6 #(
   .INIT(64'b1111111111111100111110101000100010100000100010000000000000000000)  
) LUT6_1426 (
   .O(gates_1426),
   .I0(gates_780),
   .I1(gates_779),
   .I2(gates_778),
   .I3(gates_777),
   .I4(gates_776),
   .I5(gates_775)
);
LUT6 #(
   .INIT(64'b1111111011101110111011101010100011011110111010001110110010000000)  
) LUT6_1427 (
   .O(gates_1427),
   .I0(gates_786),
   .I1(gates_785),
   .I2(gates_784),
   .I3(gates_783),
   .I4(gates_782),
   .I5(gates_781)
);
LUT6 #(
   .INIT(64'b1111111111111110111110111111000011111110111011100011000100000000)  
) LUT6_1428 (
   .O(gates_1428),
   .I0(gates_792),
   .I1(gates_791),
   .I2(gates_790),
   .I3(gates_789),
   .I4(gates_788),
   .I5(gates_787)
);
LUT6 #(
   .INIT(64'b1111111110100010111110101010001011101010101010001110101000100000)  
) LUT6_1429 (
   .O(gates_1429),
   .I0(gates_798),
   .I1(gates_797),
   .I2(gates_796),
   .I3(gates_795),
   .I4(gates_794),
   .I5(gates_793)
);
LUT6 #(
   .INIT(64'b1111111110101010111111101011100011111111111000001111101010100000)  
) LUT6_1430 (
   .O(gates_1430),
   .I0(gates_804),
   .I1(gates_803),
   .I2(gates_802),
   .I3(gates_801),
   .I4(gates_800),
   .I5(gates_799)
);
LUT6 #(
   .INIT(64'b1111111111111000110010001110000011101110110100001100000011000000)  
) LUT6_1431 (
   .O(gates_1431),
   .I0(gates_810),
   .I1(gates_809),
   .I2(gates_808),
   .I3(gates_807),
   .I4(gates_806),
   .I5(gates_805)
);
LUT6 #(
   .INIT(64'b1111111110101000111111100001000011111110000000001110100000000000)  
) LUT6_1432 (
   .O(gates_1432),
   .I0(gates_816),
   .I1(gates_815),
   .I2(gates_814),
   .I3(gates_813),
   .I4(gates_812),
   .I5(gates_811)
);
LUT6 #(
   .INIT(64'b1111101010110000111110001110000011111101111100101110000000000000)  
) LUT6_1433 (
   .O(gates_1433),
   .I0(gates_822),
   .I1(gates_821),
   .I2(gates_820),
   .I3(gates_819),
   .I4(gates_818),
   .I5(gates_817)
);
LUT6 #(
   .INIT(64'b1111111010101110111011001010100010111110101011001010100010000000)  
) LUT6_1434 (
   .O(gates_1434),
   .I0(gates_828),
   .I1(gates_827),
   .I2(gates_826),
   .I3(gates_825),
   .I4(gates_824),
   .I5(gates_823)
);
LUT6 #(
   .INIT(64'b1111111011111010111111000111100011111100110100001101000001010000)  
) LUT6_1435 (
   .O(gates_1435),
   .I0(gates_834),
   .I1(gates_833),
   .I2(gates_832),
   .I3(gates_831),
   .I4(gates_830),
   .I5(gates_829)
);
LUT6 #(
   .INIT(64'b1111111011101000101100100010000011101010111000001010000011101000)  
) LUT6_1436 (
   .O(gates_1436),
   .I0(gates_840),
   .I1(gates_839),
   .I2(gates_838),
   .I3(gates_837),
   .I4(gates_836),
   .I5(gates_835)
);
LUT6 #(
   .INIT(64'b1111110111110000111111101110100010101000100010001010101010000000)  
) LUT6_1437 (
   .O(gates_1437),
   .I0(gates_846),
   .I1(gates_845),
   .I2(gates_844),
   .I3(gates_843),
   .I4(gates_842),
   .I5(gates_841)
);
LUT6 #(
   .INIT(64'b1111111100110111111111100011000011111110111010001110110000000000)  
) LUT6_1438 (
   .O(gates_1438),
   .I0(gates_852),
   .I1(gates_851),
   .I2(gates_850),
   .I3(gates_849),
   .I4(gates_848),
   .I5(gates_847)
);
LUT6 #(
   .INIT(64'b1111111011101110111111101010111011111110111010101110000010000000)  
) LUT6_1439 (
   .O(gates_1439),
   .I0(gates_858),
   .I1(gates_857),
   .I2(gates_856),
   .I3(gates_855),
   .I4(gates_854),
   .I5(gates_853)
);
LUT6 #(
   .INIT(64'b1111111111101100111111101110100011111100110011001110100000000000)  
) LUT6_1440 (
   .O(gates_1440),
   .I0(gates_864),
   .I1(gates_863),
   .I2(gates_862),
   .I3(gates_861),
   .I4(gates_860),
   .I5(gates_859)
);
LUT6 #(
   .INIT(64'b1100110011101100111110011111110011000000110010001110001011100000)  
) LUT6_1441 (
   .O(gates_1441),
   .I0(gates_870),
   .I1(gates_869),
   .I2(gates_868),
   .I3(gates_867),
   .I4(gates_866),
   .I5(gates_865)
);
LUT6 #(
   .INIT(64'b1111111111111110111101001100000011111110110010001010100000000000)  
) LUT6_1442 (
   .O(gates_1442),
   .I0(gates_876),
   .I1(gates_875),
   .I2(gates_874),
   .I3(gates_873),
   .I4(gates_872),
   .I5(gates_871)
);
LUT6 #(
   .INIT(64'b1111111110111011111111111010001011110000100000001010000000000000)  
) LUT6_1443 (
   .O(gates_1443),
   .I0(gates_882),
   .I1(gates_881),
   .I2(gates_880),
   .I3(gates_879),
   .I4(gates_878),
   .I5(gates_877)
);
LUT6 #(
   .INIT(64'b1111111011101000111011001110010011001000100000001100000010000000)  
) LUT6_1444 (
   .O(gates_1444),
   .I0(gates_888),
   .I1(gates_887),
   .I2(gates_886),
   .I3(gates_885),
   .I4(gates_884),
   .I5(gates_883)
);
LUT6 #(
   .INIT(64'b1111111110101010010011010000000011111100100000000100100000000000)  
) LUT6_1445 (
   .O(gates_1445),
   .I0(gates_894),
   .I1(gates_893),
   .I2(gates_892),
   .I3(gates_891),
   .I4(gates_890),
   .I5(gates_889)
);
LUT6 #(
   .INIT(64'b1111111011111100110001001000000011001000100010001000000010000000)  
) LUT6_1446 (
   .O(gates_1446),
   .I0(gates_900),
   .I1(gates_899),
   .I2(gates_898),
   .I3(gates_897),
   .I4(gates_896),
   .I5(gates_895)
);
LUT6 #(
   .INIT(64'b1111101011111010111011001110100011101000101010000000000000000000)  
) LUT6_1447 (
   .O(gates_1447),
   .I0(gates_906),
   .I1(gates_905),
   .I2(gates_904),
   .I3(gates_903),
   .I4(gates_902),
   .I5(gates_901)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111010011111111111111101110101011100000)  
) LUT6_1448 (
   .O(gates_1448),
   .I0(gates_912),
   .I1(gates_911),
   .I2(gates_910),
   .I3(gates_909),
   .I4(gates_908),
   .I5(gates_907)
);
LUT6 #(
   .INIT(64'b1111111111111010111111101110101011111111111110111110101010101010)  
) LUT6_1449 (
   .O(gates_1449),
   .I0(gates_918),
   .I1(gates_917),
   .I2(gates_916),
   .I3(gates_915),
   .I4(gates_914),
   .I5(gates_913)
);
LUT6 #(
   .INIT(64'b1111111111111110000111010000100011101111111010100000110000001000)  
) LUT6_1450 (
   .O(gates_1450),
   .I0(gates_924),
   .I1(gates_923),
   .I2(gates_922),
   .I3(gates_921),
   .I4(gates_920),
   .I5(gates_919)
);
LUT6 #(
   .INIT(64'b1111111111111000111111101100100011111111111110001110111000000000)  
) LUT6_1451 (
   .O(gates_1451),
   .I0(gates_930),
   .I1(gates_929),
   .I2(gates_928),
   .I3(gates_927),
   .I4(gates_926),
   .I5(gates_925)
);
LUT6 #(
   .INIT(64'b1111111011111100101010000000000011101010111111001010000000000000)  
) LUT6_1452 (
   .O(gates_1452),
   .I0(gates_936),
   .I1(gates_935),
   .I2(gates_934),
   .I3(gates_933),
   .I4(gates_932),
   .I5(gates_931)
);
LUT6 #(
   .INIT(64'b1111110011100000110011000000000011011000101000000100000000000000)  
) LUT6_1453 (
   .O(gates_1453),
   .I0(gates_942),
   .I1(gates_941),
   .I2(gates_940),
   .I3(gates_939),
   .I4(gates_938),
   .I5(gates_937)
);
LUT6 #(
   .INIT(64'b1111111111111111111110001000100011111111111111001010000000000000)  
) LUT6_1454 (
   .O(gates_1454),
   .I0(gates_948),
   .I1(gates_947),
   .I2(gates_946),
   .I3(gates_945),
   .I4(gates_944),
   .I5(gates_943)
);
LUT6 #(
   .INIT(64'b1111111010101010111011001110100011111000100000001111100011100000)  
) LUT6_1455 (
   .O(gates_1455),
   .I0(gates_954),
   .I1(gates_953),
   .I2(gates_952),
   .I3(gates_951),
   .I4(gates_950),
   .I5(gates_949)
);
LUT6 #(
   .INIT(64'b1111111011101110111111001110100010101010111000101110000010000000)  
) LUT6_1456 (
   .O(gates_1456),
   .I0(gates_960),
   .I1(gates_959),
   .I2(gates_958),
   .I3(gates_957),
   .I4(gates_956),
   .I5(gates_955)
);
LUT6 #(
   .INIT(64'b1111111011101110101010101000100011111010101010001010001010000000)  
) LUT6_1457 (
   .O(gates_1457),
   .I0(gates_966),
   .I1(gates_965),
   .I2(gates_964),
   .I3(gates_963),
   .I4(gates_962),
   .I5(gates_961)
);
LUT6 #(
   .INIT(64'b1111111110111110111110101111101011111110101010001011110010101000)  
) LUT6_1458 (
   .O(gates_1458),
   .I0(gates_972),
   .I1(gates_971),
   .I2(gates_970),
   .I3(gates_969),
   .I4(gates_968),
   .I5(gates_967)
);
LUT6 #(
   .INIT(64'b1011101010110000101010001000000010111000100010001000100010000000)  
) LUT6_1459 (
   .O(gates_1459),
   .I0(gates_978),
   .I1(gates_977),
   .I2(gates_976),
   .I3(gates_975),
   .I4(gates_974),
   .I5(gates_973)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111110011110010011000001110000010001100)  
) LUT6_1460 (
   .O(gates_1460),
   .I0(gates_984),
   .I1(gates_983),
   .I2(gates_982),
   .I3(gates_981),
   .I4(gates_980),
   .I5(gates_979)
);
LUT6 #(
   .INIT(64'b1111101010100000111110001010000011100000000000001010000000000000)  
) LUT6_1461 (
   .O(gates_1461),
   .I0(gates_990),
   .I1(gates_989),
   .I2(gates_988),
   .I3(gates_987),
   .I4(gates_986),
   .I5(gates_985)
);
LUT6 #(
   .INIT(64'b1111111011111010111011101010000011001000110010001110101000000000)  
) LUT6_1462 (
   .O(gates_1462),
   .I0(gates_996),
   .I1(gates_995),
   .I2(gates_994),
   .I3(gates_993),
   .I4(gates_992),
   .I5(gates_991)
);
LUT6 #(
   .INIT(64'b1111111011001100111010001100110011001000000000000000000000000000)  
) LUT6_1463 (
   .O(gates_1463),
   .I0(gates_1002),
   .I1(gates_1001),
   .I2(gates_1000),
   .I3(gates_999),
   .I4(gates_998),
   .I5(gates_997)
);
LUT6 #(
   .INIT(64'b1111110011111000111010001000000011101110111110001000000010000000)  
) LUT6_1464 (
   .O(gates_1464),
   .I0(gates_1008),
   .I1(gates_1007),
   .I2(gates_1006),
   .I3(gates_1005),
   .I4(gates_1004),
   .I5(gates_1003)
);
LUT6 #(
   .INIT(64'b1111111111111010111111111111101011101110111010001111111011100000)  
) LUT6_1465 (
   .O(gates_1465),
   .I0(gates_1014),
   .I1(gates_1013),
   .I2(gates_1012),
   .I3(gates_1011),
   .I4(gates_1010),
   .I5(gates_1009)
);
LUT6 #(
   .INIT(64'b1110111111101010111010101110101011111110101011001110110010101000)  
) LUT6_1466 (
   .O(gates_1466),
   .I0(gates_1020),
   .I1(gates_1019),
   .I2(gates_1018),
   .I3(gates_1017),
   .I4(gates_1016),
   .I5(gates_1015)
);
LUT6 #(
   .INIT(64'b1110111010101010110010001000100011000100001000000000000000000000)  
) LUT6_1467 (
   .O(gates_1467),
   .I0(gates_1026),
   .I1(gates_1025),
   .I2(gates_1024),
   .I3(gates_1023),
   .I4(gates_1022),
   .I5(gates_1021)
);
LUT6 #(
   .INIT(64'b1111111011000000110111001100000011111000100000001111100011000000)  
) LUT6_1468 (
   .O(gates_1468),
   .I0(gates_1032),
   .I1(gates_1031),
   .I2(gates_1030),
   .I3(gates_1029),
   .I4(gates_1028),
   .I5(gates_1027)
);
LUT6 #(
   .INIT(64'b1111111011101110111010001100100011101010000000000000000000000000)  
) LUT6_1469 (
   .O(gates_1469),
   .I0(gates_1038),
   .I1(gates_1037),
   .I2(gates_1036),
   .I3(gates_1035),
   .I4(gates_1034),
   .I5(gates_1033)
);
LUT6 #(
   .INIT(64'b1110101010101000101010101000000010101000100000000000000000000000)  
) LUT6_1470 (
   .O(gates_1470),
   .I0(gates_1044),
   .I1(gates_1043),
   .I2(gates_1042),
   .I3(gates_1041),
   .I4(gates_1040),
   .I5(gates_1039)
);
LUT6 #(
   .INIT(64'b1111111111101010111111101110100011100000110010001110111000000000)  
) LUT6_1471 (
   .O(gates_1471),
   .I0(gates_1050),
   .I1(gates_1049),
   .I2(gates_1048),
   .I3(gates_1047),
   .I4(gates_1046),
   .I5(gates_1045)
);
LUT6 #(
   .INIT(64'b1111110010101000111110000000000011101000000000001110000000000000)  
) LUT6_1472 (
   .O(gates_1472),
   .I0(gates_1056),
   .I1(gates_1055),
   .I2(gates_1054),
   .I3(gates_1053),
   .I4(gates_1052),
   .I5(gates_1051)
);
LUT6 #(
   .INIT(64'b1111101100111011101011100011101011101111001000100010111000101000)  
) LUT6_1473 (
   .O(gates_1473),
   .I0(gates_1062),
   .I1(gates_1061),
   .I2(gates_1060),
   .I3(gates_1059),
   .I4(gates_1058),
   .I5(gates_1057)
);
LUT6 #(
   .INIT(64'b1111111011111111111010001000100011111010111110101111000000000000)  
) LUT6_1474 (
   .O(gates_1474),
   .I0(gates_1068),
   .I1(gates_1067),
   .I2(gates_1066),
   .I3(gates_1065),
   .I4(gates_1064),
   .I5(gates_1063)
);
LUT6 #(
   .INIT(64'b1111111111011111111111111111111111011111111111001111111111000100)  
) LUT6_1475 (
   .O(gates_1475),
   .I0(gates_1074),
   .I1(gates_1073),
   .I2(gates_1072),
   .I3(gates_1071),
   .I4(gates_1070),
   .I5(gates_1069)
);
LUT6 #(
   .INIT(64'b1010100011101000100000001000000010101000101000000000000000000000)  
) LUT6_1476 (
   .O(gates_1476),
   .I0(gates_1080),
   .I1(gates_1079),
   .I2(gates_1078),
   .I3(gates_1077),
   .I4(gates_1076),
   .I5(gates_1075)
);
LUT6 #(
   .INIT(64'b1110111011101111111011101010101011001010111010001110110010000000)  
) LUT6_1477 (
   .O(gates_1477),
   .I0(gates_1086),
   .I1(gates_1085),
   .I2(gates_1084),
   .I3(gates_1083),
   .I4(gates_1082),
   .I5(gates_1081)
);
LUT6 #(
   .INIT(64'b1111111111111100111111111010100011111111101010001010111010000000)  
) LUT6_1478 (
   .O(gates_1478),
   .I0(gates_1092),
   .I1(gates_1091),
   .I2(gates_1090),
   .I3(gates_1089),
   .I4(gates_1088),
   .I5(gates_1087)
);
LUT6 #(
   .INIT(64'b1111101011101100011000100010000010101100101010001010000000101000)  
) LUT6_1479 (
   .O(gates_1479),
   .I0(gates_1098),
   .I1(gates_1097),
   .I2(gates_1096),
   .I3(gates_1095),
   .I4(gates_1094),
   .I5(gates_1093)
);
LUT6 #(
   .INIT(64'b1110111011101000110010001010001010101000100010000000000000000000)  
) LUT6_1480 (
   .O(gates_1480),
   .I0(gates_1104),
   .I1(gates_1103),
   .I2(gates_1102),
   .I3(gates_1101),
   .I4(gates_1100),
   .I5(gates_1099)
);
LUT6 #(
   .INIT(64'b1111111111111111111111101100100011001100100010000000000000000000)  
) LUT6_1481 (
   .O(gates_1481),
   .I0(gates_1110),
   .I1(gates_1109),
   .I2(gates_1108),
   .I3(gates_1107),
   .I4(gates_1106),
   .I5(gates_1105)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111110011111110111010001111101011001000)  
) LUT6_1482 (
   .O(gates_1482),
   .I0(gates_1116),
   .I1(gates_1115),
   .I2(gates_1114),
   .I3(gates_1113),
   .I4(gates_1112),
   .I5(gates_1111)
);
LUT6 #(
   .INIT(64'b1110111011101100100010000000000011001000110000000000000000000000)  
) LUT6_1483 (
   .O(gates_1483),
   .I0(gates_1122),
   .I1(gates_1121),
   .I2(gates_1120),
   .I3(gates_1119),
   .I4(gates_1118),
   .I5(gates_1117)
);
LUT6 #(
   .INIT(64'b1111111111111100101100001000000011111111111111100010000000000000)  
) LUT6_1484 (
   .O(gates_1484),
   .I0(gates_1128),
   .I1(gates_1127),
   .I2(gates_1126),
   .I3(gates_1125),
   .I4(gates_1124),
   .I5(gates_1123)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111110011111111111110101111100011101000)  
) LUT6_1485 (
   .O(gates_1485),
   .I0(gates_1134),
   .I1(gates_1133),
   .I2(gates_1132),
   .I3(gates_1131),
   .I4(gates_1130),
   .I5(gates_1129)
);
LUT6 #(
   .INIT(64'b1111111111110010111011000000000011111110100000101100000000000000)  
) LUT6_1486 (
   .O(gates_1486),
   .I0(gates_1140),
   .I1(gates_1139),
   .I2(gates_1138),
   .I3(gates_1137),
   .I4(gates_1136),
   .I5(gates_1135)
);
LUT6 #(
   .INIT(64'b1110101011000100111011001110000011010000100000001100000000000000)  
) LUT6_1487 (
   .O(gates_1487),
   .I0(gates_1146),
   .I1(gates_1145),
   .I2(gates_1144),
   .I3(gates_1143),
   .I4(gates_1142),
   .I5(gates_1141)
);
LUT6 #(
   .INIT(64'b1111111011111000101100001101000011111110111010001110100010000000)  
) LUT6_1488 (
   .O(gates_1488),
   .I0(gates_1152),
   .I1(gates_1151),
   .I2(gates_1150),
   .I3(gates_1149),
   .I4(gates_1148),
   .I5(gates_1147)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111111100011101100101001101010110010101000)  
) LUT6_1489 (
   .O(gates_1489),
   .I0(gates_1158),
   .I1(gates_1157),
   .I2(gates_1156),
   .I3(gates_1155),
   .I4(gates_1154),
   .I5(gates_1153)
);
LUT6 #(
   .INIT(64'b1111111111111110111111101110110011110110111011001111110011101000)  
) LUT6_1490 (
   .O(gates_1490),
   .I0(gates_1164),
   .I1(gates_1163),
   .I2(gates_1162),
   .I3(gates_1161),
   .I4(gates_1160),
   .I5(gates_1159)
);
LUT6 #(
   .INIT(64'b1111111111111111111111111101000011011111110010001101110000000000)  
) LUT6_1491 (
   .O(gates_1491),
   .I0(gates_1170),
   .I1(gates_1169),
   .I2(gates_1168),
   .I3(gates_1167),
   .I4(gates_1166),
   .I5(gates_1165)
);
LUT6 #(
   .INIT(64'b1111111111111110111111001011110011111110101010001110100000001000)  
) LUT6_1492 (
   .O(gates_1492),
   .I0(gates_1176),
   .I1(gates_1175),
   .I2(gates_1174),
   .I3(gates_1173),
   .I4(gates_1172),
   .I5(gates_1171)
);
LUT6 #(
   .INIT(64'b1111111111111101100010000000000010111100100000001010100000000000)  
) LUT6_1493 (
   .O(gates_1493),
   .I0(gates_1182),
   .I1(gates_1181),
   .I2(gates_1180),
   .I3(gates_1179),
   .I4(gates_1178),
   .I5(gates_1177)
);
LUT6 #(
   .INIT(64'b1111111111101110111011101110100011111110101000001110110011001000)  
) LUT6_1494 (
   .O(gates_1494),
   .I0(gates_1188),
   .I1(gates_1187),
   .I2(gates_1186),
   .I3(gates_1185),
   .I4(gates_1184),
   .I5(gates_1183)
);
LUT6 #(
   .INIT(64'b1111111010101000111110101000000011111000101000001110000000000000)  
) LUT6_1495 (
   .O(gates_1495),
   .I0(gates_1194),
   .I1(gates_1193),
   .I2(gates_1192),
   .I3(gates_1191),
   .I4(gates_1190),
   .I5(gates_1189)
);
LUT6 #(
   .INIT(64'b1111111111111110111111101111111011111111111111100100110001000100)  
) LUT6_1496 (
   .O(gates_1496),
   .I0(gates_1200),
   .I1(gates_1199),
   .I2(gates_1198),
   .I3(gates_1197),
   .I4(gates_1196),
   .I5(gates_1195)
);
LUT6 #(
   .INIT(64'b1111111011111100111111001111110011101100110111001100110011001100)  
) LUT6_1497 (
   .O(gates_1497),
   .I0(gates_1206),
   .I1(gates_1205),
   .I2(gates_1204),
   .I3(gates_1203),
   .I4(gates_1202),
   .I5(gates_1201)
);
LUT6 #(
   .INIT(64'b1111110111111110111111001111000011111100111110001101100011110000)  
) LUT6_1498 (
   .O(gates_1498),
   .I0(gates_1212),
   .I1(gates_1211),
   .I2(gates_1210),
   .I3(gates_1209),
   .I4(gates_1208),
   .I5(gates_1207)
);
LUT6 #(
   .INIT(64'b1111111111111110111100111111000010000000110011000000000000000000)  
) LUT6_1499 (
   .O(gates_1499),
   .I0(gates_1218),
   .I1(gates_1217),
   .I2(gates_1216),
   .I3(gates_1215),
   .I4(gates_1214),
   .I5(gates_1213)
);
LUT6 #(
   .INIT(64'b1111110011110000100010000000000011110100111000000000000000000000)  
) LUT6_1500 (
   .O(gates_1500),
   .I0(gates_1224),
   .I1(gates_1223),
   .I2(gates_1222),
   .I3(gates_1221),
   .I4(gates_1220),
   .I5(gates_1219)
);
LUT6 #(
   .INIT(64'b1111001011100000101000001000100010100000100000000000000000000000)  
) LUT6_1501 (
   .O(gates_1501),
   .I0(gates_1230),
   .I1(gates_1229),
   .I2(gates_1228),
   .I3(gates_1227),
   .I4(gates_1226),
   .I5(gates_1225)
);
LUT6 #(
   .INIT(64'b1111100011111000111110001010000011111010101010001110000010100000)  
) LUT6_1502 (
   .O(gates_1502),
   .I0(gates_1236),
   .I1(gates_1235),
   .I2(gates_1234),
   .I3(gates_1233),
   .I4(gates_1232),
   .I5(gates_1231)
);
LUT6 #(
   .INIT(64'b1111111111101111111011001100110011001111100011001000110010001100)  
) LUT6_1503 (
   .O(gates_1503),
   .I0(gates_1242),
   .I1(gates_1241),
   .I2(gates_1240),
   .I3(gates_1239),
   .I4(gates_1238),
   .I5(gates_1237)
);
LUT6 #(
   .INIT(64'b1111111011111110111111101111111011111100111010001110110010101000)  
) LUT6_1504 (
   .O(gates_1504),
   .I0(gates_1248),
   .I1(gates_1247),
   .I2(gates_1246),
   .I3(gates_1245),
   .I4(gates_1244),
   .I5(gates_1243)
);
LUT6 #(
   .INIT(64'b1111111111001100110000001000000011101000110000001000000010000000)  
) LUT6_1505 (
   .O(gates_1505),
   .I0(gates_1254),
   .I1(gates_1253),
   .I2(gates_1252),
   .I3(gates_1251),
   .I4(gates_1250),
   .I5(gates_1249)
);
LUT6 #(
   .INIT(64'b1110111011101000110010000000000011001010100010001000100000000000)  
) LUT6_1506 (
   .O(gates_1506),
   .I0(gates_1260),
   .I1(gates_1259),
   .I2(gates_1258),
   .I3(gates_1257),
   .I4(gates_1256),
   .I5(gates_1255)
);
LUT6 #(
   .INIT(64'b1110100011100000110010001100000010001000000000001000000000000000)  
) LUT6_1507 (
   .O(gates_1507),
   .I0(gates_1266),
   .I1(gates_1265),
   .I2(gates_1264),
   .I3(gates_1263),
   .I4(gates_1262),
   .I5(gates_1261)
);
LUT6 #(
   .INIT(64'b1011111111011111111111111111101011111111011011111111111111111000)  
) LUT6_1508 (
   .O(gates_1508),
   .I0(gates_1272),
   .I1(gates_1271),
   .I2(gates_1270),
   .I3(gates_1269),
   .I4(gates_1268),
   .I5(gates_1267)
);
LUT6 #(
   .INIT(64'b1111111111111111111011101110110011101010111010001010110000100000)  
) LUT6_1509 (
   .O(gates_1509),
   .I0(gates_1278),
   .I1(gates_1277),
   .I2(gates_1276),
   .I3(gates_1275),
   .I4(gates_1274),
   .I5(gates_1273)
);
LUT6 #(
   .INIT(64'b1111111011111100111011001110000010101100111010001100100011000000)  
) LUT6_1510 (
   .O(gates_1510),
   .I0(gates_1284),
   .I1(gates_1283),
   .I2(gates_1282),
   .I3(gates_1281),
   .I4(gates_1280),
   .I5(gates_1279)
);
LUT6 #(
   .INIT(64'b1111111111101100110101010000000011111110111010001100010000000000)  
) LUT6_1511 (
   .O(gates_1511),
   .I0(gates_1290),
   .I1(gates_1289),
   .I2(gates_1288),
   .I3(gates_1287),
   .I4(gates_1286),
   .I5(gates_1285)
);
LUT6 #(
   .INIT(64'b1111110011101000111111011000000010101000100010001000100000000000)  
) LUT6_1512 (
   .O(gates_1512),
   .I0(gates_1296),
   .I1(gates_1295),
   .I2(gates_1294),
   .I3(gates_1293),
   .I4(gates_1292),
   .I5(gates_1291)
);
LUT6 #(
   .INIT(64'b1111111111101110111111111100000011101010100010001100000000000000)  
) LUT6_1513 (
   .O(gates_1513),
   .I0(gates_1302),
   .I1(gates_1301),
   .I2(gates_1300),
   .I3(gates_1299),
   .I4(gates_1298),
   .I5(gates_1297)
);
LUT6 #(
   .INIT(64'b1111111111111110111010100100100011111010111010001000100010000000)  
) LUT6_1514 (
   .O(gates_1514),
   .I0(gates_1308),
   .I1(gates_1307),
   .I2(gates_1306),
   .I3(gates_1305),
   .I4(gates_1304),
   .I5(gates_1303)
);
LUT6 #(
   .INIT(64'b1111101011100000111001001100000011100010100000001000000010000000)  
) LUT6_1515 (
   .O(gates_1515),
   .I0(gates_1314),
   .I1(gates_1313),
   .I2(gates_1312),
   .I3(gates_1311),
   .I4(gates_1310),
   .I5(gates_1309)
);
LUT6 #(
   .INIT(64'b1111111110001000111111001000000011101100100010001010000010000000)  
) LUT6_1516 (
   .O(gates_1516),
   .I0(gates_1320),
   .I1(gates_1319),
   .I2(gates_1318),
   .I3(gates_1317),
   .I4(gates_1316),
   .I5(gates_1315)
);
LUT6 #(
   .INIT(64'b1111110111111100111010001110100011110000000000001000000010000000)  
) LUT6_1517 (
   .O(gates_1517),
   .I0(gates_1326),
   .I1(gates_1325),
   .I2(gates_1324),
   .I3(gates_1323),
   .I4(gates_1322),
   .I5(gates_1321)
);
LUT6 #(
   .INIT(64'b1111111011100000111110101000000011101010001010001011000010000000)  
) LUT6_1518 (
   .O(gates_1518),
   .I0(gates_1332),
   .I1(gates_1331),
   .I2(gates_1330),
   .I3(gates_1329),
   .I4(gates_1328),
   .I5(gates_1327)
);
LUT6 #(
   .INIT(64'b1111111011101000111010001000000011101000100000001000000000000000)  
) LUT6_1519 (
   .O(gates_1519),
   .I0(gates_1338),
   .I1(gates_1337),
   .I2(gates_1336),
   .I3(gates_1335),
   .I4(gates_1334),
   .I5(gates_1333)
);
LUT6 #(
   .INIT(64'b1111111011101000111011001100100011001110100000001000000000000000)  
) LUT6_1520 (
   .O(gates_1520),
   .I0(gates_1344),
   .I1(gates_1343),
   .I2(gates_1342),
   .I3(gates_1341),
   .I4(gates_1340),
   .I5(gates_1339)
);
LUT6 #(
   .INIT(64'b1111111010101000101010001010100011101010100010001000100010000000)  
) LUT6_1521 (
   .O(gates_1521),
   .I0(gates_1350),
   .I1(gates_1349),
   .I2(gates_1348),
   .I3(gates_1347),
   .I4(gates_1346),
   .I5(gates_1345)
);
LUT6 #(
   .INIT(64'b1111111010001000111010001000000011101010000000001000000000000000)  
) LUT6_1522 (
   .O(gates_1522),
   .I0(gates_1356),
   .I1(gates_1355),
   .I2(gates_1354),
   .I3(gates_1353),
   .I4(gates_1352),
   .I5(gates_1351)
);
LUT6 #(
   .INIT(64'b1111110011111100111111001010000011101100110000001100100000000000)  
) LUT6_1523 (
   .O(gates_1523),
   .I0(gates_1362),
   .I1(gates_1361),
   .I2(gates_1360),
   .I3(gates_1359),
   .I4(gates_1358),
   .I5(gates_1357)
);
LUT6 #(
   .INIT(64'b1111111011101000111111101110000010100000100000001000000010000000)  
) LUT6_1524 (
   .O(gates_1524),
   .I0(gates_1368),
   .I1(gates_1367),
   .I2(gates_1366),
   .I3(gates_1365),
   .I4(gates_1364),
   .I5(gates_1363)
);
LUT6 #(
   .INIT(64'b1110111011101000101010001010000011101000101010001000000010000000)  
) LUT6_1525 (
   .O(gates_1525),
   .I0(gates_1374),
   .I1(gates_1373),
   .I2(gates_1372),
   .I3(gates_1371),
   .I4(gates_1370),
   .I5(gates_1369)
);
LUT6 #(
   .INIT(64'b1111111011101000111110000000000011111000111000001000000000000000)  
) LUT6_1526 (
   .O(gates_1526),
   .I0(gates_1380),
   .I1(gates_1379),
   .I2(gates_1378),
   .I3(gates_1377),
   .I4(gates_1376),
   .I5(gates_1375)
);
LUT6 #(
   .INIT(64'b1111111111101000111110001000000011111100100000001111100000000000)  
) LUT6_1527 (
   .O(gates_1527),
   .I0(gates_1386),
   .I1(gates_1385),
   .I2(gates_1384),
   .I3(gates_1383),
   .I4(gates_1382),
   .I5(gates_1381)
);
LUT6 #(
   .INIT(64'b1111111011111000111111101000000011101110100010001110000000000000)  
) LUT6_1528 (
   .O(gates_1528),
   .I0(gates_1392),
   .I1(gates_1391),
   .I2(gates_1390),
   .I3(gates_1389),
   .I4(gates_1388),
   .I5(gates_1387)
);
LUT6 #(
   .INIT(64'b1111111011101100111010001000000011101110110010001100000000000000)  
) LUT6_1529 (
   .O(gates_1529),
   .I0(gates_1398),
   .I1(gates_1397),
   .I2(gates_1396),
   .I3(gates_1395),
   .I4(gates_1394),
   .I5(gates_1393)
);
LUT6 #(
   .INIT(64'b1111111111111110111011101000000011111100101010001010000000000000)  
) LUT6_1530 (
   .O(gates_1530),
   .I0(gates_1404),
   .I1(gates_1403),
   .I2(gates_1402),
   .I3(gates_1401),
   .I4(gates_1400),
   .I5(gates_1399)
);
LUT6 #(
   .INIT(64'b1111111111101010111010101010000011111000101000001010000010000000)  
) LUT6_1531 (
   .O(gates_1531),
   .I0(gates_1410),
   .I1(gates_1409),
   .I2(gates_1408),
   .I3(gates_1407),
   .I4(gates_1406),
   .I5(gates_1405)
);
LUT6 #(
   .INIT(64'b1111111011101000111011001000000011111100100010001100100000000000)  
) LUT6_1532 (
   .O(gates_1532),
   .I0(gates_1416),
   .I1(gates_1415),
   .I2(gates_1414),
   .I3(gates_1413),
   .I4(gates_1412),
   .I5(gates_1411)
);
LUT6 #(
   .INIT(64'b1111111011101000111011001000100010111000100000001000100010000000)  
) LUT6_1533 (
   .O(gates_1533),
   .I0(gates_1422),
   .I1(gates_1421),
   .I2(gates_1420),
   .I3(gates_1419),
   .I4(gates_1418),
   .I5(gates_1417)
);
LUT6 #(
   .INIT(64'b1111111111111000111111001110000011111100101000001110100010000000)  
) LUT6_1534 (
   .O(gates_1534),
   .I0(gates_1428),
   .I1(gates_1427),
   .I2(gates_1426),
   .I3(gates_1425),
   .I4(gates_1424),
   .I5(gates_1423)
);
LUT6 #(
   .INIT(64'b1111111011110100111010001110000011111110110000001100010000000000)  
) LUT6_1535 (
   .O(gates_1535),
   .I0(gates_1434),
   .I1(gates_1433),
   .I2(gates_1432),
   .I3(gates_1431),
   .I4(gates_1430),
   .I5(gates_1429)
);
LUT6 #(
   .INIT(64'b1111100010100000111010000000000010100000000000001000100000000000)  
) LUT6_1536 (
   .O(gates_1536),
   .I0(gates_1440),
   .I1(gates_1439),
   .I2(gates_1438),
   .I3(gates_1437),
   .I4(gates_1436),
   .I5(gates_1435)
);
LUT6 #(
   .INIT(64'b1111111111111110111110101010000011111010111100001010000010000000)  
) LUT6_1537 (
   .O(gates_1537),
   .I0(gates_1446),
   .I1(gates_1445),
   .I2(gates_1444),
   .I3(gates_1443),
   .I4(gates_1442),
   .I5(gates_1441)
);
LUT6 #(
   .INIT(64'b1111110011101000101010001000000011101000100010001000000010000000)  
) LUT6_1538 (
   .O(gates_1538),
   .I0(gates_1452),
   .I1(gates_1451),
   .I2(gates_1450),
   .I3(gates_1449),
   .I4(gates_1448),
   .I5(gates_1447)
);
LUT6 #(
   .INIT(64'b1111111011101100111010001000000011111100100000001000000000000000)  
) LUT6_1539 (
   .O(gates_1539),
   .I0(gates_1458),
   .I1(gates_1457),
   .I2(gates_1456),
   .I3(gates_1455),
   .I4(gates_1454),
   .I5(gates_1453)
);
LUT6 #(
   .INIT(64'b1111111111101100111011001100000011111110100000001110000000000000)  
) LUT6_1540 (
   .O(gates_1540),
   .I0(gates_1464),
   .I1(gates_1463),
   .I2(gates_1462),
   .I3(gates_1461),
   .I4(gates_1460),
   .I5(gates_1459)
);
LUT6 #(
   .INIT(64'b1111111111101110111010001000100011101000100000001000000010000000)  
) LUT6_1541 (
   .O(gates_1541),
   .I0(gates_1470),
   .I1(gates_1469),
   .I2(gates_1468),
   .I3(gates_1467),
   .I4(gates_1466),
   .I5(gates_1465)
);
LUT6 #(
   .INIT(64'b1111111011101000110010001010000011101000100000001000000000000000)  
) LUT6_1542 (
   .O(gates_1542),
   .I0(gates_1476),
   .I1(gates_1475),
   .I2(gates_1474),
   .I3(gates_1473),
   .I4(gates_1472),
   .I5(gates_1471)
);
LUT6 #(
   .INIT(64'b1111111111101000111111001110000011101100100000001100100000000000)  
) LUT6_1543 (
   .O(gates_1543),
   .I0(gates_1482),
   .I1(gates_1481),
   .I2(gates_1480),
   .I3(gates_1479),
   .I4(gates_1478),
   .I5(gates_1477)
);
LUT6 #(
   .INIT(64'b1111111111111110111111000100000011111010110010001100000000000000)  
) LUT6_1544 (
   .O(gates_1544),
   .I0(gates_1488),
   .I1(gates_1487),
   .I2(gates_1486),
   .I3(gates_1485),
   .I4(gates_1484),
   .I5(gates_1483)
);
LUT6 #(
   .INIT(64'b1111111111111100111011101000100011101100100010001000000000000000)  
) LUT6_1545 (
   .O(gates_1545),
   .I0(gates_1494),
   .I1(gates_1493),
   .I2(gates_1492),
   .I3(gates_1491),
   .I4(gates_1490),
   .I5(gates_1489)
);
LUT6 #(
   .INIT(64'b1111111011101000111010001100100011111010100010001100000010000000)  
) LUT6_1546 (
   .O(gates_1546),
   .I0(gates_1500),
   .I1(gates_1499),
   .I2(gates_1498),
   .I3(gates_1497),
   .I4(gates_1496),
   .I5(gates_1495)
);
LUT6 #(
   .INIT(64'b1111111011111000111110001110100011101110111010001110100010101000)  
) LUT6_1547 (
   .O(gates_1547),
   .I0(gates_1506),
   .I1(gates_1505),
   .I2(gates_1504),
   .I3(gates_1503),
   .I4(gates_1502),
   .I5(gates_1501)
);
LUT6 #(
   .INIT(64'b1111111111101100111011101100000011101000100000001000100010000000)  
) LUT6_1548 (
   .O(gates_1548),
   .I0(gates_1512),
   .I1(gates_1511),
   .I2(gates_1510),
   .I3(gates_1509),
   .I4(gates_1508),
   .I5(gates_1507)
);
LUT6 #(
   .INIT(64'b1111111011100010111011001000000011111100101010001100110000000000)  
) LUT6_1549 (
   .O(gates_1549),
   .I0(gates_1518),
   .I1(gates_1517),
   .I2(gates_1516),
   .I3(gates_1515),
   .I4(gates_1514),
   .I5(gates_1513)
);
LUT6 #(
   .INIT(64'b1111111011101000111110101101100011111000000000001110000000000000)  
) LUT6_1550 (
   .O(gates_1550),
   .I0(gates_1524),
   .I1(gates_1523),
   .I2(gates_1522),
   .I3(gates_1521),
   .I4(gates_1520),
   .I5(gates_1519)
);
LUT6 #(
   .INIT(64'b1111111111111010111110110010100011101110110001000010000000000000)  
) LUT6_1551 (
   .O(gates_1551),
   .I0(gates_1530),
   .I1(gates_1529),
   .I2(gates_1528),
   .I3(gates_1527),
   .I4(gates_1526),
   .I5(gates_1525)
);
LUT6 #(
   .INIT(64'b1111111011111000111110101100000011101000111010101100000000000000)  
) LUT6_1552 (
   .O(gates_1552),
   .I0(gates_1536),
   .I1(gates_1535),
   .I2(gates_1534),
   .I3(gates_1533),
   .I4(gates_1532),
   .I5(gates_1531)
);
LUT6 #(
   .INIT(64'b1111111011111100111110001110100011111110110000001000100000000000)  
) LUT6_1553 (
   .O(gates_1553),
   .I0(gates_1542),
   .I1(gates_1541),
   .I2(gates_1540),
   .I3(gates_1539),
   .I4(gates_1538),
   .I5(gates_1537)
);
LUT6 #(
   .INIT(64'b1111111110101010111010011000100010111000111000001000100010000000)  
) LUT6_1554 (
   .O(gates_1554),
   .I0(gates_1548),
   .I1(gates_1547),
   .I2(gates_1546),
   .I3(gates_1545),
   .I4(gates_1544),
   .I5(gates_1543)
);
LUT6 #(
   .INIT(64'b1110111011110000111110001000000011111110101100001110001010000000)  
) LUT6_1555 (
   .O(gates_1555),
   .I0(gates_1554),
   .I1(gates_1553),
   .I2(gates_1552),
   .I3(gates_1551),
   .I4(gates_1550),
   .I5(gates_1549)
);



endmodule