module lut_5level_tree5(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [576:0] data_in,
                       input       data_valid,
                       output      data_out     
                       );
wire    [576:0] InputBits;
wire    gates_1, gates_2, gates_3, gates_4, gates_5, gates_6, gates_7, gates_8, gates_9, gates_10, gates_11, gates_12, gates_13, gates_14, gates_15, gates_16, gates_17, gates_18, gates_19, gates_20, gates_21, gates_22, gates_23, gates_24, gates_25, gates_26, gates_27, gates_28, gates_29, gates_30, gates_31, gates_32, gates_33, gates_34, gates_35, gates_36, gates_37, gates_38, gates_39, gates_40, gates_41, gates_42, gates_43, gates_44, gates_45, gates_46, gates_47, gates_48, gates_49, gates_50, gates_51, gates_52, gates_53, gates_54, gates_55, gates_56, gates_57, gates_58, gates_59, gates_60, gates_61, gates_62, gates_63, gates_64, gates_65, gates_66, gates_67, gates_68, gates_69, gates_70, gates_71, gates_72, gates_73, gates_74, gates_75, gates_76, gates_77, gates_78, gates_79, gates_80, gates_81, gates_82, gates_83, gates_84, gates_85, gates_86, gates_87, gates_88, gates_89, gates_90, gates_91, gates_92, gates_93, gates_94, gates_95, gates_96, gates_97, gates_98, gates_99, gates_100, gates_101, gates_102, gates_103, gates_104, gates_105, gates_106, gates_107, gates_108, gates_109, gates_110, gates_111, gates_112, gates_113, gates_114, gates_115, gates_116, gates_117, gates_118, gates_119, gates_120, gates_121, gates_122, gates_123, gates_124, gates_125, gates_126, gates_127, gates_128, gates_129, gates_130, gates_131, gates_132, gates_133, gates_134, gates_135, gates_136, gates_137, gates_138, gates_139, gates_140, gates_141, gates_142, gates_143, gates_144, gates_145, gates_146, gates_147, gates_148, gates_149, gates_150, gates_151, gates_152, gates_153, gates_154, gates_155, gates_156, gates_157, gates_158, gates_159, gates_160, gates_161, gates_162, gates_163, gates_164, gates_165, gates_166, gates_167, gates_168, gates_169, gates_170, gates_171, gates_172, gates_173, gates_174, gates_175, gates_176, gates_177, gates_178, gates_179, gates_180, gates_181, gates_182, gates_183, gates_184, gates_185, gates_186, gates_187, gates_188, gates_189, gates_190, gates_191, gates_192, gates_193, gates_194, gates_195, gates_196, gates_197, gates_198, gates_199, gates_200, gates_201, gates_202, gates_203, gates_204, gates_205, gates_206, gates_207, gates_208, gates_209, gates_210, gates_211, gates_212, gates_213, gates_214, gates_215, gates_216, gates_217, gates_218, gates_219, gates_220, gates_221, gates_222, gates_223, gates_224, gates_225, gates_226, gates_227, gates_228, gates_229, gates_230, gates_231, gates_232, gates_233, gates_234, gates_235, gates_236, gates_237, gates_238, gates_239, gates_240, gates_241, gates_242, gates_243, gates_244, gates_245, gates_246, gates_247, gates_248, gates_249, gates_250, gates_251, gates_252, gates_253, gates_254, gates_255, gates_256, gates_257, gates_258, gates_259, gates_260, gates_261, gates_262, gates_263, gates_264, gates_265, gates_266, gates_267, gates_268, gates_269, gates_270, gates_271, gates_272, gates_273, gates_274, gates_275, gates_276, gates_277, gates_278, gates_279, gates_280, gates_281, gates_282, gates_283, gates_284, gates_285, gates_286, gates_287, gates_288, gates_289, gates_290, gates_291, gates_292, gates_293, gates_294, gates_295, gates_296, gates_297, gates_298, gates_299, gates_300, gates_301, gates_302, gates_303, gates_304, gates_305, gates_306, gates_307, gates_308, gates_309, gates_310, gates_311, gates_312, gates_313, gates_314, gates_315, gates_316, gates_317, gates_318, gates_319, gates_320, gates_321, gates_322, gates_323, gates_324, gates_325, gates_326, gates_327, gates_328, gates_329, gates_330, gates_331, gates_332, gates_333, gates_334, gates_335, gates_336, gates_337, gates_338, gates_339, gates_340, gates_341, gates_342, gates_343, gates_344, gates_345, gates_346, gates_347, gates_348, gates_349, gates_350, gates_351, gates_352, gates_353, gates_354, gates_355, gates_356, gates_357, gates_358, gates_359, gates_360, gates_361, gates_362, gates_363, gates_364, gates_365, gates_366, gates_367, gates_368, gates_369, gates_370, gates_371, gates_372, gates_373, gates_374, gates_375, gates_376, gates_377, gates_378, gates_379, gates_380, gates_381, gates_382, gates_383, gates_384, gates_385, gates_386, gates_387, gates_388, gates_389, gates_390, gates_391, gates_392, gates_393, gates_394, gates_395, gates_396, gates_397, gates_398, gates_399, gates_400, gates_401, gates_402, gates_403, gates_404, gates_405, gates_406, gates_407, gates_408, gates_409, gates_410, gates_411, gates_412, gates_413, gates_414, gates_415, gates_416, gates_417, gates_418, gates_419, gates_420, gates_421, gates_422, gates_423, gates_424, gates_425, gates_426, gates_427, gates_428, gates_429, gates_430, gates_431, gates_432, gates_433, gates_434, gates_435, gates_436, gates_437, gates_438, gates_439, gates_440, gates_441, gates_442, gates_443, gates_444, gates_445, gates_446, gates_447, gates_448, gates_449, gates_450, gates_451, gates_452, gates_453, gates_454, gates_455, gates_456, gates_457, gates_458, gates_459, gates_460, gates_461, gates_462, gates_463, gates_464, gates_465, gates_466, gates_467, gates_468, gates_469, gates_470, gates_471, gates_472, gates_473, gates_474, gates_475, gates_476, gates_477, gates_478, gates_479, gates_480, gates_481, gates_482, gates_483, gates_484, gates_485, gates_486, gates_487, gates_488, gates_489, gates_490, gates_491, gates_492, gates_493, gates_494, gates_495, gates_496, gates_497, gates_498, gates_499, gates_500, gates_501, gates_502, gates_503, gates_504, gates_505, gates_506, gates_507, gates_508, gates_509, gates_510, gates_511, gates_512, gates_513, gates_514, gates_515, gates_516, gates_517, gates_518, gates_519, gates_520, gates_521, gates_522, gates_523, gates_524, gates_525, gates_526, gates_527, gates_528, gates_529, gates_530, gates_531, gates_532, gates_533, gates_534, gates_535, gates_536, gates_537, gates_538, gates_539, gates_540, gates_541, gates_542, gates_543, gates_544, gates_545, gates_546, gates_547, gates_548, gates_549, gates_550, gates_551, gates_552, gates_553, gates_554, gates_555, gates_556, gates_557, gates_558, gates_559, gates_560, gates_561, gates_562, gates_563, gates_564, gates_565, gates_566, gates_567, gates_568, gates_569, gates_570, gates_571, gates_572, gates_573, gates_574, gates_575, gates_576, gates_577, gates_578, gates_579, gates_580, gates_581, gates_582, gates_583, gates_584, gates_585, gates_586, gates_587, gates_588, gates_589, gates_590, gates_591, gates_592, gates_593, gates_594, gates_595, gates_596, gates_597, gates_598, gates_599, gates_600, gates_601, gates_602, gates_603, gates_604, gates_605, gates_606, gates_607, gates_608, gates_609, gates_610, gates_611, gates_612, gates_613, gates_614, gates_615, gates_616, gates_617, gates_618, gates_619, gates_620, gates_621, gates_622, gates_623, gates_624, gates_625, gates_626, gates_627, gates_628, gates_629, gates_630, gates_631, gates_632, gates_633, gates_634, gates_635, gates_636, gates_637, gates_638, gates_639, gates_640, gates_641, gates_642, gates_643, gates_644, gates_645, gates_646, gates_647, gates_648, gates_649, gates_650, gates_651, gates_652, gates_653, gates_654, gates_655, gates_656, gates_657, gates_658, gates_659, gates_660, gates_661, gates_662, gates_663, gates_664, gates_665, gates_666, gates_667, gates_668, gates_669, gates_670, gates_671, gates_672, gates_673, gates_674, gates_675, gates_676, gates_677, gates_678, gates_679, gates_680, gates_681, gates_682, gates_683, gates_684, gates_685, gates_686, gates_687, gates_688, gates_689, gates_690, gates_691, gates_692, gates_693, gates_694, gates_695, gates_696, gates_697, gates_698, gates_699, gates_700, gates_701, gates_702, gates_703, gates_704, gates_705, gates_706, gates_707, gates_708, gates_709, gates_710, gates_711, gates_712, gates_713, gates_714, gates_715, gates_716, gates_717, gates_718, gates_719, gates_720, gates_721, gates_722, gates_723, gates_724, gates_725, gates_726, gates_727, gates_728, gates_729, gates_730, gates_731, gates_732, gates_733, gates_734, gates_735, gates_736, gates_737, gates_738, gates_739, gates_740, gates_741, gates_742, gates_743, gates_744, gates_745, gates_746, gates_747, gates_748, gates_749, gates_750, gates_751, gates_752, gates_753, gates_754, gates_755, gates_756, gates_757, gates_758, gates_759, gates_760, gates_761, gates_762, gates_763, gates_764, gates_765, gates_766, gates_767, gates_768, gates_769, gates_770, gates_771, gates_772, gates_773, gates_774, gates_775, gates_776, gates_777, gates_778, gates_779, gates_780, gates_781, gates_782, gates_783, gates_784, gates_785, gates_786, gates_787, gates_788, gates_789, gates_790, gates_791, gates_792, gates_793, gates_794, gates_795, gates_796, gates_797, gates_798, gates_799, gates_800, gates_801, gates_802, gates_803, gates_804, gates_805, gates_806, gates_807, gates_808, gates_809, gates_810, gates_811, gates_812, gates_813, gates_814, gates_815, gates_816, gates_817, gates_818, gates_819, gates_820, gates_821, gates_822, gates_823, gates_824, gates_825, gates_826, gates_827, gates_828, gates_829, gates_830, gates_831, gates_832, gates_833, gates_834, gates_835, gates_836, gates_837, gates_838, gates_839, gates_840, gates_841, gates_842, gates_843, gates_844, gates_845, gates_846, gates_847, gates_848, gates_849, gates_850, gates_851, gates_852, gates_853, gates_854, gates_855, gates_856, gates_857, gates_858, gates_859, gates_860, gates_861, gates_862, gates_863, gates_864, gates_865, gates_866, gates_867, gates_868, gates_869, gates_870, gates_871, gates_872, gates_873, gates_874, gates_875, gates_876, gates_877, gates_878, gates_879, gates_880, gates_881, gates_882, gates_883, gates_884, gates_885, gates_886, gates_887, gates_888, gates_889, gates_890, gates_891, gates_892, gates_893, gates_894, gates_895, gates_896, gates_897, gates_898, gates_899, gates_900, gates_901, gates_902, gates_903, gates_904, gates_905, gates_906, gates_907, gates_908, gates_909, gates_910, gates_911, gates_912, gates_913, gates_914, gates_915, gates_916, gates_917, gates_918, gates_919, gates_920, gates_921, gates_922, gates_923, gates_924, gates_925, gates_926, gates_927, gates_928, gates_929, gates_930, gates_931, gates_932, gates_933, gates_934, gates_935, gates_936, gates_937, gates_938, gates_939, gates_940, gates_941, gates_942, gates_943, gates_944, gates_945, gates_946, gates_947, gates_948, gates_949, gates_950, gates_951, gates_952, gates_953, gates_954, gates_955, gates_956, gates_957, gates_958, gates_959, gates_960, gates_961, gates_962, gates_963, gates_964, gates_965, gates_966, gates_967, gates_968, gates_969, gates_970, gates_971, gates_972, gates_973, gates_974, gates_975, gates_976, gates_977, gates_978, gates_979, gates_980, gates_981, gates_982, gates_983, gates_984, gates_985, gates_986, gates_987, gates_988, gates_989, gates_990, gates_991, gates_992, gates_993, gates_994, gates_995, gates_996, gates_997, gates_998, gates_999, gates_1000, gates_1001, gates_1002, gates_1003, gates_1004, gates_1005, gates_1006, gates_1007, gates_1008, gates_1009, gates_1010, gates_1011, gates_1012, gates_1013, gates_1014, gates_1015, gates_1016, gates_1017, gates_1018, gates_1019, gates_1020, gates_1021, gates_1022, gates_1023, gates_1024, gates_1025, gates_1026, gates_1027, gates_1028, gates_1029, gates_1030, gates_1031, gates_1032, gates_1033, gates_1034, gates_1035, gates_1036, gates_1037, gates_1038, gates_1039, gates_1040, gates_1041, gates_1042, gates_1043, gates_1044, gates_1045, gates_1046, gates_1047, gates_1048, gates_1049, gates_1050, gates_1051, gates_1052, gates_1053, gates_1054, gates_1055, gates_1056, gates_1057, gates_1058, gates_1059, gates_1060, gates_1061, gates_1062, gates_1063, gates_1064, gates_1065, gates_1066, gates_1067, gates_1068, gates_1069, gates_1070, gates_1071, gates_1072, gates_1073, gates_1074, gates_1075, gates_1076, gates_1077, gates_1078, gates_1079, gates_1080, gates_1081, gates_1082, gates_1083, gates_1084, gates_1085, gates_1086, gates_1087, gates_1088, gates_1089, gates_1090, gates_1091, gates_1092, gates_1093, gates_1094, gates_1095, gates_1096, gates_1097, gates_1098, gates_1099, gates_1100, gates_1101, gates_1102, gates_1103, gates_1104, gates_1105, gates_1106, gates_1107, gates_1108, gates_1109, gates_1110, gates_1111, gates_1112, gates_1113, gates_1114, gates_1115, gates_1116, gates_1117, gates_1118, gates_1119, gates_1120, gates_1121, gates_1122, gates_1123, gates_1124, gates_1125, gates_1126, gates_1127, gates_1128, gates_1129, gates_1130, gates_1131, gates_1132, gates_1133, gates_1134, gates_1135, gates_1136, gates_1137, gates_1138, gates_1139, gates_1140, gates_1141, gates_1142, gates_1143, gates_1144, gates_1145, gates_1146, gates_1147, gates_1148, gates_1149, gates_1150, gates_1151, gates_1152, gates_1153, gates_1154, gates_1155, gates_1156, gates_1157, gates_1158, gates_1159, gates_1160, gates_1161, gates_1162, gates_1163, gates_1164, gates_1165, gates_1166, gates_1167, gates_1168, gates_1169, gates_1170, gates_1171, gates_1172, gates_1173, gates_1174, gates_1175, gates_1176, gates_1177, gates_1178, gates_1179, gates_1180, gates_1181, gates_1182, gates_1183, gates_1184, gates_1185, gates_1186, gates_1187, gates_1188, gates_1189, gates_1190, gates_1191, gates_1192, gates_1193, gates_1194, gates_1195, gates_1196, gates_1197, gates_1198, gates_1199, gates_1200, gates_1201, gates_1202, gates_1203, gates_1204, gates_1205, gates_1206, gates_1207, gates_1208, gates_1209, gates_1210, gates_1211, gates_1212, gates_1213, gates_1214, gates_1215, gates_1216, gates_1217, gates_1218, gates_1219, gates_1220, gates_1221, gates_1222, gates_1223, gates_1224, gates_1225, gates_1226, gates_1227, gates_1228, gates_1229, gates_1230, gates_1231, gates_1232, gates_1233, gates_1234, gates_1235, gates_1236, gates_1237, gates_1238, gates_1239, gates_1240, gates_1241, gates_1242, gates_1243, gates_1244, gates_1245, gates_1246, gates_1247, gates_1248, gates_1249, gates_1250, gates_1251, gates_1252, gates_1253, gates_1254, gates_1255, gates_1256, gates_1257, gates_1258, gates_1259, gates_1260, gates_1261, gates_1262, gates_1263, gates_1264, gates_1265, gates_1266, gates_1267, gates_1268, gates_1269, gates_1270, gates_1271, gates_1272, gates_1273, gates_1274, gates_1275, gates_1276, gates_1277, gates_1278, gates_1279, gates_1280, gates_1281, gates_1282, gates_1283, gates_1284, gates_1285, gates_1286, gates_1287, gates_1288, gates_1289, gates_1290, gates_1291, gates_1292, gates_1293, gates_1294, gates_1295, gates_1296, gates_1297, gates_1298, gates_1299, gates_1300, gates_1301, gates_1302, gates_1303, gates_1304, gates_1305, gates_1306, gates_1307, gates_1308, gates_1309, gates_1310, gates_1311, gates_1312, gates_1313, gates_1314, gates_1315, gates_1316, gates_1317, gates_1318, gates_1319, gates_1320, gates_1321, gates_1322, gates_1323, gates_1324, gates_1325, gates_1326, gates_1327, gates_1328, gates_1329, gates_1330, gates_1331, gates_1332, gates_1333, gates_1334, gates_1335, gates_1336, gates_1337, gates_1338, gates_1339, gates_1340, gates_1341, gates_1342, gates_1343, gates_1344, gates_1345, gates_1346, gates_1347, gates_1348, gates_1349, gates_1350, gates_1351, gates_1352, gates_1353, gates_1354, gates_1355, gates_1356, gates_1357, gates_1358, gates_1359, gates_1360, gates_1361, gates_1362, gates_1363, gates_1364, gates_1365, gates_1366, gates_1367, gates_1368, gates_1369, gates_1370, gates_1371, gates_1372, gates_1373, gates_1374, gates_1375, gates_1376, gates_1377, gates_1378, gates_1379, gates_1380, gates_1381, gates_1382, gates_1383, gates_1384, gates_1385, gates_1386, gates_1387, gates_1388, gates_1389, gates_1390, gates_1391, gates_1392, gates_1393, gates_1394, gates_1395, gates_1396, gates_1397, gates_1398, gates_1399, gates_1400, gates_1401, gates_1402, gates_1403, gates_1404, gates_1405, gates_1406, gates_1407, gates_1408, gates_1409, gates_1410, gates_1411, gates_1412, gates_1413, gates_1414, gates_1415, gates_1416, gates_1417, gates_1418, gates_1419, gates_1420, gates_1421, gates_1422, gates_1423, gates_1424, gates_1425, gates_1426, gates_1427, gates_1428, gates_1429, gates_1430, gates_1431, gates_1432, gates_1433, gates_1434, gates_1435, gates_1436, gates_1437, gates_1438, gates_1439, gates_1440, gates_1441, gates_1442, gates_1443, gates_1444, gates_1445, gates_1446, gates_1447, gates_1448, gates_1449, gates_1450, gates_1451, gates_1452, gates_1453, gates_1454, gates_1455, gates_1456, gates_1457, gates_1458, gates_1459, gates_1460, gates_1461, gates_1462, gates_1463, gates_1464, gates_1465, gates_1466, gates_1467, gates_1468, gates_1469, gates_1470, gates_1471, gates_1472, gates_1473, gates_1474, gates_1475, gates_1476, gates_1477, gates_1478, gates_1479, gates_1480, gates_1481, gates_1482, gates_1483, gates_1484, gates_1485, gates_1486, gates_1487, gates_1488, gates_1489, gates_1490, gates_1491, gates_1492, gates_1493, gates_1494, gates_1495, gates_1496, gates_1497, gates_1498, gates_1499, gates_1500, gates_1501, gates_1502, gates_1503, gates_1504, gates_1505, gates_1506, gates_1507, gates_1508, gates_1509, gates_1510, gates_1511, gates_1512, gates_1513, gates_1514, gates_1515, gates_1516, gates_1517, gates_1518, gates_1519, gates_1520, gates_1521, gates_1522, gates_1523, gates_1524, gates_1525, gates_1526, gates_1527, gates_1528, gates_1529, gates_1530, gates_1531, gates_1532, gates_1533, gates_1534, gates_1535, gates_1536, gates_1537, gates_1538, gates_1539, gates_1540, gates_1541, gates_1542, gates_1543, gates_1544, gates_1545, gates_1546, gates_1547, gates_1548, gates_1549, gates_1550, gates_1551, gates_1552, gates_1553, gates_1554, gates_1555;

assign  InputBits = data_in;
//assign  data_out = data_valid & gates[807];
assign  data_out = data_valid & gates_408;

LUT6 #(
   .INIT(64'b0110000111010101111101101010101110101011010000111110100111101010)  
) LUT6_1 (
   .O(gates_819),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0010001001001010100000010011011001101011011000011011110000101101)  
) LUT6_2 (
   .O(gates_46),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1011010001100000011101011001011011011111101100001001100010110100)  
) LUT6_3 (
   .O(gates_1179),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1110011101011100110001111111011100110001011011000100110010011110)  
) LUT6_4 (
   .O(gates_1528),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0100111110111100011111101001010000010000000001100000010111000001)  
) LUT6_5 (
   .O(gates_307),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0110111110000011111001111010001000010010100110000001001010001111)  
) LUT6_6 (
   .O(gates_297),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1001000111110001110100101111010000100110110110000010111010110001)  
) LUT6_7 (
   .O(gates_1517),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0001101110001101000101000110000010001110101101111100111101011110)  
) LUT6_8 (
   .O(gates_907),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0100111110111110100101100001011000110011010110000111011000011101)  
) LUT6_9 (
   .O(gates_106),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1010001011010100101000110100100110000111101010001000111110101100)  
) LUT6_10 (
   .O(gates_948),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1011100010001010101101110100010100001101001010110111111000100101)  
) LUT6_11 (
   .O(gates_1144),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0110011110111110011010010010101000001001101010110100011101011010)  
) LUT6_12 (
   .O(gates_619),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1111010110000100001100000000010010110000001001110001010010011100)  
) LUT6_13 (
   .O(gates_1414),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0111011010010011000000011110111111000110011100000110011111101110)  
) LUT6_14 (
   .O(gates_801),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1100111010001001001110100000001110010101101100000010111111000111)  
) LUT6_15 (
   .O(gates_1378),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0011111001100100010000001111110011001111101111000010010011110011)  
) LUT6_16 (
   .O(gates_1397),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b1000100011101011000001010101110001001111010111110111000000010110)  
) LUT6_17 (
   .O(gates_1415),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1101101111101101001100000101011100001101001111001101100111000001)  
) LUT6_18 (
   .O(gates_1470),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0001010111101100011111000000011000111100000011110001000100001010)  
) LUT6_19 (
   .O(gates_740),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0110011100001011000010011000001111000011011000111111111000101000)  
) LUT6_20 (
   .O(gates_1463),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0000001101111001000100011001011111100001100111110010100110010110)  
) LUT6_21 (
   .O(gates_1530),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0101110000001111100111001010010010100110110101011111001110010011)  
) LUT6_22 (
   .O(gates_341),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0100110010100100101011001101111010111000110101000011001011011000)  
) LUT6_23 (
   .O(gates_1367),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0001110101100101110011001101111101001111110101000110001011011101)  
) LUT6_24 (
   .O(gates_1428),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1101010101001110101101011001100111110000010011110110100101001100)  
) LUT6_25 (
   .O(gates_1408),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0011001000111011110100010101101011010000110110101001111001001001)  
) LUT6_26 (
   .O(gates_998),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1001100011111101100110110011100100111100100001101111110100110000)  
) LUT6_27 (
   .O(gates_1240),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1000010000001001001001111101110110111001001000100101011100100110)  
) LUT6_28 (
   .O(gates_577),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1000000000011100101000100000110100100001111101111101011010101010)  
) LUT6_29 (
   .O(gates_960),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1010111000100111111110111101001100001010001010010101101011101101)  
) LUT6_30 (
   .O(gates_318),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1111000000111010001100011110011101110101001001100100111010110111)  
) LUT6_31 (
   .O(gates_449),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0011000000101000100111000101011111011101100111001011001010110100)  
) LUT6_32 (
   .O(gates_830),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0100011110000111101100110010000010100101101101010100100111010100)  
) LUT6_33 (
   .O(gates_1088),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1110010000110011100111011111001110100000011011111010100010011101)  
) LUT6_34 (
   .O(gates_1262),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0111000111011010111101011111011010101010101101000100000010011010)  
) LUT6_35 (
   .O(gates_327),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0101110000111010001010111111110101110011001010110110010101010001)  
) LUT6_36 (
   .O(gates_964),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1000001101001101010111100011111101010101001000000111001000100101)  
) LUT6_37 (
   .O(gates_1009),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0001111110001111110101111110101001011101110100011110100000101001)  
) LUT6_38 (
   .O(gates_97),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0101011100100011101110101110011001100111111000001001111100101000)  
) LUT6_39 (
   .O(gates_1555),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1000000010111101000111010011011001110011111001111001010101101110)  
) LUT6_40 (
   .O(gates_175),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0011001111101100111011011110011010011111100110011011000100100000)  
) LUT6_41 (
   .O(gates_202),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0000011101000101010011110000010111001000100001110101111000011111)  
) LUT6_42 (
   .O(gates_188),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0110000110001100100010001111111001100111110010111010110100111000)  
) LUT6_43 (
   .O(gates_293),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1010101100101100000110011001111001000111101010111111001100001001)  
) LUT6_44 (
   .O(gates_1315),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0010001110010000011011111000100111001111111010010101111110111011)  
) LUT6_45 (
   .O(gates_1329),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0000000111000111110001010000001011001110010111100011111011111100)  
) LUT6_46 (
   .O(gates_1098),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1110101110110101110011101101110001110101001110100111000001001000)  
) LUT6_47 (
   .O(gates_868),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0001101110000111100011010111101110110001001011111100000001011110)  
) LUT6_48 (
   .O(gates_250),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1001011110011100001001101100111010110000101111110011011100001101)  
) LUT6_49 (
   .O(gates_378),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1011110101100001101110000111010010010111100100100001110100000110)  
) LUT6_50 (
   .O(gates_1137),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0000100111101111110000101000010000101000011000000101010010100000)  
) LUT6_51 (
   .O(gates_539),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0010111111111110101111110011101111011000010110001100111100110101)  
) LUT6_52 (
   .O(gates_1418),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1111111011100101011100110011100110100101011000110111110100011010)  
) LUT6_53 (
   .O(gates_817),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1001110000000100110010010110001101101000101000110000110000010010)  
) LUT6_54 (
   .O(gates_970),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0011110011111111011000001101111100100010011010101001100010001101)  
) LUT6_55 (
   .O(gates_637),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0110011111010110100001001010101011011100110100000011011101000010)  
) LUT6_56 (
   .O(gates_947),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1101000010111000101011111111111100000101110110101110011110010100)  
) LUT6_57 (
   .O(gates_683),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0110001011001111010010011100000010011100011011001100011100001110)  
) LUT6_58 (
   .O(gates_1343),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1101110101011000000100000100001000010000100111110110101100010001)  
) LUT6_59 (
   .O(gates_1152),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1101100010101110100011001111101001000101010110000111001001011000)  
) LUT6_60 (
   .O(gates_747),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0000110100100111100010011100000001011011011111001110000100000101)  
) LUT6_61 (
   .O(gates_275),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1100100101010011011011011111101111000100000101101000100010101100)  
) LUT6_62 (
   .O(gates_1177),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1110101100100011100000010000101101010001001000101010001101010111)  
) LUT6_63 (
   .O(gates_411),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0110110000010101000000001011001000111000000010010101001101110101)  
) LUT6_64 (
   .O(gates_1122),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0010101011011101101010101001011110101010101011101111010101001101)  
) LUT6_65 (
   .O(gates_1158),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1100010110010011110000010100101011111101010100110111010100001110)  
) LUT6_66 (
   .O(gates_1545),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1010100011011000100100010101001100111100100110011010001111111101)  
) LUT6_67 (
   .O(gates_460),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1111100011111001000101100101001010101000010010101101010000110010)  
) LUT6_68 (
   .O(gates_1146),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1100110110010000000010100101000100011011100111111001111101000101)  
) LUT6_69 (
   .O(gates_593),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0010011110101000110101000111011011010100111110010000010011100110)  
) LUT6_70 (
   .O(gates_7),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1001010111110011000001111100001111010010010001101011010010011011)  
) LUT6_71 (
   .O(gates_911),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0100101110001010010101010000111010011101111100110111101100100101)  
) LUT6_72 (
   .O(gates_980),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1011110001010001110111011011000100100001000001011010010100010010)  
) LUT6_73 (
   .O(gates_315),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1110010010110111011000101010001011001000111110111011101011110000)  
) LUT6_74 (
   .O(gates_1033),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1001010000001101011001111001110011000111010000000010110100000101)  
) LUT6_75 (
   .O(gates_548),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1001110111101110110001100101111001111111000000100111101110011101)  
) LUT6_76 (
   .O(gates_1149),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b0100100110000110000001100110001000111110111001001100100101110100)  
) LUT6_77 (
   .O(gates_549),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0000101101011010010100000001100010000000010100011100010101010111)  
) LUT6_78 (
   .O(gates_312),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0101100010101000100111010010111110000110010101101101010000000000)  
) LUT6_79 (
   .O(gates_771),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0100011101101111001100000000010101011001101010001110111101110010)  
) LUT6_80 (
   .O(gates_617),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0001010010101100101011110111000110111011001010100000101101001100)  
) LUT6_81 (
   .O(gates_1446),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1010010101111001111001101011111010010101101101110110111101110011)  
) LUT6_82 (
   .O(gates_601),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1010001111000100111000100101001011100001010111110001111001100011)  
) LUT6_83 (
   .O(gates_1365),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0011010001111110110100100011010000010110101010000101000111100011)  
) LUT6_84 (
   .O(gates_977),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0111110110001110110101000001010010111001100011000011110110000111)  
) LUT6_85 (
   .O(gates_64),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0001010111000100001110110100010111101101010011010111100100110101)  
) LUT6_86 (
   .O(gates_459),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1111001100100001100111111101100111011011101100000101111011111110)  
) LUT6_87 (
   .O(gates_141),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1101100011010000011010011101111010110111010101000101111110100011)  
) LUT6_88 (
   .O(gates_655),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1101111100011100010011001110101000010111111011111011111001110010)  
) LUT6_89 (
   .O(gates_30),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1011100101011000011001001110000001011010001101100100000110100111)  
) LUT6_90 (
   .O(gates_1290),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b1111011100011100100101111001011111111011000011101101101111000001)  
) LUT6_91 (
   .O(gates_1362),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0100011011111011000100100010100110000111101000011111010100001010)  
) LUT6_92 (
   .O(gates_8),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0111101101101000000000101000111010100100100111110101101111110011)  
) LUT6_93 (
   .O(gates_353),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1001101110011010110111000101101001010110101001001101111001100111)  
) LUT6_94 (
   .O(gates_4),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1111011001100010010100011111111111011000000111000001011100100001)  
) LUT6_95 (
   .O(gates_57),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0000101001111000111011011001111110110110100001101111010000110100)  
) LUT6_96 (
   .O(gates_452),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1101010001111001001001000011101110001110011011111000011010000010)  
) LUT6_97 (
   .O(gates_1001),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1100000101111110101101100010011000111111010011001110101010010011)  
) LUT6_98 (
   .O(gates_301),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1010111100100111101110100101111110111000100010101111100111111100)  
) LUT6_99 (
   .O(gates_567),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0100000100110100011111001000111110111101100000100111111010001110)  
) LUT6_100 (
   .O(gates_1167),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0101101101000100101110001111011110000010111001000111110000011000)  
) LUT6_101 (
   .O(gates_1082),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1001001110111001010011101101000100000111001001100101010000011110)  
) LUT6_102 (
   .O(gates_406),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0110000110100100101010101010110001000111011001100100110101010100)  
) LUT6_103 (
   .O(gates_641),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0000001110000101100011001110100110110010110100000101010000100000)  
) LUT6_104 (
   .O(gates_1204),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0001111101000010001001111010000001111001110010001001110100011001)  
) LUT6_105 (
   .O(gates_1048),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1001111100000111000001001100010001011001101111111111001111001101)  
) LUT6_106 (
   .O(gates_335),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0011111111100010100100011100011001111011101101001101000000111011)  
) LUT6_107 (
   .O(gates_1221),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b1011011101000110011000100100011100101111110000110000110100110011)  
) LUT6_108 (
   .O(gates_381),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0010011110101111100010110011111010010001010111110001110001111000)  
) LUT6_109 (
   .O(gates_935),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0111111010011110000111001110101001011001010110110000111101000111)  
) LUT6_110 (
   .O(gates_159),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1111010001111110100000011101010000001101110010100000011110101001)  
) LUT6_111 (
   .O(gates_69),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0011110010110100000011000111111010110001100111101010010100011110)  
) LUT6_112 (
   .O(gates_1010),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b1100101111001010010101111000001011110010000001101100011010000100)  
) LUT6_113 (
   .O(gates_1021),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1101100110000000101001011000000111001011111111101011100100011000)  
) LUT6_114 (
   .O(gates_1169),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0001111010011010101110000110110101110001100001001110100001010010)  
) LUT6_115 (
   .O(gates_455),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1010010110011110001000001101100101001011101000101001011111110000)  
) LUT6_116 (
   .O(gates_1032),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1100100000011111011111100101110100111111110011001110101110110100)  
) LUT6_117 (
   .O(gates_937),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0100110011111001111001111111100111110001110011101110011001010001)  
) LUT6_118 (
   .O(gates_992),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0000101100101111010011000100000101000011011000100010010000001100)  
) LUT6_119 (
   .O(gates_1368),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0110100101001000111000010110100010011000011010011110101001011010)  
) LUT6_120 (
   .O(gates_1159),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1010011010101111100010001000000000100101011110000001100110001001)  
) LUT6_121 (
   .O(gates_922),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0011011011100001101011100001000110000100101110101001110011000011)  
) LUT6_122 (
   .O(gates_147),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1110010111011111100101111110110100000101001000101100010100110101)  
) LUT6_123 (
   .O(gates_514),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1110110101111011011011001001011110010011111111100010101101010100)  
) LUT6_124 (
   .O(gates_432),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0010001001100100110101100010101001001000001110001110011011010111)  
) LUT6_125 (
   .O(gates_527),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1000011101101110010100000011001000101011110111000100111000000111)  
) LUT6_126 (
   .O(gates_521),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1000011010111100010011100111011011111101000110011010111111111000)  
) LUT6_127 (
   .O(gates_1278),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1100001010001010000100011110010100010101111010000000010010010000)  
) LUT6_128 (
   .O(gates_768),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1010010100101101010011011010101111001101011011101110111010110110)  
) LUT6_129 (
   .O(gates_1244),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0010110011010111001011101000101010100010111111001000001001011101)  
) LUT6_130 (
   .O(gates_916),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0000010000000100010101101110101100111110000100001100000010010011)  
) LUT6_131 (
   .O(gates_909),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0011000111011100010101000010101001100010010101010011101100010001)  
) LUT6_132 (
   .O(gates_859),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1001100011101001111100101110100001001010100101110011001110111111)  
) LUT6_133 (
   .O(gates_242),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b1001100100100011100010001101110000001110100101011110011110100010)  
) LUT6_134 (
   .O(gates_1261),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0100110110110101100111111010110100110000101100111001100011011010)  
) LUT6_135 (
   .O(gates_238),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1001010010101010000100011110111001011110111001110110000010110000)  
) LUT6_136 (
   .O(gates_1350),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0000000010000100010010011111100101100110011111001001011100001110)  
) LUT6_137 (
   .O(gates_725),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1110010101011011100010100110001000000101011001100100011100010101)  
) LUT6_138 (
   .O(gates_59),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0100010001110000010110100000011111000111000100101111011110100110)  
) LUT6_139 (
   .O(gates_1464),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0100100011010000010111011011001011110000010011110100010111000000)  
) LUT6_140 (
   .O(gates_79),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1000110100010110101110111000100000101001011110111000110000010111)  
) LUT6_141 (
   .O(gates_506),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1001100101111110000110101110010100100011010010010011110011001111)  
) LUT6_142 (
   .O(gates_1134),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1100100001110100100100010100011111111000001101010110001010011100)  
) LUT6_143 (
   .O(gates_930),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1010100010101001001010110110011101010000001001000100110110011110)  
) LUT6_144 (
   .O(gates_1482),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0000011010010100011111000000101110000100000101011011011110100000)  
) LUT6_145 (
   .O(gates_1385),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0011111110100100101111110000111100010110100101000010100100011100)  
) LUT6_146 (
   .O(gates_498),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1000111011011110010000111101011000111111011001001100000110111100)  
) LUT6_147 (
   .O(gates_393),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0111101010100011101011110100101001011111111011110100101010010111)  
) LUT6_148 (
   .O(gates_1197),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b0010001000010001001100101101111100101010100011010101001100011100)  
) LUT6_149 (
   .O(gates_656),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0010101100001100011110001101101110001110001001010110010001100001)  
) LUT6_150 (
   .O(gates_1431),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1100110010110110011010010011101001101110100011100100000000101110)  
) LUT6_151 (
   .O(gates_580),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0100100001000110000101000010110010111001101000001101001010010110)  
) LUT6_152 (
   .O(gates_1136),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b0111100010000010111010100101001011100101101110001110101001110010)  
) LUT6_153 (
   .O(gates_524),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1011011110001011010010100001010010011000000110011000100011100101)  
) LUT6_154 (
   .O(gates_778),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0010101100101011000001001001010100111110101001101010001100010010)  
) LUT6_155 (
   .O(gates_763),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1110000110001010001110010111000011011000100111101110111000000011)  
) LUT6_156 (
   .O(gates_444),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b1011010010011010100000011111011001100011110011100001110001011100)  
) LUT6_157 (
   .O(gates_757),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0001011111000001011110101011011000110111011101101101011111100111)  
) LUT6_158 (
   .O(gates_181),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0001100101110010010010100001110001101010000110101000011000101001)  
) LUT6_159 (
   .O(gates_906),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0010110011010010011101001111100001110011101000110111010111111100)  
) LUT6_160 (
   .O(gates_1388),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0101101110100100000100001111010010101111101000000111110011101111)  
) LUT6_161 (
   .O(gates_636),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0010000001001010100010001000000111010000101101100000010101101100)  
) LUT6_162 (
   .O(gates_485),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0000110010110011100101000110011001110011011110100100010110011111)  
) LUT6_163 (
   .O(gates_581),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1111001011101010000000010100010110111001110010100010101101110000)  
) LUT6_164 (
   .O(gates_1539),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0100100000000010111010111101101100011011110011011000011011000111)  
) LUT6_165 (
   .O(gates_1391),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1110011111110011111001010110101010101111001001101110111101110110)  
) LUT6_166 (
   .O(gates_1489),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1001111110110001011111111001010100110101001001101011001010111001)  
) LUT6_167 (
   .O(gates_1299),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b1001110110001100000101111011010001110101100011100110010010010000)  
) LUT6_168 (
   .O(gates_457),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0110000000100100011110001101000011001110010001001011101000101100)  
) LUT6_169 (
   .O(gates_407),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0101110011010101010111010111010011010111110110111100011011111010)  
) LUT6_170 (
   .O(gates_1521),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0010000100101110110111110110111111110101110011100001001011110101)  
) LUT6_171 (
   .O(gates_811),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1101110101011001011111110101110011101001101100011010001101011011)  
) LUT6_172 (
   .O(gates_1027),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b0000100101100110101011000000001101001011111000110101101101100010)  
) LUT6_173 (
   .O(gates_1379),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b1010000000111100110011000111010100111111011000100000110111010010)  
) LUT6_174 (
   .O(gates_1436),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b1100011010110010110011110001111100110000110001010110001010100100)  
) LUT6_175 (
   .O(gates_372),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1101000101010101111110011111000001110100011001011111111111100010)  
) LUT6_176 (
   .O(gates_1234),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0001110110001011010100010101111100100010000100011010100000011101)  
) LUT6_177 (
   .O(gates_1230),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1010001101111111111011110001011111100011111010100011001111000001)  
) LUT6_178 (
   .O(gates_1284),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1011010110100111000000110100100001110101100110011111011100101000)  
) LUT6_179 (
   .O(gates_174),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0101011100110100010010111000110110011010100000000110110001111000)  
) LUT6_180 (
   .O(gates_261),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0100111010110111000110101110111101111001101100100100111111001010)  
) LUT6_181 (
   .O(gates_788),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0011000110011101001101100101011011011000000001011100100100101000)  
) LUT6_182 (
   .O(gates_1120),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1010000001110001110110110000010100110010110010111111110001111101)  
) LUT6_183 (
   .O(gates_17),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0010010011001001110101000011101011010001101110001001110101011011)  
) LUT6_184 (
   .O(gates_793),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1001100101000101111000100100111100011110000110001101111010111100)  
) LUT6_185 (
   .O(gates_673),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1011000111011011011000011001100011101010101101001011011111101110)  
) LUT6_186 (
   .O(gates_446),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0011001011010101010011011110101111000110101001000011011111101001)  
) LUT6_187 (
   .O(gates_433),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0110111000100111010010011001100100001000111101110111010100100001)  
) LUT6_188 (
   .O(gates_1387),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0111010101001111000001100101011101001101010111111010000111001001)  
) LUT6_189 (
   .O(gates_1324),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1001001100110110101001111011011110101101010111011111111110010010)  
) LUT6_190 (
   .O(gates_724),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0001110110110001101011101010000111000000011000000111001001000101)  
) LUT6_191 (
   .O(gates_837),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0110110100000001111101110110111001101110111110001101111001011000)  
) LUT6_192 (
   .O(gates_1425),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1010101011010100011100110011101111011010100001111011011000011000)  
) LUT6_193 (
   .O(gates_1335),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1011011101010000100100101000101111000001001000001110011010011101)  
) LUT6_194 (
   .O(gates_1228),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1110111010100101100110111100101110011100110001010111001101000100)  
) LUT6_195 (
   .O(gates_728),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0101101010011100000001111011001100111010000011111110010011001010)  
) LUT6_196 (
   .O(gates_163),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0111010100010111001000011110101100011100010010100111010111111100)  
) LUT6_197 (
   .O(gates_649),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1110011001001110111000110110010011111110000010001101111111010111)  
) LUT6_198 (
   .O(gates_928),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0111100100111011111111100111000000010010100110101010001100010110)  
) LUT6_199 (
   .O(gates_1318),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1100101011000100000100001001010101001011111010001000001110100111)  
) LUT6_200 (
   .O(gates_1256),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1011000011010011101001100000001000000000111001010110011000000110)  
) LUT6_201 (
   .O(gates_78),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1100110110111110000001011111001001100101010000100001101000010101)  
) LUT6_202 (
   .O(gates_1044),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1000100110010101110101000001001001001010101011111010011101001101)  
) LUT6_203 (
   .O(gates_183),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b1110110001000010100111001100010010101110001011001011000111010011)  
) LUT6_204 (
   .O(gates_594),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1111100011100010010110110101000001010011111111100100011110011010)  
) LUT6_205 (
   .O(gates_697),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0000001011001110110000110111011000100001011101011110100001101111)  
) LUT6_206 (
   .O(gates_775),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0111100110011001000010101000101000101101001010110000110101110100)  
) LUT6_207 (
   .O(gates_1178),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1000111101100111101110001100100010000110011010001001100110000011)  
) LUT6_208 (
   .O(gates_699),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0001111010000100111000001110010010110010010000101010001010000100)  
) LUT6_209 (
   .O(gates_565),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1100010101001100011101101000001001110000111000110110101111001000)  
) LUT6_210 (
   .O(gates_1166),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1111110110010110000101111001010110100100111101100010101010110101)  
) LUT6_211 (
   .O(gates_628),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0101110000101000000111100111101101001010010110000010001100111100)  
) LUT6_212 (
   .O(gates_629),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1000111010001110101001111000110000011100011011000011010100001001)  
) LUT6_213 (
   .O(gates_1493),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0100110000110111101110100111101001011111010100010010100011100101)  
) LUT6_214 (
   .O(gates_688),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b1010011111011111001111000101100111011001010011111100000101001110)  
) LUT6_215 (
   .O(gates_764),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0100101110110111111100110000001100101101011101001000111010001000)  
) LUT6_216 (
   .O(gates_815),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1011100110111111011110100110010011010000011100011010000100001110)  
) LUT6_217 (
   .O(gates_612),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1101100010010110010101111000100100100111101100100110011101111111)  
) LUT6_218 (
   .O(gates_1352),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0010001011000101000101010001010010011111110011001100100111100101)  
) LUT6_219 (
   .O(gates_1116),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b0110111001100000010011101101001000100101001100000111100001000011)  
) LUT6_220 (
   .O(gates_394),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0011111010000111110101110011001100000000101101011111010111100001)  
) LUT6_221 (
   .O(gates_285),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1100100111110110111101011110000010011111110100101011100101000011)  
) LUT6_222 (
   .O(gates_1481),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1101100101111000000001000010111000011011010111001011010010101110)  
) LUT6_223 (
   .O(gates_1488),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1001011010100100110000010101010001000011010011010001011111010001)  
) LUT6_224 (
   .O(gates_831),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1001100000111101011100101000000101001000001111101111111101101101)  
) LUT6_225 (
   .O(gates_1483),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0110100101000110101101110001111101001011011001010110001100011010)  
) LUT6_226 (
   .O(gates_1499),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b1011011010010000110110111111110111011101110110100001011000000101)  
) LUT6_227 (
   .O(gates_709),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1000001110000111010010100111011010100011100111011101110011101100)  
) LUT6_228 (
   .O(gates_1449),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b0110110101111101101011011101111111001111110001110001111010010111)  
) LUT6_229 (
   .O(gates_929),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b1001100100001011010011010101101110000111100111010001010001001111)  
) LUT6_230 (
   .O(gates_1515),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1100011111000110000000110010101110111111101010000000110011000011)  
) LUT6_231 (
   .O(gates_23),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0101001010110011111001001000101010110010110100011100111111111010)  
) LUT6_232 (
   .O(gates_1163),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0010111011011110011111000001001101000110010000100101000001010000)  
) LUT6_233 (
   .O(gates_858),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0011110001110100111000111001100100101010010011100000111111100100)  
) LUT6_234 (
   .O(gates_1422),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0110000101101000011110000111001111000101110101100010100000001111)  
) LUT6_235 (
   .O(gates_1147),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001000000011000110110100000101111000010101101111001000000000101)  
) LUT6_236 (
   .O(gates_43),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1100101110111100100101011001011011111001010100110111100011011110)  
) LUT6_237 (
   .O(gates_726),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0011010111001001101100111001001100001000101110111010001110001010)  
) LUT6_238 (
   .O(gates_1496),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1000011101010111010101100011001010111000110000110010100001111011)  
) LUT6_239 (
   .O(gates_475),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1000111001101111111010101111100110111000001101011100100100110000)  
) LUT6_240 (
   .O(gates_752),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1000111110111000000000000000110111000110011001010011011110011110)  
) LUT6_241 (
   .O(gates_1330),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1010010110111000000011101010111101011101111001101011101110100010)  
) LUT6_242 (
   .O(gates_177),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0101111111010110100101011000110001100010111110111100111000010100)  
) LUT6_243 (
   .O(gates_468),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1010010110010010100101001010101111001101000100000111011111110010)  
) LUT6_244 (
   .O(gates_1487),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1010010111000011110001011010101010001100011110101111000110000110)  
) LUT6_245 (
   .O(gates_823),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1001100001000100011111100101101000101011011001001100100010011101)  
) LUT6_246 (
   .O(gates_185),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1011001110101101001101011001101101110011001001101010011101110110)  
) LUT6_247 (
   .O(gates_219),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1100001100100001000010010010100100110111000010010000101110110101)  
) LUT6_248 (
   .O(gates_70),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b0011111100000110011000111111110011011001111101010001111011010111)  
) LUT6_249 (
   .O(gates_1382),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0000101110101010110110111110001110011100110001000010101000110111)  
) LUT6_250 (
   .O(gates_1239),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1110101100101011101011100110011010110111111111010100101100101010)  
) LUT6_251 (
   .O(gates_1452),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0011000010001100111000100000011010101110001100110111100101011110)  
) LUT6_252 (
   .O(gates_1401),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b1011011101011010000010111110111110110010011001110101101001011000)  
) LUT6_253 (
   .O(gates_745),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1000101000000100011100110100011000011000011000000101011101101111)  
) LUT6_254 (
   .O(gates_1506),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0111011110001000011000000011110110000010010001101001000101010111)  
) LUT6_255 (
   .O(gates_533),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b1011001100001000000010000110001010111110011100111010111001100011)  
) LUT6_256 (
   .O(gates_1014),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0011000101101010110100001111101101111011000111011100111110011111)  
) LUT6_257 (
   .O(gates_95),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1111100100011101010111110110110111100010110100000101101001001010)  
) LUT6_258 (
   .O(gates_642),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1100110111111111000000010011011110000011010001000111010010111000)  
) LUT6_259 (
   .O(gates_543),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1111110111010001101110001010111000101110110101001001000100001101)  
) LUT6_260 (
   .O(gates_1375),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1100011000001000001011000001100100100001000000100111111110000001)  
) LUT6_261 (
   .O(gates_1220),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0001110010101010110010011110100000000100111110100100110011000011)  
) LUT6_262 (
   .O(gates_718),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1010010100000000000010100111001110010010100100110001101100011001)  
) LUT6_263 (
   .O(gates_166),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0011110011000101101111111000001101001011101100101010011101110000)  
) LUT6_264 (
   .O(gates_324),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1100111110101000011000000001100001100111100101010000000001011001)  
) LUT6_265 (
   .O(gates_158),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0011101000110111001110011011010101011000101011111010100101110100)  
) LUT6_266 (
   .O(gates_622),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001011110100111101100010110101001110010101110101011000110011011)  
) LUT6_267 (
   .O(gates_537),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1111011000010011100101011000110000000101001000001000100011101100)  
) LUT6_268 (
   .O(gates_263),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1111000000011101111010000010111000001001000010010110111101001011)  
) LUT6_269 (
   .O(gates_1052),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0100111110011110111001011010111011001110000001011111111111101000)  
) LUT6_270 (
   .O(gates_1316),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0001101101000101000000100011011011000111111010101100110001001010)  
) LUT6_271 (
   .O(gates_1351),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0110011001001100011100011100111010100000000000010001110001100000)  
) LUT6_272 (
   .O(gates_150),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0010110010011011011111110111111111111010000011110110010000110110)  
) LUT6_273 (
   .O(gates_1175),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0000101110100010010101101101111101011110100101000111010100100110)  
) LUT6_274 (
   .O(gates_260),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0101011100110000000110000011101101010001100000011001000111001100)  
) LUT6_275 (
   .O(gates_1064),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0011111011101001000011010100000011100101000110100111110011111111)  
) LUT6_276 (
   .O(gates_927),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1011011011110011100101011110100000001110110000011001010101100100)  
) LUT6_277 (
   .O(gates_1491),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1011010100101011011110111011000001101110000101011001100111110011)  
) LUT6_278 (
   .O(gates_963),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1110010100011111011111101101011010010000100101010001010111001010)  
) LUT6_279 (
   .O(gates_1182),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0010111001111000011000000011000001000001010011000101110101000011)  
) LUT6_280 (
   .O(gates_574),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0100010101000001000101111100101001011110011010101010001101100001)  
) LUT6_281 (
   .O(gates_1236),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1011001011100011000100110111111101011001111101011110000000011000)  
) LUT6_282 (
   .O(gates_555),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b1011010100011000101011110110101001011101011000011101111100110010)  
) LUT6_283 (
   .O(gates_1522),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1011111001110110001011011100101101101111110101010000111001011111)  
) LUT6_284 (
   .O(gates_1008),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1111110111101111001000100100110110000101001000011010111010100001)  
) LUT6_285 (
   .O(gates_503),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1000000101110100011001110110101010111011110011001101011101110000)  
) LUT6_286 (
   .O(gates_735),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0111001000100100011100111000001010001111010111101000001111000000)  
) LUT6_287 (
   .O(gates_520),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1100000010001000101101100111011011010100101010110111110001011101)  
) LUT6_288 (
   .O(gates_1276),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1011001100111100110110110001110011001001101111010000100111001010)  
) LUT6_289 (
   .O(gates_1012),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1110110110111110101001010110110011001010101100001001111110100100)  
) LUT6_290 (
   .O(gates_447),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0111111101101100010000111000000010110011011011101001111111001010)  
) LUT6_291 (
   .O(gates_784),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1111010000011001011101110100100001011101001100101111101100001100)  
) LUT6_292 (
   .O(gates_679),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0010110011011101101110100001001110100100101000001000100010011011)  
) LUT6_293 (
   .O(gates_497),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1000101111000001110010001010010001100011010010110101100000000001)  
) LUT6_294 (
   .O(gates_891),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0100000000011101101100111001010100111001100110000110001001001000)  
) LUT6_295 (
   .O(gates_19),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1110100000111010100100011100111100010110001001010011101000100110)  
) LUT6_296 (
   .O(gates_1125),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1001110111010010010101101010011110100010101100110000010010000001)  
) LUT6_297 (
   .O(gates_779),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1001101111001000101111010100100010010101110001100101111010110011)  
) LUT6_298 (
   .O(gates_1469),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0011111100010111011101100011110101111110000111011010100001000101)  
) LUT6_299 (
   .O(gates_405),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0100110011000101000110010111011011000000100000101110001000001001)  
) LUT6_300 (
   .O(gates_1461),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0010001001110101010000111101110101010101010111010101001100101010)  
) LUT6_301 (
   .O(gates_1281),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0001110010001110100001111100111100101011101001011000010001100001)  
) LUT6_302 (
   .O(gates_780),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0111011111111101100111001000101111001001001001011100001100110000)  
) LUT6_303 (
   .O(gates_1078),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1010111111101001110110011100101001010000010010000001000001101111)  
) LUT6_304 (
   .O(gates_442),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b1010011110110011111000001011011100010100010010010011110010001001)  
) LUT6_305 (
   .O(gates_1550),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1011111110100111110010101001001111110010100101100101010100001101)  
) LUT6_306 (
   .O(gates_1484),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1001110001000101010010101111111101000101100000001010001101000000)  
) LUT6_307 (
   .O(gates_988),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1001001101100110000000011111010010111010010001001010101000011011)  
) LUT6_308 (
   .O(gates_1430),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1010010100011111110001001101001000101110110110101101001110111110)  
) LUT6_309 (
   .O(gates_722),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1101101101111100000010011001010101001110011001010011000010101110)  
) LUT6_310 (
   .O(gates_1536),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0111110111100010111101010011001010101100110010001001000111010001)  
) LUT6_311 (
   .O(gates_923),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0111000010001111010110100111101111100101001011100110101011010000)  
) LUT6_312 (
   .O(gates_309),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0110011011001100111011110111011101001101100000111011110001100100)  
) LUT6_313 (
   .O(gates_401),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1110111010111001011010100000010101110011000001000111010101110000)  
) LUT6_314 (
   .O(gates_1371),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1101011011011101000100110101110100010111111101001001110100010100)  
) LUT6_315 (
   .O(gates_846),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1010110110100101111001110110110011001011001000110100110101000110)  
) LUT6_316 (
   .O(gates_995),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1011011000110001111110011101000011011011111011111000011010101110)  
) LUT6_317 (
   .O(gates_867),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0111100001111001011101100011111001110010111101111010110001011111)  
) LUT6_318 (
   .O(gates_695),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0000001001011001110101010000011011011111110000010010110101010110)  
) LUT6_319 (
   .O(gates_154),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1110100100000001000011100110110111001011100000000100100111110010)  
) LUT6_320 (
   .O(gates_1113),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0101001000000000000000000000010000100000111000100111100010010101)  
) LUT6_321 (
   .O(gates_1003),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0010010011111000000001011011101001000001111000010000001011001101)  
) LUT6_322 (
   .O(gates_1059),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b1111000100011010010110100101001111100001111101011001011111101011)  
) LUT6_323 (
   .O(gates_1187),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0010100011010111000010111010010110010000011010000010101000000000)  
) LUT6_324 (
   .O(gates_999),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b0110010110001110001000000100011011100000011110010010000110001111)  
) LUT6_325 (
   .O(gates_65),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b1101011000100001000001101101011010101000000010010101101100110010)  
) LUT6_326 (
   .O(gates_711),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0110110111100100011011001111011111000110100111100110011011100101)  
) LUT6_327 (
   .O(gates_1031),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0000110000100101100110101101011010100100010111110011000001010001)  
) LUT6_328 (
   .O(gates_1226),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0001010010101001110000011100010101110011010110001101101011111001)  
) LUT6_329 (
   .O(gates_294),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0101111111110111101001000101001100101000010011010111001000110000)  
) LUT6_330 (
   .O(gates_1444),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b1110011110100000111100000001110111010110010100011100001100000110)  
) LUT6_331 (
   .O(gates_873),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001001110110101101100001001000010111111010001010000111011011001)  
) LUT6_332 (
   .O(gates_1288),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1000000010001101111001010101000000100111001001111001000010000110)  
) LUT6_333 (
   .O(gates_663),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0111010100101110010100101100011100001100100010000011111110100110)  
) LUT6_334 (
   .O(gates_1344),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1011011110101110001010101011111011001100001101111000011001000010)  
) LUT6_335 (
   .O(gates_1202),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1010010111111111011000101000100010010101001110010100110000100100)  
) LUT6_336 (
   .O(gates_1176),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0101011001001111011110111011010111101110000101001010110100101110)  
) LUT6_337 (
   .O(gates_161),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1100111111001010000110010001011001011110010101101100000111101110)  
) LUT6_338 (
   .O(gates_1447),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0000101000011110001001000000110001110010011110010111001000101111)  
) LUT6_339 (
   .O(gates_344),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1110110000000000011011000000110000110010110100010100001010110011)  
) LUT6_340 (
   .O(gates_634),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b0101111010101010010011101000110100101111011100001111011100000111)  
) LUT6_341 (
   .O(gates_93),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0011011011011110110101111111011110111111011000010011100010111001)  
) LUT6_342 (
   .O(gates_1248),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0110000000110000111001100101001100010101001111101100001100000010)  
) LUT6_343 (
   .O(gates_1513),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1100010001001110101100110111001111110010100001000010010111010011)  
) LUT6_344 (
   .O(gates_501),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1101001110111010011010010100010000011011011010011000101111100101)  
) LUT6_345 (
   .O(gates_379),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1001100011101000001010100110011100000010111011001110010001110110)  
) LUT6_346 (
   .O(gates_1277),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1001110011000011110110000010110010110000010011010110001110011000)  
) LUT6_347 (
   .O(gates_368),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0001011010110011001111001011100010011000111111001001101001101010)  
) LUT6_348 (
   .O(gates_665),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0010011010110101000110110000111010001010010101101110100111111110)  
) LUT6_349 (
   .O(gates_621),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0011101001100101001011100111010000010110100100101000110011000100)  
) LUT6_350 (
   .O(gates_1231),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1101011100011111101110110001110111011001111010011111000001100101)  
) LUT6_351 (
   .O(gates_569),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0101011110110010011101110000110010100001011010110001100001110101)  
) LUT6_352 (
   .O(gates_1337),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b1100100011000010110110111110011011001000010001000111111010111010)  
) LUT6_353 (
   .O(gates_208),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0110000011110011101111101111011001101110101101010001011100111111)  
) LUT6_354 (
   .O(gates_11),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0100101100110001101001101001000111011001111100001001101010101100)  
) LUT6_355 (
   .O(gates_1005),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1100001100010100101011100011111001100111101010000100101011000100)  
) LUT6_356 (
   .O(gates_1282),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0000111000101110111011110010101000001100111011100010010010111100)  
) LUT6_357 (
   .O(gates_412),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1100100100111100111110101111011100011100101101111100111110001100)  
) LUT6_358 (
   .O(gates_616),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000111011001101100010100111010010111101111000001011100110110101)  
) LUT6_359 (
   .O(gates_536),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0100010001000110001011101001111110101101011110000111011010101011)  
) LUT6_360 (
   .O(gates_813),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1101000111001010101101010110011010000001000100011111011110010000)  
) LUT6_361 (
   .O(gates_72),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1110110000101101010101100010011101001111001110111101110010011010)  
) LUT6_362 (
   .O(gates_1164),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001100100100011101001110010111010001000110000011001001010011110)  
) LUT6_363 (
   .O(gates_1145),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1111000101000110011101100000010110111111110001000011110000011000)  
) LUT6_364 (
   .O(gates_954),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1010100011100001001011001100100101100001100010001110001010100000)  
) LUT6_365 (
   .O(gates_857),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b1000110000101101011110101011111001111001000110100101111001011100)  
) LUT6_366 (
   .O(gates_640),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b1110001101110001011000000111000001000000011001000111001100011001)  
) LUT6_367 (
   .O(gates_262),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1011011101101100100001101010010010110100011000110100100001000001)  
) LUT6_368 (
   .O(gates_1404),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0101110100100011111001000100010110001001111110110110011101101000)  
) LUT6_369 (
   .O(gates_1395),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1111010100001111011101010100010101011110010110000111101111101000)  
) LUT6_370 (
   .O(gates_967),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0000001001010110111101011111110110110100100001000010000010010000)  
) LUT6_371 (
   .O(gates_959),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0100010100100100100110101000010010000011000110011110110111100111)  
) LUT6_372 (
   .O(gates_1172),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1001111100001101011110001100010110011101010111100000101111011011)  
) LUT6_373 (
   .O(gates_919),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0001001001001100011011011010010101011001010000110001000101111011)  
) LUT6_374 (
   .O(gates_1541),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1000111010001000010111101100101010100010010110111101110000011110)  
) LUT6_375 (
   .O(gates_917),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1001010010001100100101110000000001111111101110110011110001111110)  
) LUT6_376 (
   .O(gates_463),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1010001000110110011100111001000011000110100100010100101001111010)  
) LUT6_377 (
   .O(gates_707),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0001000010010111101111100011100011000001001110001000010010111100)  
) LUT6_378 (
   .O(gates_860),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b1111100101100010001111110000010000101000010000001101101110011010)  
) LUT6_379 (
   .O(gates_703),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1101101111001100001011101011110011101001100101111010011101100111)  
) LUT6_380 (
   .O(gates_1523),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0111011001011100000010001000010000100110100111010101001100000001)  
) LUT6_381 (
   .O(gates_1336),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0010100111001101010101000000111110100100101011100110000011011010)  
) LUT6_382 (
   .O(gates_291),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1110110101000110100001010110100000010011111011001000111011010010)  
) LUT6_383 (
   .O(gates_1507),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0011010101100111011001010101001001101100010011011111011110100111)  
) LUT6_384 (
   .O(gates_1300),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1111100111001011111001001000001010101101001010001111010110010110)  
) LUT6_385 (
   .O(gates_886),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0110001110010101100000001001010101010101010010110101100000111101)  
) LUT6_386 (
   .O(gates_1474),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0110011001011000001001010100001011011001000011000101010010000011)  
) LUT6_387 (
   .O(gates_646),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1100111100011010000011011010000011110010101110000111100110101001)  
) LUT6_388 (
   .O(gates_1127),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0111001101100000110001010111000110111010000110110100100011000100)  
) LUT6_389 (
   .O(gates_1265),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1101110010001000110101001011011101111000100000001100001001010010)  
) LUT6_390 (
   .O(gates_320),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1111001000010100010110111011111010000100110000111011100000011101)  
) LUT6_391 (
   .O(gates_659),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0010000000100001001110101011111010000001011100010000000011100000)  
) LUT6_392 (
   .O(gates_1527),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0011000011100110110010110111000110010011110111101001111101000001)  
) LUT6_393 (
   .O(gates_739),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1110100100100111100101100101000111111001100111101001011100001100)  
) LUT6_394 (
   .O(gates_557),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0001100101110111111010010001000110110011100110001011001101110011)  
) LUT6_395 (
   .O(gates_3),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0101100000110101100001111001100010001000101111111001101001101111)  
) LUT6_396 (
   .O(gates_1095),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1100100100001110001010010111000010111011000100101111101100111111)  
) LUT6_397 (
   .O(gates_789),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0100100000100010110100000111100110111011001111100100111111101110)  
) LUT6_398 (
   .O(gates_1062),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1001100010111101000011110100001010100100001100101001100101101000)  
) LUT6_399 (
   .O(gates_897),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1101001110011101110001110100101111110011001111011000010101100111)  
) LUT6_400 (
   .O(gates_1057),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b1110011001001111100000110110001011111110101010110010010010111100)  
) LUT6_401 (
   .O(gates_354),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1100011011011011000010110010111101100010000111011010010001001110)  
) LUT6_402 (
   .O(gates_329),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1101011010101110011111110010001100000011011010000010110101010000)  
) LUT6_403 (
   .O(gates_105),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1100101000110111011110010001100111110001101110100101111001100100)  
) LUT6_404 (
   .O(gates_560),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1000001000100110001111111010111101101100111010010010011100101110)  
) LUT6_405 (
   .O(gates_839),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1010010101011111001100011101001001000010011000001101010001001101)  
) LUT6_406 (
   .O(gates_633),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0101110100101100100101111001111100010111101010100111011011111111)  
) LUT6_407 (
   .O(gates_544),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0110001100001011110000000110001011011000111011001111000001010101)  
) LUT6_408 (
   .O(gates_1466),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0000101000111111011011111000010001010010000001000011010101001111)  
) LUT6_409 (
   .O(gates_102),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1010110100011001101111000100110000111000111111011000011111011110)  
) LUT6_410 (
   .O(gates_690),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0110110100111100111001010111000010110101010001101001010111011011)  
) LUT6_411 (
   .O(gates_357),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1000101111100001001111010010111000110100011111011001101010010100)  
) LUT6_412 (
   .O(gates_731),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0000101001011001001110000111110111101101100001011111010101110110)  
) LUT6_413 (
   .O(gates_670),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0101100011000111101110101111111000011100000010101011101011011000)  
) LUT6_414 (
   .O(gates_1298),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0001011010100101001010111100110101000000100000110100110011010111)  
) LUT6_415 (
   .O(gates_441),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1101110110110010011101101101001101101100101000110010110101110111)  
) LUT6_416 (
   .O(gates_1497),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1110111110101111000101010010111111000110011010000110100111111101)  
) LUT6_417 (
   .O(gates_138),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1010100101001011011101001111100001101001011001011100110101100001)  
) LUT6_418 (
   .O(gates_483),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0100111011001111110100011010101000110011001010001111000100100001)  
) LUT6_419 (
   .O(gates_647),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1100001001101100010111011010010011001111011100011100010111100010)  
) LUT6_420 (
   .O(gates_84),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1001000111101101100111111011011000100101111111111100010111010000)  
) LUT6_421 (
   .O(gates_113),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0001011110111000111110101110101100001100101001101000010000001000)  
) LUT6_422 (
   .O(gates_568),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1110101000110010010111001010110001111100110111101111100101110011)  
) LUT6_423 (
   .O(gates_173),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0111111011101001010011111110100000000010111110101110110100100101)  
) LUT6_424 (
   .O(gates_797),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0010110010000000101001111001100000000001101000100011110101000011)  
) LUT6_425 (
   .O(gates_350),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0011010010010110110001000011000010001110110110011111001110000010)  
) LUT6_426 (
   .O(gates_267),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b1010110100001111011000100000011001111100010011010010100000111010)  
) LUT6_427 (
   .O(gates_1420),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0000101110111110110001010001111001100000001011011001101111010010)  
) LUT6_428 (
   .O(gates_608),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0000010010001110100000011101000010011111111111001101001000000000)  
) LUT6_429 (
   .O(gates_6),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1000001100001110001100000010010000001110101001001010110010110111)  
) LUT6_430 (
   .O(gates_103),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1101111101011000110001011000100111100100110001001110111000110010)  
) LUT6_431 (
   .O(gates_871),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0101001000001110101101010001100100010100101110111111000101111011)  
) LUT6_432 (
   .O(gates_597),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0100101000001100010011000000100000111111011000111000010101011111)  
) LUT6_433 (
   .O(gates_599),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0001000101100000101011010101000011010000011001111101111010010101)  
) LUT6_434 (
   .O(gates_675),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1100001110110011011111000101011100101111001000100001010110011000)  
) LUT6_435 (
   .O(gates_806),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0011011110100100011111111001100111100010001000010101101011010100)  
) LUT6_436 (
   .O(gates_228),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1100100100001110101100111111001101110101001000010100010010000111)  
) LUT6_437 (
   .O(gates_1104),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0100010100001001110100111010000100111011111101101011010011111000)  
) LUT6_438 (
   .O(gates_1504),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1001111110101101011000100011010000110001100010111010101011011101)  
) LUT6_439 (
   .O(gates_359),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0110010111000010110001100010011011011000100100110101100111110101)  
) LUT6_440 (
   .O(gates_1100),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1001011000011001110000010101111100111101111000110010011111000101)  
) LUT6_441 (
   .O(gates_799),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1000000010010001110100000000101100000010111011000010110010111011)  
) LUT6_442 (
   .O(gates_802),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1001010001100010010011000101100111100000001111011000001111011111)  
) LUT6_443 (
   .O(gates_1473),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1110001111100010001010001001000101001110101001111001011110101000)  
) LUT6_444 (
   .O(gates_142),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0001100111011001111100110100001011101101001110111110010000100001)  
) LUT6_445 (
   .O(gates_1546),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1010111111010110100110001011001110101001100000111111110011100011)  
) LUT6_446 (
   .O(gates_1101),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1111100011001001100110111001010100101111000101111101010001000111)  
) LUT6_447 (
   .O(gates_717),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0111100010000010101000101001000100001101110101101100001011001010)  
) LUT6_448 (
   .O(gates_336),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0111011010001011111100000011111000010001001011001000000101110100)  
) LUT6_449 (
   .O(gates_479),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1101100001011110100000101000010111011001000001010101001111011110)  
) LUT6_450 (
   .O(gates_426),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1100001001101111000000111100011001011001001100011110011100011110)  
) LUT6_451 (
   .O(gates_332),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b0000110001110000000111100000111100110010011000000000111010011000)  
) LUT6_452 (
   .O(gates_1069),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1110010010000000001101101111100001011110101011101111000000001101)  
) LUT6_453 (
   .O(gates_721),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0100001001111011110110111100100100101011101101101000100011000101)  
) LUT6_454 (
   .O(gates_1267),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0101100010011110010000110000010100110100110000001010000111101001)  
) LUT6_455 (
   .O(gates_625),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b1100010111010101100110011010110100011011110101001101100101010100)  
) LUT6_456 (
   .O(gates_272),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0111111110011010001011110100100011001001011101011001110110000101)  
) LUT6_457 (
   .O(gates_345),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0110101000011010110010100101001111111001010010001011100100011010)  
) LUT6_458 (
   .O(gates_805),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0110100101111011100011110001111010110111001011111011010110100010)  
) LUT6_459 (
   .O(gates_1198),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1111101011111000101111100010001001110110101101101101110100110000)  
) LUT6_460 (
   .O(gates_504),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1010101101001100011011001110101011011011010010010100111010011110)  
) LUT6_461 (
   .O(gates_1325),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0111110010000110011100100000001010101100111011010010010101101100)  
) LUT6_462 (
   .O(gates_1097),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b1100011000010000111001111100001011111011000010101111010100100110)  
) LUT6_463 (
   .O(gates_415),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0100111000000010101111110100110100011011010100001101100101100100)  
) LUT6_464 (
   .O(gates_1170),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0001010010110001101000011001100111001111111100110100001110110010)  
) LUT6_465 (
   .O(gates_1406),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1011010011010101111000010100111000110010110111100101011001110000)  
) LUT6_466 (
   .O(gates_1448),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1100110100100110111001001000100101010110101100110110111011111011)  
) LUT6_467 (
   .O(gates_316),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0100000110011110110001100010101101000000111011011011110101100110)  
) LUT6_468 (
   .O(gates_667),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0000111011011001011001101100001000001010111100001111101000100010)  
) LUT6_469 (
   .O(gates_448),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0111100001101100000100001111100111000010110101001111000111101011)  
) LUT6_470 (
   .O(gates_1355),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1010111011100001000010011000110010100100010111111111101100011001)  
) LUT6_471 (
   .O(gates_614),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0010011011111001000110101110011111000111101000010110111010101010)  
) LUT6_472 (
   .O(gates_687),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1111110000100101000111101011000011100011001100110001101010101100)  
) LUT6_473 (
   .O(gates_264),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1111011101111000110011100111101001101111111011001100011010001100)  
) LUT6_474 (
   .O(gates_1106),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b1110101000000001011101001101001000010011000101100100010100010101)  
) LUT6_475 (
   .O(gates_638),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1010000111000001110000000010011110101010001100110111000011111110)  
) LUT6_476 (
   .O(gates_531),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0011011111000010110001001111011111100110000101001111010011111111)  
) LUT6_477 (
   .O(gates_1389),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0010110110111000100111001100011010011010101000000110000010110011)  
) LUT6_478 (
   .O(gates_306),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0100100100110101111110110101110000110110001001011101101011001100)  
) LUT6_479 (
   .O(gates_118),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0001100011001111111110011000110101011111101001110110110110001001)  
) LUT6_480 (
   .O(gates_326),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1110000010010011010001110010000011100111110101010110101001100101)  
) LUT6_481 (
   .O(gates_877),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0100001010001011100110001101010100101101000011100000000011111110)  
) LUT6_482 (
   .O(gates_825),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0111010010110110001101000101101011111011000010000000110000000001)  
) LUT6_483 (
   .O(gates_237),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1001000110101011110001001011111011011111101011000101000011100110)  
) LUT6_484 (
   .O(gates_1495),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1001011001111000001101001100111101101011010000111010111101100110)  
) LUT6_485 (
   .O(gates_1041),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0101000100101010100111011000010010011100010101001110110110110011)  
) LUT6_486 (
   .O(gates_51),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1100100110100100000111101010110010011100011001101110011011000000)  
) LUT6_487 (
   .O(gates_169),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0011001001100100000101100111111000010110000111101110011111100111)  
) LUT6_488 (
   .O(gates_666),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1011000100110001001000110001011100100001001011001001110110110100)  
) LUT6_489 (
   .O(gates_639),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0010110110001110010001110101010111001000011010101001010000101101)  
) LUT6_490 (
   .O(gates_197),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1110011110100110010001010110000010101111111101111111110000100110)  
) LUT6_491 (
   .O(gates_38),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b1110000001100101100011111001010101010110001010011001011100101110)  
) LUT6_492 (
   .O(gates_912),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1111100101011110010000000010110110000111100011100000011100001010)  
) LUT6_493 (
   .O(gates_938),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0011110101011101101101000110110110110001010111010001101011000100)  
) LUT6_494 (
   .O(gates_1255),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1101111100000010110101111001110001000001100010000101001001001111)  
) LUT6_495 (
   .O(gates_1099),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0101111110111100111000100001001011000110110100000110110001010100)  
) LUT6_496 (
   .O(gates_1372),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b1111111011011011100000001001011000111001001111101011101001001110)  
) LUT6_497 (
   .O(gates_592),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1011010001001110110111010000100011001100111011111010011000011100)  
) LUT6_498 (
   .O(gates_1199),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1000101100101000000000010011001110110000010000111110110001111000)  
) LUT6_499 (
   .O(gates_1215),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0100010111001000000001110011101110100001010110110110101111000001)  
) LUT6_500 (
   .O(gates_681),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1000100101001100011000100010000001110010100000011101110000100111)  
) LUT6_501 (
   .O(gates_289),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0100101001101101101100001111011101001010001001111111100101110111)  
) LUT6_502 (
   .O(gates_1227),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b1010111111010111010101101010001110001010010110010011001101011111)  
) LUT6_503 (
   .O(gates_1357),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b1110010010000101011001011010011001010110101000000100110110111010)  
) LUT6_504 (
   .O(gates_210),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0001101111110011001100101110011011100100010100010010110101101011)  
) LUT6_505 (
   .O(gates_1128),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1001000000101001011000010101001110010100100101001110111111011100)  
) LUT6_506 (
   .O(gates_895),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1111010111110010110001011010111011000101100010011010000101110101)  
) LUT6_507 (
   .O(gates_630),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b0001001011101011100111010000110111000110010111110010010100001101)  
) LUT6_508 (
   .O(gates_865),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1101100111110110101001000010000000111110100001010011110011101010)  
) LUT6_509 (
   .O(gates_528),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0100100001000100011110111111011010110111100100001110111011010011)  
) LUT6_510 (
   .O(gates_477),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0010000110010011111110010010000111100000100101011111110000100001)  
) LUT6_511 (
   .O(gates_1055),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0100011011000001010101111100000111011110111111110101101101010001)  
) LUT6_512 (
   .O(gates_1364),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0000110111100100000110101011110110111110000000000011111010010010)  
) LUT6_513 (
   .O(gates_400),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1011101001100001111010001100111000000000000001110001110111001000)  
) LUT6_514 (
   .O(gates_1219),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0000101100111010001011001001011000001111101011011001000010011011)  
) LUT6_515 (
   .O(gates_1542),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0100010011000011010110010010101000110001100010000011101110100001)  
) LUT6_516 (
   .O(gates_116),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1111001100101000010110011010100110000011111100000001000000011111)  
) LUT6_517 (
   .O(gates_976),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0001110011001101111011111011101100110001110110110110001101001011)  
) LUT6_518 (
   .O(gates_1434),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1010100000101110010100011011000001110110011110010001110111101011)  
) LUT6_519 (
   .O(gates_1253),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0000101100011101000010000110000100000100000011011111001100001011)  
) LUT6_520 (
   .O(gates_429),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0001111000000011011000111111111001100001100011010011101101010111)  
) LUT6_521 (
   .O(gates_60),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1011001110101110111000010010110100101100110011000001000011000001)  
) LUT6_522 (
   .O(gates_546),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0101000011001010111100001001010000100110111100000000011111001101)  
) LUT6_523 (
   .O(gates_767),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1010101100101110101001110001110100110111001000000110111110110001)  
) LUT6_524 (
   .O(gates_63),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1010110001001001010111111110100101000010000111010101001011100001)  
) LUT6_525 (
   .O(gates_1023),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1010001111001100001100011111000001011011000110011001000111001100)  
) LUT6_526 (
   .O(gates_29),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1000111000111100101101111111000111011000011000111000110101001110)  
) LUT6_527 (
   .O(gates_874),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0011100000011001011011001110001100011011110111101111011011100110)  
) LUT6_528 (
   .O(gates_677),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1000100100000101101011101010111000101011011100001010011010000110)  
) LUT6_529 (
   .O(gates_1140),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0101010011001110101100010011000010000100010000001001011011000110)  
) LUT6_530 (
   .O(gates_466),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0001110111001000001010011000000000001101111001101111101100111100)  
) LUT6_531 (
   .O(gates_126),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1010001111000001111101011011100000000101001001111100011000001010)  
) LUT6_532 (
   .O(gates_321),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1101001010110000010100010001000010011111001011010100000010110101)  
) LUT6_533 (
   .O(gates_456),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1000001100101110110100001001101011100001110000000110110000101011)  
) LUT6_534 (
   .O(gates_975),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0001111011001011010010110011110011000111000001001001110111100101)  
) LUT6_535 (
   .O(gates_1063),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0110000100111010001011011100101101000001101001010101000001010000)  
) LUT6_536 (
   .O(gates_875),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1100011011101010011000000011100111010110001010001100001001000000)  
) LUT6_537 (
   .O(gates_254),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0110001110100101000010010001011000010001010010101100101001110001)  
) LUT6_538 (
   .O(gates_809),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1000101010111110100101101000010001000010001100011111000100101010)  
) LUT6_539 (
   .O(gates_61),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1111110100111101010001101000110001100001001011100011010101001110)  
) LUT6_540 (
   .O(gates_576),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0101100110101100100010111001000011110101101010110100011110010101)  
) LUT6_541 (
   .O(gates_1510),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0010110001001100101011010110011011010010100011101100101011001011)  
) LUT6_542 (
   .O(gates_894),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1101100001101000000011010101001111011100101001001001000111011000)  
) LUT6_543 (
   .O(gates_712),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b1111000000001001100011010010001100011110010110111011110011001111)  
) LUT6_544 (
   .O(gates_710),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0100001010011000111101101000011010001010110110000011100110100100)  
) LUT6_545 (
   .O(gates_1287),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1110110011110101011100001011101101100110001110111111011011001101)  
) LUT6_546 (
   .O(gates_283),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0011111101111110010001110001111110110111001100110010100011000011)  
) LUT6_547 (
   .O(gates_785),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b0011110100111111011000000011100001010011000010011101110110000111)  
) LUT6_548 (
   .O(gates_792),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0000010111110111100111010000111101111111001111001000000001100000)  
) LUT6_549 (
   .O(gates_1074),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1111111101011001110100111111010100000111001011001000001001001110)  
) LUT6_550 (
   .O(gates_1117),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1111100111010111100000000011000010110100011111101000101101111011)  
) LUT6_551 (
   .O(gates_1486),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0011001010100110100100000010110000011011111110001100100110001101)  
) LUT6_552 (
   .O(gates_1065),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1000101000101111111000110010010001001111011010111111001101011011)  
) LUT6_553 (
   .O(gates_1292),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1011000010110111100010110000110011001111010000110110110001100000)  
) LUT6_554 (
   .O(gates_402),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001010100100010111000001000110101111101000101111111111000101110)  
) LUT6_555 (
   .O(gates_1135),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0100001100010111010101000000100110010101110111101111111110000111)  
) LUT6_556 (
   .O(gates_1121),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1111101001110110101100100111111111010101111011111000001100100100)  
) LUT6_557 (
   .O(gates_879),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0011110101000010101111111000001000111000110101010000110001010001)  
) LUT6_558 (
   .O(gates_340),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0101010101100010001111010001101110100100110101101110101010100010)  
) LUT6_559 (
   .O(gates_510),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1111111111000000000000001100100110000100011001101001100011000111)  
) LUT6_560 (
   .O(gates_1080),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b1111010001001100001001111100010000111000101000000001100101111011)  
) LUT6_561 (
   .O(gates_417),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0101111011101011010000010100001000101001001101001111010100100011)  
) LUT6_562 (
   .O(gates_472),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0010001010001100010101011100100001111111101100110111110011110111)  
) LUT6_563 (
   .O(gates_200),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0101001110101110100111000111101000100101001001001011110010000101)  
) LUT6_564 (
   .O(gates_346),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1010011110101000111010010001010011110101101100011110000000010011)  
) LUT6_565 (
   .O(gates_553),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1011100110001111011010001011001110001101011101010010100010010010)  
) LUT6_566 (
   .O(gates_1180),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1100110001011000001111001110011100110101010111000010101000011000)  
) LUT6_567 (
   .O(gates_486),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1111100110001011110100000110011011010001100000010010011000100101)  
) LUT6_568 (
   .O(gates_686),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0110101110010001110110001111111011111011010111100000011110110000)  
) LUT6_569 (
   .O(gates_1084),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1101111011010001001010110011101100110011010101010000000000111100)  
) LUT6_570 (
   .O(gates_564),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0110101110110000110001100101011101001111100000101101100101100100)  
) LUT6_571 (
   .O(gates_719),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1100010000101100110101000110001110000100011110101011101010100010)  
) LUT6_572 (
   .O(gates_632),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b0111111000010101001110011100000001100111000111110110111110111100)  
) LUT6_573 (
   .O(gates_1390),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1000100011110111110001010011001111011011110110111101011000101010)  
) LUT6_574 (
   .O(gates_1285),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1111111000111010100000010111101101110010001010001101101100011010)  
) LUT6_575 (
   .O(gates_435),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1010111100110011100010000011010011001101101101100101101100100010)  
) LUT6_576 (
   .O(gates_1537),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1110011111101010011010011000110101001110011110000010011110110101)  
) LUT6_577 (
   .O(gates_80),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1101011111111110100101011001100110101011000000111111010111000110)  
) LUT6_578 (
   .O(gates_812),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1110010001010100011111010011110010000011101101000100010100100110)  
) LUT6_579 (
   .O(gates_824),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0111001101111111010101101111001100110101110100001110101010010100)  
) LUT6_580 (
   .O(gates_866),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1100100111010011001000100001101000011101001001000100111110101010)  
) LUT6_581 (
   .O(gates_1413),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0110011011011000001000111110001000011111000010101000011000011011)  
) LUT6_582 (
   .O(gates_1529),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1011001101010011011111011010100110100001000101100011001000011000)  
) LUT6_583 (
   .O(gates_221),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1101101111111011010001011001011011010100100111100110111110100100)  
) LUT6_584 (
   .O(gates_883),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0010011100011000010000011001110010011101101011100000111111001001)  
) LUT6_585 (
   .O(gates_74),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0011010011000110011011110011001111000000101001010110000000100001)  
) LUT6_586 (
   .O(gates_155),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0000100010001010010101111100110101100110001001011101100110000110)  
) LUT6_587 (
   .O(gates_266),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b1101111000001011001100011110001100110110111010100100010100111011)  
) LUT6_588 (
   .O(gates_1247),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0101110001110010011100000011111111000110000000000000010110000100)  
) LUT6_589 (
   .O(gates_438),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0011100111111110100001011011000001010000100110101101110111100000)  
) LUT6_590 (
   .O(gates_782),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0011100000110101001001010011101110101101000000000010110010000010)  
) LUT6_591 (
   .O(gates_1118),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0101000110001010011101011100110111001001010111010110101111000010)  
) LUT6_592 (
   .O(gates_589),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0000100110111001011100000100000110011010110010011010111101100101)  
) LUT6_593 (
   .O(gates_278),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0100100111100000011101001110001110000010101110110011110111111100)  
) LUT6_594 (
   .O(gates_1310),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0110011110101100010011000100101100001110010000010001111011111110)  
) LUT6_595 (
   .O(gates_882),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0111010110001111011111110101100011000001011111100001000101101000)  
) LUT6_596 (
   .O(gates_985),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1011101010101000100100011000111110011000010100010000101100111100)  
) LUT6_597 (
   .O(gates_684),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0011100011111001100000001001011000100101011101010111011101101110)  
) LUT6_598 (
   .O(gates_1131),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b1011111101001100111111110100001101101011101011001001011011010110)  
) LUT6_599 (
   .O(gates_25),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b1011001001000010010101100010100000001010110111011100101101000000)  
) LUT6_600 (
   .O(gates_89),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1111111011010011100110000100001101101011100000010100000010000111)  
) LUT6_601 (
   .O(gates_199),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1100111100100001101011010010011101011110011111111100110110000001)  
) LUT6_602 (
   .O(gates_669),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0100111110000101011100110000100000100110100011110000000100001100)  
) LUT6_603 (
   .O(gates_465),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1111100001011001110011110111101110111001000011110010010111000000)  
) LUT6_604 (
   .O(gates_171),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0000110001010000000110000001101100100010110101001101011110100000)  
) LUT6_605 (
   .O(gates_295),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0010111001010110101011010000100000110100111000100011100000000110)  
) LUT6_606 (
   .O(gates_136),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1000010101110100101011110011110110100110001011000000010101010111)  
) LUT6_607 (
   .O(gates_698),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0111001111110111010010001111001011011001000100110011010101010001)  
) LUT6_608 (
   .O(gates_1000),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0110101111001100010011001110111111011100000110010100111011100101)  
) LUT6_609 (
   .O(gates_1369),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1011100100001011110000010001101100000001001101101001110110110111)  
) LUT6_610 (
   .O(gates_204),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0000100000010100100011001011101010111111010111111011010100100111)  
) LUT6_611 (
   .O(gates_10),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1010000011001110101001111000011000001100001000100010011011000101)  
) LUT6_612 (
   .O(gates_840),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1110011110000100010110100001001101000110110100011000110010111100)  
) LUT6_613 (
   .O(gates_1002),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0001110110101001111100111101110111111001001110101011110110000011)  
) LUT6_614 (
   .O(gates_1342),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0000110000001110010101100101111000000001100011001110001000001010)  
) LUT6_615 (
   .O(gates_1323),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0011100011110101100101011101111100001011110011111000111100101010)  
) LUT6_616 (
   .O(gates_781),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0100101110110001001011110111101101101011111010010000010101100010)  
) LUT6_617 (
   .O(gates_723),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1101111110101000101010111010110111101011100111011101110111100111)  
) LUT6_618 (
   .O(gates_1139),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b1001100001111011100010110001000001100000011100101111011100000111)  
) LUT6_619 (
   .O(gates_578),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0100011010010110010110111000000001100100000010010101000100001101)  
) LUT6_620 (
   .O(gates_1308),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1100100000111001000100111100010011001011010100100001111001110100)  
) LUT6_621 (
   .O(gates_365),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1110011001010010010010011010100001010001110110111010100001000100)  
) LUT6_622 (
   .O(gates_814),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1110000101111110010010110111111110000101011111101011001110111001)  
) LUT6_623 (
   .O(gates_885),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0110110111110110010101110000110010010000010000110100001100101101)  
) LUT6_624 (
   .O(gates_370),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0000111101110100001010110001111001011010000111001100111011101100)  
) LUT6_625 (
   .O(gates_1076),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1001001010100001011101101111001100001011101000101110000101101100)  
) LUT6_626 (
   .O(gates_1260),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0001011010011001011010001110111010110110001101011101001101100011)  
) LUT6_627 (
   .O(gates_1188),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0010010010000000111011011011010010110010110100001101100010010100)  
) LUT6_628 (
   .O(gates_855),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b0000100110010011110010101001100111010101101000111111001111010010)  
) LUT6_629 (
   .O(gates_281),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1101100001101101101011001000001111100011111101000010000101100000)  
) LUT6_630 (
   .O(gates_157),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1000000000000001000111101011010011101001011001001110110001001110)  
) LUT6_631 (
   .O(gates_870),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0010000010100000010101001011000010000011010101011111111000010010)  
) LUT6_632 (
   .O(gates_144),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1110000100011111101001001010010101010010101111000110111111010110)  
) LUT6_633 (
   .O(gates_249),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1011101000101000011111011011110001001000011111011001110010011111)  
) LUT6_634 (
   .O(gates_436),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0010001010000100010010010110110000110010000010000111010111111000)  
) LUT6_635 (
   .O(gates_744),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0011001001111011100100101011101110010100011010100111101000001001)  
) LUT6_636 (
   .O(gates_1458),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0011100010010100001010001111111111110001010010010100000110111101)  
) LUT6_637 (
   .O(gates_1543),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0001100110111000000110010001011001100111000010001011001001111100)  
) LUT6_638 (
   .O(gates_268),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0101011101101011111001110011101111001000010011101001000110010100)  
) LUT6_639 (
   .O(gates_635),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b1101011110101110001110001110000001011000101100010011111011111101)  
) LUT6_640 (
   .O(gates_1028),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b1111010001000111010111111100000001110011010100101000001010111111)  
) LUT6_641 (
   .O(gates_1360),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0101101001001011001011010001110010110100000011010001111010001011)  
) LUT6_642 (
   .O(gates_822),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1001111111000111101010101001111100001001111001010101000011000111)  
) LUT6_643 (
   .O(gates_1006),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1100110010101001011100000001111001111101010111101001001011010010)  
) LUT6_644 (
   .O(gates_1303),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1011001010000010011000111010111000101101101010000000001101011011)  
) LUT6_645 (
   .O(gates_273),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0100110110011000111110010101101001101000101010011111000111110001)  
) LUT6_646 (
   .O(gates_55),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1000110101000111101000011111111001010101100100101001000101111110)  
) LUT6_647 (
   .O(gates_360),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0001101010110000111100110101000101000111100001010001001010010110)  
) LUT6_648 (
   .O(gates_205),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1000110011011010000000111100101001010101100100101010010100011111)  
) LUT6_649 (
   .O(gates_668),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1000111111011110000001111010100100111000110011010010101110010111)  
) LUT6_650 (
   .O(gates_997),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0110010001001101111001100110001110000011010011100010000010100101)  
) LUT6_651 (
   .O(gates_1383),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0100101100111011011001000110001000010101001111101011111111011000)  
) LUT6_652 (
   .O(gates_1346),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1100111100010101001110111001101001110010101110001111010110011101)  
) LUT6_653 (
   .O(gates_1025),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0010000101111000100101011010000101100001111000110001011111000010)  
) LUT6_654 (
   .O(gates_1036),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0011011011101100111110010101111101101010000011010011110001101110)  
) LUT6_655 (
   .O(gates_253),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0110000110111001011100010000011100111111011110010101000101101111)  
) LUT6_656 (
   .O(gates_1271),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b1011001110111101001010000000111000011110110011011001110000011011)  
) LUT6_657 (
   .O(gates_1142),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1010011100011111111010101111101001110100100000111101101110100111)  
) LUT6_658 (
   .O(gates_494),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1011100100110011001010111010111001110111110100110111110101001001)  
) LUT6_659 (
   .O(gates_482),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0101011100010110101010001100111011100100110001101000110001110111)  
) LUT6_660 (
   .O(gates_349),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0101111000000111101110101011011100101000011000001111001111011000)  
) LUT6_661 (
   .O(gates_1274),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0100000001011100110011100011000100010110101101010001010010110100)  
) LUT6_662 (
   .O(gates_716),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1110101100100110111000010010010101101010111010110000000101000110)  
) LUT6_663 (
   .O(gates_206),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0010111101000000000101001001101111001000001011001101010101000100)  
) LUT6_664 (
   .O(gates_109),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1001100011111000010010000000010100101100010101100101111010000111)  
) LUT6_665 (
   .O(gates_1061),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0001000111101000001001011010111010100101111101000011010100000010)  
) LUT6_666 (
   .O(gates_821),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0100000010011110011101001101111000111100111011100110100011111111)  
) LUT6_667 (
   .O(gates_383),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1110111010100101011001101100111011101011001111001010000110010100)  
) LUT6_668 (
   .O(gates_1195),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1000011011011100111100011110000001111110011110011010000010111110)  
) LUT6_669 (
   .O(gates_1454),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0110011111010101100100011010110010001010011010001001110000110101)  
) LUT6_670 (
   .O(gates_787),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0110001011101100000001010101101010110100011001111011011111100110)  
) LUT6_671 (
   .O(gates_696),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0001001100001100010110110101110010111110000110111000000101111010)  
) LUT6_672 (
   .O(gates_88),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1110001011000001101010001001011100111101000101101111101101000000)  
) LUT6_673 (
   .O(gates_876),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1111011100010010100010110010111111111100111010011010010111010000)  
) LUT6_674 (
   .O(gates_994),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1001111110111000100110010011110010001101011100010111011000100011)  
) LUT6_675 (
   .O(gates_192),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0000010100111001010001100110010111000000000001110101110111111011)  
) LUT6_676 (
   .O(gates_1011),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0001000001010111100100011101011111011100011011101100001101111100)  
) LUT6_677 (
   .O(gates_111),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1110101111011110001110110110101011000010001000001111100011101110)  
) LUT6_678 (
   .O(gates_458),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1101001000101111001010000010110001010001000011011100100000110111)  
) LUT6_679 (
   .O(gates_286),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0101100001101000011110000110000101001011001001111000110000001100)  
) LUT6_680 (
   .O(gates_445),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1110001000011000100110010100110101100001100010000010010110101011)  
) LUT6_681 (
   .O(gates_1302),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0001100011011101100110111001000010000001100110000000100101100100)  
) LUT6_682 (
   .O(gates_924),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1110111001111111100010001100101000010011111111001001111111001111)  
) LUT6_683 (
   .O(gates_990),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0001010111011100110001010011010010100001011010001110100111101100)  
) LUT6_684 (
   .O(gates_689),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1101110101111101100000010001001010111110000111100011110000001100)  
) LUT6_685 (
   .O(gates_1114),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b1010011001001111100000010100100100111010000101101010000010100101)  
) LUT6_686 (
   .O(gates_376),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1001011101010010010101110111110010001000010001100000011101110000)  
) LUT6_687 (
   .O(gates_404),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1001010011101001110010001010001110111110000101110100101001100000)  
) LUT6_688 (
   .O(gates_1126),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0001101110100001110000110111101101010101010011010100100110011100)  
) LUT6_689 (
   .O(gates_863),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0011000101101011001000001001110100101101101111111110011000011010)  
) LUT6_690 (
   .O(gates_1174),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0110101000111010010000010011101010010111011101111110100001000000)  
) LUT6_691 (
   .O(gates_762),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1100001010101011101100011001011101011001000010110100110110111011)  
) LUT6_692 (
   .O(gates_852),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0111100101000000101010110010110011010010101101100111111000110110)  
) LUT6_693 (
   .O(gates_949),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0100000010111001011010100011000101001110111000101001001001000011)  
) LUT6_694 (
   .O(gates_1519),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0000111111001011010110001100010011010110000001100111000111110001)  
) LUT6_695 (
   .O(gates_905),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0101110001001011111111110011110110001000000001000101001000100011)  
) LUT6_696 (
   .O(gates_953),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0101110100010101111001001001000000011111000110100011000100110101)  
) LUT6_697 (
   .O(gates_1229),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1001001011000110011111011001101001111011101100111011111001000101)  
) LUT6_698 (
   .O(gates_508),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1101001111101101001101001000001111001110010011000011111011110101)  
) LUT6_699 (
   .O(gates_310),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1000000011000000001111110001111100100000100110100101001011100100)  
) LUT6_700 (
   .O(gates_572),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1111100110110010000010011001100010011000010000110101010010001010)  
) LUT6_701 (
   .O(gates_481),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0011010000001001110000011110011111010101101001111001110010100010)  
) LUT6_702 (
   .O(gates_333),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1111111010010111000101110110110000011000111101011110010100110100)  
) LUT6_703 (
   .O(gates_1191),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0101001001011011001000110111101000111001101011000001101101011000)  
) LUT6_704 (
   .O(gates_148),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1101100001011000011010001111001101100101110111101011110100101111)  
) LUT6_705 (
   .O(gates_1394),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1100101001000010011100111110011101101011101011111000010110001011)  
) LUT6_706 (
   .O(gates_186),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0111010111001110101110010111100110101010010011110100001001100001)  
) LUT6_707 (
   .O(gates_418),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1110010001100101100010111011111111011010011010100111100111000011)  
) LUT6_708 (
   .O(gates_478),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1000011110011110011101000101111110000111000000101101101011101100)  
) LUT6_709 (
   .O(gates_1094),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0000101111001001110111010000110110011010110001000111011011110111)  
) LUT6_710 (
   .O(gates_931),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1100001001100101010100111111001110000110001101111111011001100111)  
) LUT6_711 (
   .O(gates_991),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0010010001001000110100101100100001110101001110101000000011011111)  
) LUT6_712 (
   .O(gates_1450),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0001100101100101111111011101101000010111100100100100011101110011)  
) LUT6_713 (
   .O(gates_434),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1110101011010010111101111110000110010001111101110011110101111011)  
) LUT6_714 (
   .O(gates_1419),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0110110101101001101011011001110000000110001001011010010000110111)  
) LUT6_715 (
   .O(gates_382),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1100001011011000100110011100011001010000000100111111000010101100)  
) LUT6_716 (
   .O(gates_1465),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0011001001100001100110100110101010011100110011001100011011010010)  
) LUT6_717 (
   .O(gates_127),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0110111100000101111001010111000100101100101100110001111100111000)  
) LUT6_718 (
   .O(gates_783),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1101001011111101000101010101000110111011110110111111100001100011)  
) LUT6_719 (
   .O(gates_187),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0011111111000100001001100000110011101111000111101100101010001111)  
) LUT6_720 (
   .O(gates_1034),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0101010001101110101000010000110111000011010010001100010111111011)  
) LUT6_721 (
   .O(gates_36),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1101011010111000010111100011000011011011010010110100001010101101)  
) LUT6_722 (
   .O(gates_913),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b0000010100000001100100100000111110110100100100100101010111011111)  
) LUT6_723 (
   .O(gates_416),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1001001001110011011011000110101111111101011110010101000011001001)  
) LUT6_724 (
   .O(gates_1270),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b0111101011011001000111001101010110001101110000011111010001111111)  
) LUT6_725 (
   .O(gates_904),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0011111111111101100111000110011100011000100101100011000110100001)  
) LUT6_726 (
   .O(gates_339),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0010000111111100011100010011100010010111100011001111011001000011)  
) LUT6_727 (
   .O(gates_535),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1101110111011111000100110000101100110011000100001001101100011000)  
) LUT6_728 (
   .O(gates_1123),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1100001011001111110101100011000010110111111110001111001001001110)  
) LUT6_729 (
   .O(gates_881),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1111100100000010110001010111000000111111000011100001010011110010)  
) LUT6_730 (
   .O(gates_1279),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0010010001000011100011100100010010011100000111111010110010110001)  
) LUT6_731 (
   .O(gates_631),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1010110000111101001100100111010110010101010000001101001101101100)  
) LUT6_732 (
   .O(gates_692),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b1100100010000111000100000111101111011001010000100010111011001100)  
) LUT6_733 (
   .O(gates_1259),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1100000001000001001010011111110110110100110100100010100011011001)  
) LUT6_734 (
   .O(gates_880),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0001011100010101010101110101000100101010110010101000110110010111)  
) LUT6_735 (
   .O(gates_550),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0101010011010110001010111100011101000011011100110110100011001010)  
) LUT6_736 (
   .O(gates_1492),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0000110001001111000101011011110111110001011011111000101001110001)  
) LUT6_737 (
   .O(gates_67),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1010111001011100001101011111100111001001111000011010101011000101)  
) LUT6_738 (
   .O(gates_1250),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1110000111000000001001101100011111101111001110101010110111001011)  
) LUT6_739 (
   .O(gates_135),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1001110101010000011101101000110100101000010100100110000110111101)  
) LUT6_740 (
   .O(gates_108),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0001111101000010000000000100010110111000001011011011001101100010)  
) LUT6_741 (
   .O(gates_178),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1110110010101110110110011010000000011000011001000011001100101100)  
) LUT6_742 (
   .O(gates_1338),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0101010101110010010010000001010001000001101011010111100100101010)  
) LUT6_743 (
   .O(gates_623),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b1011010001011101000110100001111110111000011111111110101001001111)  
) LUT6_744 (
   .O(gates_230),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1110110111010010101100010110101010111011101011110011011111100110)  
) LUT6_745 (
   .O(gates_440),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0001000110100110100110110100010111100011100100011101111110100001)  
) LUT6_746 (
   .O(gates_604),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0010100011000010100010010001011101110000101011001101100111111001)  
) LUT6_747 (
   .O(gates_1471),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0011011010000011101101101001001100010110101000110111101011100101)  
) LUT6_748 (
   .O(gates_743),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1010101010110001110001101101011111010100110000011000000100011101)  
) LUT6_749 (
   .O(gates_1019),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b1001101010111010011110011001001010011111010011001100111011011010)  
) LUT6_750 (
   .O(gates_220),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b1110111111001000011010110100001111001111101111000010101110001100)  
) LUT6_751 (
   .O(gates_484),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1000000011100000011111100100010011000110100100010001000110001001)  
) LUT6_752 (
   .O(gates_391),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0110010011111100100010001100011101000000110000001101101001001101)  
) LUT6_753 (
   .O(gates_1212),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0000001011010010010000100110111100001111001000000001010000111011)  
) LUT6_754 (
   .O(gates_1509),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0011110001101100000110110110000010111110101111010001001010011110)  
) LUT6_755 (
   .O(gates_749),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0111000101111011110001100011101011101001101010010110011001101000)  
) LUT6_756 (
   .O(gates_342),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1101111010101000001111001111001110111001111100001001001000111111)  
) LUT6_757 (
   .O(gates_942),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1010010100111111100000101100110111100100010000011110110100010011)  
) LUT6_758 (
   .O(gates_189),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b0100010100011100001011101101000101100110010111001111000011100011)  
) LUT6_759 (
   .O(gates_92),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0111000111100101000110111100111110111111100111101101110001000010)  
) LUT6_760 (
   .O(gates_1045),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0000001111011001111101001001101001010000100011001000111001110111)  
) LUT6_761 (
   .O(gates_45),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1111000000000111111001010111000001000001010101001101011110000000)  
) LUT6_762 (
   .O(gates_738),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0101011110001101100011111101100001110100111010111111010010011100)  
) LUT6_763 (
   .O(gates_562),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1000101001110110001010100100000111010110110010101111000111001011)  
) LUT6_764 (
   .O(gates_1181),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1100000100010111001011000100010011110101111001010001011011001111)  
) LUT6_765 (
   .O(gates_1046),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1010100100010001110010010000100111101011010110110110010011111011)  
) LUT6_766 (
   .O(gates_1200),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0001100111001001110110110001101010001100111111111101101110111100)  
) LUT6_767 (
   .O(gates_1112),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1101011110010011100010010000101110011110100101010011101011110110)  
) LUT6_768 (
   .O(gates_955),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1011110111111010001111101111110110111000111111100101110110101111)  
) LUT6_769 (
   .O(gates_1102),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0001000000111001101111111010010000010011110101110111100110110111)  
) LUT6_770 (
   .O(gates_369),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0110101000100001011110001000110001011010010010000101011100000110)  
) LUT6_771 (
   .O(gates_661),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0110111101110101010001011111001101101110011001001100011100110000)  
) LUT6_772 (
   .O(gates_556),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0011001010011110110110111010000010110001011011100111000101101111)  
) LUT6_773 (
   .O(gates_509),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1100111111101101110001111111000110100001101000010010011000010001)  
) LUT6_774 (
   .O(gates_245),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1001101101001111100010111110111000000100101001100110010101000001)  
) LUT6_775 (
   .O(gates_1505),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1100000001000010111000100000111110000001000010010010100010111001)  
) LUT6_776 (
   .O(gates_311),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0001010011001011110111111100000000011101100011001100111100010001)  
) LUT6_777 (
   .O(gates_984),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1000100101001100011110010001000011101111100110011010001010101011)  
) LUT6_778 (
   .O(gates_137),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1100101110100101111110100111110010010110010010000101100100111100)  
) LUT6_779 (
   .O(gates_454),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0010101110100100011100111110111100011001101001011110100000001110)  
) LUT6_780 (
   .O(gates_375),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1110011111100010000101011100001110101101001101010011000010101010)  
) LUT6_781 (
   .O(gates_1460),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b1000101011010001101101011000111111010001100011001010000110110011)  
) LUT6_782 (
   .O(gates_1157),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0101100001100000101010111100100000111110000000000111110001001011)  
) LUT6_783 (
   .O(gates_1258),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0110000000100001000101101101101011010100101010111001010101010101)  
) LUT6_784 (
   .O(gates_1502),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0110010001100100010100011100110111001111000001000111101001100100)  
) LUT6_785 (
   .O(gates_611),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0000010000100010111000001111000111000101010111000111100110100011)  
) LUT6_786 (
   .O(gates_76),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0101111000101000000001011011100000110100011011011111101010101100)  
) LUT6_787 (
   .O(gates_715),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1111111010110011101110010010101110000001101111010101100110000101)  
) LUT6_788 (
   .O(gates_1374),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0010011000110111110001010010111111110000110100111100100111001011)  
) LUT6_789 (
   .O(gates_1462),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0010000000011111001100101000111000101001000000000001011111010001)  
) LUT6_790 (
   .O(gates_888),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0011011001100000101110010111100010100101010000011011111111110110)  
) LUT6_791 (
   .O(gates_1073),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0011011000100111100111010101110011001110101111011011010101001110)  
) LUT6_792 (
   .O(gates_1358),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0101001010000110010001010011101011110000001111011100110101111111)  
) LUT6_793 (
   .O(gates_1218),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0110000100011111110100111011111110001000011001011000011000000001)  
) LUT6_794 (
   .O(gates_119),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0100011101001110111010111111011110100001100111011010111000001001)  
) LUT6_795 (
   .O(gates_1410),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b0011111011100110101011011011111010111111110111110111110001010111)  
) LUT6_796 (
   .O(gates_1205),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0010010001001011101111011100010001000001010000000010111010011100)  
) LUT6_797 (
   .O(gates_588),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0110111101011111011100010100111110100000001000110000001001001000)  
) LUT6_798 (
   .O(gates_32),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0001011001110100000010010000001000101110111101100110010110101100)  
) LUT6_799 (
   .O(gates_796),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0000001100101001111101100010111011100010111001111101010111100100)  
) LUT6_800 (
   .O(gates_198),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1011000110100111100100111111000001110011110101000111100110101110)  
) LUT6_801 (
   .O(gates_1232),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1010011000011100010110110110110100011001011110001011010111000100)  
) LUT6_802 (
   .O(gates_773),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0011001000001010011100011100000110010000111010100000001110011001)  
) LUT6_803 (
   .O(gates_31),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0101110011110101001110010100010101001111010011010110011001001010)  
) LUT6_804 (
   .O(gates_672),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1010001000100111011100100110101000001110111101000001011011001110)  
) LUT6_805 (
   .O(gates_1111),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0110101010111111010011010011110001100011100100101011000000110111)  
) LUT6_806 (
   .O(gates_844),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1010010001010100000110100100001011000000110011111010010000110000)  
) LUT6_807 (
   .O(gates_901),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0001111100100001001101111010010110011110001100110010110001001101)  
) LUT6_808 (
   .O(gates_833),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1110010010010001010110010110110101110010100000000111000111100001)  
) LUT6_809 (
   .O(gates_1349),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010010000011001111111111101011001101101001100101111111011000100)  
) LUT6_810 (
   .O(gates_1525),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0100101101101011100111101100011000010000111101000111111001100001)  
) LUT6_811 (
   .O(gates_363),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0010111110110011110001000110000101110011101000111110010001000011)  
) LUT6_812 (
   .O(gates_618),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1000011110010011100101111001000100110111011110101111111100110001)  
) LUT6_813 (
   .O(gates_644),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0111000000001010111111111110110101010000011001101111001001101001)  
) LUT6_814 (
   .O(gates_519),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1100111101100010100000111000011110001000010000010110101100111011)  
) LUT6_815 (
   .O(gates_1442),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0001101011001110000101010011111000101110001000010101110010110011)  
) LUT6_816 (
   .O(gates_854),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1101000011001011111101101010111111011010111001100010011010111111)  
) LUT6_817 (
   .O(gates_44),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1101101000001100011100101010011010000000000100001011110110011000)  
) LUT6_818 (
   .O(gates_1096),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1011010000100111111100101111011011001000110101110000101111011101)  
) LUT6_819 (
   .O(gates_471),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0011110100111110000111101101110101000110001110100011110010100011)  
) LUT6_820 (
   .O(gates_769),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1100010000000111000011111110111101111100000010110000110110011110)  
) LUT6_821 (
   .O(gates_853),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0111111011111001111010000110000101101010111101010001000001111100)  
) LUT6_822 (
   .O(gates_241),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1011110100110001101110001000011101111011011110101101001101000101)  
) LUT6_823 (
   .O(gates_1185),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1001011001110010000010101010110011110000011111010011100001010111)  
) LUT6_824 (
   .O(gates_1313),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1111100111100001100111111101010111011011000011111111010001000001)  
) LUT6_825 (
   .O(gates_1007),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1011000000001111100001111110101101001100011011001001001111010010)  
) LUT6_826 (
   .O(gates_603),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0110010000000111101101000101101001000000010100110010011101110101)  
) LUT6_827 (
   .O(gates_1138),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1011100010011101111011001011010100111100011000111001010111000100)  
) LUT6_828 (
   .O(gates_849),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b1110010100101010110010011100011010010111100001100000110001010011)  
) LUT6_829 (
   .O(gates_280),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1000110001100010111111111111111001100011100010100011001001001001)  
) LUT6_830 (
   .O(gates_660),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0101100001000000010011010010111010010110111111110101000100010010)  
) LUT6_831 (
   .O(gates_1514),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0001001011101011100001101111001110111010101011111100001100101101)  
) LUT6_832 (
   .O(gates_1035),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b1001101100100111111001000001111011000000011000000010011001011011)  
) LUT6_833 (
   .O(gates_934),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1110001100110100011110011011100100011000000010001010010000001101)  
) LUT6_834 (
   .O(gates_602),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0010000111100100100001000001110001000110100010000111100100010000)  
) LUT6_835 (
   .O(gates_1377),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b0000011101010101111011100000000000001111011101100000100000101100)  
) LUT6_836 (
   .O(gates_298),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0110100011100100101010100011110011000111100000100111001101101011)  
) LUT6_837 (
   .O(gates_643),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1001111011011000100000010000001001100010011111100110100101000101)  
) LUT6_838 (
   .O(gates_1475),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1010101101000100011110110001110110100101110110100110010000111111)  
) LUT6_839 (
   .O(gates_164),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b1001111001011110110000010100010011100110011100100010110010011100)  
) LUT6_840 (
   .O(gates_190),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000011111110000010001011010001011001011110000100100000000111011)  
) LUT6_841 (
   .O(gates_1467),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1000011001101010111011011011111010101001100010111111100011000000)  
) LUT6_842 (
   .O(gates_605),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0011100111100111010100100110110001110111001101100000111110000111)  
) LUT6_843 (
   .O(gates_706),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1101001001100001110001100110110110110100110001010011001100111100)  
) LUT6_844 (
   .O(gates_1203),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1001010111010011101100100000000110000111101001111101110000110011)  
) LUT6_845 (
   .O(gates_1249),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0010001001001000100100010010111111011110100100111101011100001101)  
) LUT6_846 (
   .O(gates_579),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b1110001110011010100000101011100011111101111110011101110011011010)  
) LUT6_847 (
   .O(gates_343),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1001011000111110001001111001010000010100011010100110100010110111)  
) LUT6_848 (
   .O(gates_1058),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0100101101010110101111111100000001001110011100000101000110100110)  
) LUT6_849 (
   .O(gates_1380),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1001101111111001011010100101100101001110010110000000001101000000)  
) LUT6_850 (
   .O(gates_21),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1001110000000110010001101000110110011001011000110011000010111010)  
) LUT6_851 (
   .O(gates_810),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b1111110111110010110110111100100101000001000001010111011100101001)  
) LUT6_852 (
   .O(gates_1451),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0011010110000100010000101000101101111101001001001000100110101111)  
) LUT6_853 (
   .O(gates_52),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0011000010001010010011100010110100100111011101010110010010100010)  
) LUT6_854 (
   .O(gates_575),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b0100100001111100110011111000110000110001001100001001101010101110)  
) LUT6_855 (
   .O(gates_226),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1010101111011101111011001100000001110110011011111001011101110110)  
) LUT6_856 (
   .O(gates_986),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0110000000101101101100111101111100100111100101100011010101010011)  
) LUT6_857 (
   .O(gates_1105),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0110011110000001111000010000000001000111111110110011100000111111)  
) LUT6_858 (
   .O(gates_583),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0010000011100111101111001111111101100111110010001101101111111001)  
) LUT6_859 (
   .O(gates_98),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1000100000011010101110111010111111110111010010001100101000111111)  
) LUT6_860 (
   .O(gates_1407),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1001111000101001100000011111001000100100000111011100010000100100)  
) LUT6_861 (
   .O(gates_693),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0100011000101001100110111101101010101100111101011001101110000011)  
) LUT6_862 (
   .O(gates_258),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1110000101001000000101111101010110010110100111110111001100001011)  
) LUT6_863 (
   .O(gates_48),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0010101100011110011100000011001101000110111010101101100000010000)  
) LUT6_864 (
   .O(gates_1087),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1111001101011111110000110011011010001011011010111010100001011001)  
) LUT6_865 (
   .O(gates_1345),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1101100000010100010000111100110111010000100011111010000100010111)  
) LUT6_866 (
   .O(gates_20),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1010110111010010100100000111010001010100001001111110111011111111)  
) LUT6_867 (
   .O(gates_915),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0001101010101100011001010010001001010010000000000100011010001000)  
) LUT6_868 (
   .O(gates_322),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1010101001101110100001011101001010001000110111110111010110100100)  
) LUT6_869 (
   .O(gates_750),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0010001001101100110001111011101101101101000000000111011110010001)  
) LUT6_870 (
   .O(gates_211),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1110011011000101000111101000110111111101000110100011011100111001)  
) LUT6_871 (
   .O(gates_1207),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1110001100011010111101011010111101000110000101111010101001010100)  
) LUT6_872 (
   .O(gates_246),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1001110100011101000111111010101011001110000101010110111010101100)  
) LUT6_873 (
   .O(gates_276),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0110110100000000111100010100010010101001000101110111011001100001)  
) LUT6_874 (
   .O(gates_304),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b1000111101010010101011011110000101010011000011111111011011110010)  
) LUT6_875 (
   .O(gates_1083),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0101100010000001011001110110011000111000000111101000110100100110)  
) LUT6_876 (
   .O(gates_502),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0010011101111111100101000111001010110011111011001010000110100101)  
) LUT6_877 (
   .O(gates_409),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0001010010100111001100111111100000010011000101101101111011010011)  
) LUT6_878 (
   .O(gates_1213),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1101011110110100101010001101101010111011110011011000001100001111)  
) LUT6_879 (
   .O(gates_290),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0110010000000110111010010110011100110101011101100110110100000010)  
) LUT6_880 (
   .O(gates_1068),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0100100110011011100100001110000111100001111000010111111101101010)  
) LUT6_881 (
   .O(gates_85),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1010111111111110101011000011111111000110010001011000101011011010)  
) LUT6_882 (
   .O(gates_170),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1110101000010101111101011111111011000101001101010000100111100001)  
) LUT6_883 (
   .O(gates_1535),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0110000010111010001101011110101010011000100001111000001110000010)  
) LUT6_884 (
   .O(gates_664),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0100111010000000110101110100001000010111011100111001011011011100)  
) LUT6_885 (
   .O(gates_86),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1001110011011010010000101110110101101111100110001101001100001010)  
) LUT6_886 (
   .O(gates_26),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0010010011111110010000110110110001001101111011100001001001010100)  
) LUT6_887 (
   .O(gates_981),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b1101110110111001101111000101100010000000100110111000000000011010)  
) LUT6_888 (
   .O(gates_338),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1111100101000111011010110011000110101101100100010001110000001001)  
) LUT6_889 (
   .O(gates_351),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0011010001011100011111110101110100001101111111111001110111010010)  
) LUT6_890 (
   .O(gates_22),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1010101000111001011000000111000100001100001010111011101111000110)  
) LUT6_891 (
   .O(gates_1269),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1001111011000100010111001000011110101100100100111011001000111100)  
) LUT6_892 (
   .O(gates_1457),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1000111100101000111101001101011001011010001001001010110101111000)  
) LUT6_893 (
   .O(gates_1405),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1001011101100111100101010011110000101100011100001010010100110011)  
) LUT6_894 (
   .O(gates_1359),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0111110101101000101000011000010010101110101100111011010100011010)  
) LUT6_895 (
   .O(gates_832),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1110000000100010110011001101010110101001010101101000010001011000)  
) LUT6_896 (
   .O(gates_1266),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0000101010011000111101100011100101010010100111001111100111111001)  
) LUT6_897 (
   .O(gates_1165),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1111110100001010110010110000111000010010110100100000010101110111)  
) LUT6_898 (
   .O(gates_974),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0101011011111101011000010001010101111111011100101101011001001011)  
) LUT6_899 (
   .O(gates_1275),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1011001000101001011001000010101111011101100100101101101011001001)  
) LUT6_900 (
   .O(gates_1403),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1010100110001010010001010011011111010101100100000011110001101100)  
) LUT6_901 (
   .O(gates_1538),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0001110000111100100010011101100110111110101011010001110011000101)  
) LUT6_902 (
   .O(gates_81),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0001011010100000111101000010010010101010010000110011100101111011)  
) LUT6_903 (
   .O(gates_134),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1010110100101011100111010110000111110110001100110000001000001100)  
) LUT6_904 (
   .O(gates_702),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1011111001111010100101110101010010110111001110101010110001110110)  
) LUT6_905 (
   .O(gates_705),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1000001010000010101000111010101000100101000001110101001000100010)  
) LUT6_906 (
   .O(gates_1402),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b1001110000100010100101010010010001110110001101010011111001100001)  
) LUT6_907 (
   .O(gates_515),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0110111101001010100111000101011001101011110111110110100101110101)  
) LUT6_908 (
   .O(gates_384),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0110110000111110011110100100010001000000110000110000101000000000)  
) LUT6_909 (
   .O(gates_884),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0111000010101010000111111001001101010101111000000110001011000011)  
) LUT6_910 (
   .O(gates_1017),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1111011101110101011111100000111100010110000010101110111001111110)  
) LUT6_911 (
   .O(gates_554),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0000110010010111100111110010001001111000000010011001100111000011)  
) LUT6_912 (
   .O(gates_951),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0001101001001011010101110110111101100111010010101110100100010111)  
) LUT6_913 (
   .O(gates_1319),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0111011000100110000001101111111100010000010011100011111010011110)  
) LUT6_914 (
   .O(gates_737),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1011000100001001000001100001111001001010011111101011110110011101)  
) LUT6_915 (
   .O(gates_573),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1111100000000010111110101101110101001000000101001001001010101101)  
) LUT6_916 (
   .O(gates_517),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1010111101000000010100011101000101011100011111000011001011110100)  
) LUT6_917 (
   .O(gates_1071),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0101101110111101100001000000001011111011001010111011011110000110)  
) LUT6_918 (
   .O(gates_24),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0011100010111110101111101100001110011110100011010101000110011111)  
) LUT6_919 (
   .O(gates_1376),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1100000100110011000001001001000100101101111001000110011110001110)  
) LUT6_920 (
   .O(gates_671),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1000001000000100110001011101011100010001100111000110000100111110)  
) LUT6_921 (
   .O(gates_39),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0010001011110110010101111110000100010010100010000010111000111000)  
) LUT6_922 (
   .O(gates_244),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1110000011000101101100110101011011110111000101110101111100101111)  
) LUT6_923 (
   .O(gates_1208),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0001111000101110110000001010000010011111100110100000011101000011)  
) LUT6_924 (
   .O(gates_12),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0010110100101010010110001010101110100010001110101010101110110010)  
) LUT6_925 (
   .O(gates_1520),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0010110100010001001110111110010011111000010100101011011100011010)  
) LUT6_926 (
   .O(gates_818),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0010100000000001011100011100001000100110111101100110010100000110)  
) LUT6_927 (
   .O(gates_759),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0110000001000100111000000000001111000011011100100111000110011001)  
) LUT6_928 (
   .O(gates_499),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0110110111001101101011111110110001101010111110110110010001000010)  
) LUT6_929 (
   .O(gates_83),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0011111101111111011000000101111101000000011100100101100011011110)  
) LUT6_930 (
   .O(gates_130),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0101111010010100110110010111001010101110100000001000000010001001)  
) LUT6_931 (
   .O(gates_1524),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1001110010110111011010010000111000101110001011000110011101011011)  
) LUT6_932 (
   .O(gates_496),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1001100111101100111000001010000101011000010010001001000101101010)  
) LUT6_933 (
   .O(gates_1494),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0010101110110000001000010000111101110010100101001001101110100100)  
) LUT6_934 (
   .O(gates_751),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0011001111100101100110110000000100011001001110011000011011011100)  
) LUT6_935 (
   .O(gates_505),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0011100100000101001001111011110110010100010101100110110010111001)  
) LUT6_936 (
   .O(gates_287),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0010111000111110000101101010000000101110001001001100001011001100)  
) LUT6_937 (
   .O(gates_662),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0111000110001101110101011111000101111001111100100001110000000001)  
) LUT6_938 (
   .O(gates_180),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0010001001011111011101000000000010001110001110111011010101100000)  
) LUT6_939 (
   .O(gates_1477),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0000011101101111011100110111110000011111101001000101000101101001)  
) LUT6_940 (
   .O(gates_1189),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1100110010110101101000110100101000101100100001011100100100100000)  
) LUT6_941 (
   .O(gates_305),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b1001000001110111001101010001101100001010110100101010111110000010)  
) LUT6_942 (
   .O(gates_1427),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0100001000111001001011000101000011011010010001111011101111100110)  
) LUT6_943 (
   .O(gates_355),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0001101110110110110000011111001011011001000010000100000001111001)  
) LUT6_944 (
   .O(gates_325),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b1101011011001010110110100110111000000000111110100110011001000110)  
) LUT6_945 (
   .O(gates_397),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1000000000110110011110110111101100011101001100101101110101000111)  
) LUT6_946 (
   .O(gates_282),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0001010010111110000111100001110111001101000110100100011011000000)  
) LUT6_947 (
   .O(gates_1554),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b1000010000011001100101111110001111111101101100100011111110000101)  
) LUT6_948 (
   .O(gates_168),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1001111111111100101001000010100111001110100001101100010011111011)  
) LUT6_949 (
   .O(gates_1322),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1000110100101000010011100000011010000001100100101111101100000011)  
) LUT6_950 (
   .O(gates_492),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1011000010010101101000011110011100100001010110100010010111010100)  
) LUT6_951 (
   .O(gates_940),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0111100101100000110010000001110100000001101111101001011010001111)  
) LUT6_952 (
   .O(gates_1432),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1101001001011011000101111010000001011100110100001100010011101100)  
) LUT6_953 (
   .O(gates_274),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1010001000111000111010010010101110110010101010011101010110110011)  
) LUT6_954 (
   .O(gates_1480),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0000010111001110011111111011000101001000110110011100111001010000)  
) LUT6_955 (
   .O(gates_889),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1110100001001110110011011000010011000110011111101011000010111101)  
) LUT6_956 (
   .O(gates_748),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1010000100110100011111000011101001001110001001101001001110100011)  
) LUT6_957 (
   .O(gates_758),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0011011000011010111010111010110111100000101100010110100111010111)  
) LUT6_958 (
   .O(gates_331),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0001101110101110000000000001001011011101100000100001111111110100)  
) LUT6_959 (
   .O(gates_1238),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1101100101011110001111101110000100101110101000000000011111001010)  
) LUT6_960 (
   .O(gates_957),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b0001110000000011000000001111111000101010011000011000010001000111)  
) LUT6_961 (
   .O(gates_965),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0011010111001101001110101101100101010111000111100001010011101011)  
) LUT6_962 (
   .O(gates_872),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0101100100001110001100000111001010001111111110111111111000011000)  
) LUT6_963 (
   .O(gates_566),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b0011100000001101100000000001011111110000100001010101000110001101)  
) LUT6_964 (
   .O(gates_1085),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0001000000110101101011110100110111000111110000100101111110011101)  
) LUT6_965 (
   .O(gates_1334),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1110010100010100101000111011010000001011001111110111000111001101)  
) LUT6_966 (
   .O(gates_191),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1110100111000011101100001010001000010100011111011101101011011011)  
) LUT6_967 (
   .O(gates_1192),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0011101111010001010111010111001010110110110111000101111001101100)  
) LUT6_968 (
   .O(gates_1399),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0100011100001100010111001111000000001100000000001100010010100000)  
) LUT6_969 (
   .O(gates_893),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0100110101100000001110010100100100000111101100011100110000100100)  
) LUT6_970 (
   .O(gates_626),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0000101100000000111101101110000011111001101001010011101010011010)  
) LUT6_971 (
   .O(gates_1173),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0111111010001011000011100110100110000000110010011000110001111011)  
) LUT6_972 (
   .O(gates_836),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0010000111101101110001010001010111001100001100111101100111010100)  
) LUT6_973 (
   .O(gates_798),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0011000001011111110100111110000110110011001110011100001010110100)  
) LUT6_974 (
   .O(gates_896),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0110100111011010011100000011100100101111101001100101100000111011)  
) LUT6_975 (
   .O(gates_584),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1110101000111000110100000100101101111111011010101110100001000001)  
) LUT6_976 (
   .O(gates_1532),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0101011011011001100100111101111100010010011111110000100011101000)  
) LUT6_977 (
   .O(gates_399),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1011000100101001010010011010011010100111001111000011100100010001)  
) LUT6_978 (
   .O(gates_413),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1111011101010000001000010101110100000010001101010001010110011001)  
) LUT6_979 (
   .O(gates_1443),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0001101010011111001111101011100111001100110001001000011000010011)  
) LUT6_980 (
   .O(gates_1081),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1001001000000100110101011001011100110111100111100011101111110100)  
) LUT6_981 (
   .O(gates_613),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1010101110101110001111101111011100010010000000100010011010001111)  
) LUT6_982 (
   .O(gates_1013),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0101101011000010110000100110010111101100000110001100010000001100)  
) LUT6_983 (
   .O(gates_16),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b1011110011010111101110111110101111111100110101010010111111100001)  
) LUT6_984 (
   .O(gates_1366),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0011001011011100001000110110010011100000001100011000101010010101)  
) LUT6_985 (
   .O(gates_862),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0010011010101110100110110000011011100011011100001101010101110111)  
) LUT6_986 (
   .O(gates_54),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0101110001110100111011110101001000111001001001000010000010000111)  
) LUT6_987 (
   .O(gates_1476),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1110000100011101110010001001000000111011011000001101010001010001)  
) LUT6_988 (
   .O(gates_691),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0111000001100111000000010101001010101111100000001000111101011010)  
) LUT6_989 (
   .O(gates_131),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1010001010000111010101000000001101010011011000101111101100001001)  
) LUT6_990 (
   .O(gates_890),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1001000001011000001010100110000110010110011110110011110111000101)  
) LUT6_991 (
   .O(gates_730),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1000111100111111000100110001011001000111100010010101001010000011)  
) LUT6_992 (
   .O(gates_944),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0111010100010001100110001000110001001100011101000111110111111101)  
) LUT6_993 (
   .O(gates_453),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0000011110000001110110100001101101101101010010101100100101100001)  
) LUT6_994 (
   .O(gates_1241),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0010110001100010101111010100000000000101001000010001001010001101)  
) LUT6_995 (
   .O(gates_1547),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1000111111001100111100000100110111010101111000111010010111110100)  
) LUT6_996 (
   .O(gates_777),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1100110101100101100110111101000101011000001110010100100001011010)  
) LUT6_997 (
   .O(gates_1040),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0000000110011111100011010110011100011111011111110111101010001011)  
) LUT6_998 (
   .O(gates_1456),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0001111000010010000100010010101110100100010000111111010100110011)  
) LUT6_999 (
   .O(gates_1305),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1110111001001011011100101101001100000110101011101001111001010111)  
) LUT6_1000 (
   .O(gates_920),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0001001100011001010100100000011111010111100100010111101000110011)  
) LUT6_1001 (
   .O(gates_523),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1111000000001110000011101000101110010001001101000000000001011000)  
) LUT6_1002 (
   .O(gates_414),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0010011001100101101101100000000111001011110011100011110110110001)  
) LUT6_1003 (
   .O(gates_145),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1010111011101011111000110111111001100010100111010011110011100010)  
) LUT6_1004 (
   .O(gates_1217),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1101100100011111100001110100111010101010010001100011101011011000)  
) LUT6_1005 (
   .O(gates_1301),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0001101010101100001011100110100000100110101000100110010100010100)  
) LUT6_1006 (
   .O(gates_252),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0111011010000111111000001100100000100110101001100101110110100000)  
) LUT6_1007 (
   .O(gates_474),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b0011000100110000110110101010111000011000010100000011110110111010)  
) LUT6_1008 (
   .O(gates_1424),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0001110010001100000110011111101011110111100110100101100010011100)  
) LUT6_1009 (
   .O(gates_534),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0111100000001100111110111000011011100111111001110000100011110101)  
) LUT6_1010 (
   .O(gates_1151),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1010100010010000111011100101110100001110101011000010101010100001)  
) LUT6_1011 (
   .O(gates_259),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0001111101101001010100111011010011001111110110111111101101011010)  
) LUT6_1012 (
   .O(gates_609),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1011001100011111001010110101110001101111000100010010101111111010)  
) LUT6_1013 (
   .O(gates_648),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b0111001100000110010101000100000010000111100100101001111011101001)  
) LUT6_1014 (
   .O(gates_235),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1101010000001110011101110010100011011110100010100010111011101010)  
) LUT6_1015 (
   .O(gates_1143),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1101001001000001101101110000001100010010001111100100011000000110)  
) LUT6_1016 (
   .O(gates_1439),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1011111010101101111000000010010011101101111010000000100110000010)  
) LUT6_1017 (
   .O(gates_490),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0110101100000101000111101110000110100111111011100001000011001111)  
) LUT6_1018 (
   .O(gates_256),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0000100101010110111000001101010001000110110111010011111001100101)  
) LUT6_1019 (
   .O(gates_966),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1010100000010001000101011100010000111010101011010010100110001100)  
) LUT6_1020 (
   .O(gates_1075),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0011011101111101111000010000001111010100101010110111010101111010)  
) LUT6_1021 (
   .O(gates_358),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0111100101000100110001101010100100000100100111011000010101001101)  
) LUT6_1022 (
   .O(gates_803),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0100011011100010111010101000010011101011101110001000110110100010)  
) LUT6_1023 (
   .O(gates_308),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0010111000011010010101111011100101111110011110111100111010000001)  
) LUT6_1024 (
   .O(gates_366),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b1000001000111000111101110011100111111110110010111000110000100001)  
) LUT6_1025 (
   .O(gates_431),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0101000100010101010011001000000011110001000011010111111001100001)  
) LUT6_1026 (
   .O(gates_195),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1110111101000100101101110101011001000110001011110010010101100101)  
) LUT6_1027 (
   .O(gates_425),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1100001000000111110010010100000101000001000000010110010101111101)  
) LUT6_1028 (
   .O(gates_714),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1011010001011101011001100111100001011011100101000001111001111100)  
) LUT6_1029 (
   .O(gates_114),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0100001110011000010101010111101110011000100010001100101100000011)  
) LUT6_1030 (
   .O(gates_184),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1010010000001001110100000001110101000101000001111110011100010010)  
) LUT6_1031 (
   .O(gates_222),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0101010110111000001101000000001111100000101100010111110011100000)  
) LUT6_1032 (
   .O(gates_1518),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0110100001100011110100100011000000011110100101001111011110111011)  
) LUT6_1033 (
   .O(gates_1026),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b0010111011010100000110000001101111011111011110110011101000011111)  
) LUT6_1034 (
   .O(gates_90),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1000001101100010101010101000110010110110010000100110100111111000)  
) LUT6_1035 (
   .O(gates_615),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0001011100111110010000000011010000111111100101010000100011010111)  
) LUT6_1036 (
   .O(gates_1225),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b0010111001000011001001100110011011100111001101011100110100000000)  
) LUT6_1037 (
   .O(gates_827),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0010110011101011111000000111000100101110000011001000000000011110)  
) LUT6_1038 (
   .O(gates_480),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0001111000011001011001000001110000110001101001110010110000011011)  
) LUT6_1039 (
   .O(gates_469),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0011010010110110011110101011001101001011011110010101001000110001)  
) LUT6_1040 (
   .O(gates_1440),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0100000111110110100101000001110000000111011110111011001111011010)  
) LUT6_1041 (
   .O(gates_804),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b0001101110001010001010110010101010111001010010000010011010100011)  
) LUT6_1042 (
   .O(gates_115),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b1000010111010010000110100110100110100011000100101111110110110101)  
) LUT6_1043 (
   .O(gates_302),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0111100110001111010000001101001100011000101100000010010100111011)  
) LUT6_1044 (
   .O(gates_971),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0111110001000010111100101100011101100011011001111001011010010100)  
) LUT6_1045 (
   .O(gates_1511),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0000011010010110110110111111010100111110011011111010001001001110)  
) LUT6_1046 (
   .O(gates_1246),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1101010011100010000101001000111101110110100111010100010110111011)  
) LUT6_1047 (
   .O(gates_1363),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b0111100011010101010101111000010110100101011110111011100101101111)  
) LUT6_1048 (
   .O(gates_530),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b1001110101101011010110001001011110101011001111111110000000001110)  
) LUT6_1049 (
   .O(gates_600),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0011010010111000100011000100010110011110010100001000011101111100)  
) LUT6_1050 (
   .O(gates_284),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0001111100110000101001000001100101111011100011011110001100100001)  
) LUT6_1051 (
   .O(gates_770),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0111101111101111010101001111000111100100110101111101001001000000)  
) LUT6_1052 (
   .O(gates_34),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1010011000000101000101010011100110011111111010011010000111101000)  
) LUT6_1053 (
   .O(gates_165),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0011011111110011100100100000001111101111111010010001111010110010)  
) LUT6_1054 (
   .O(gates_193),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b0100110110010001111111001101101001111011001001001001011111111100)  
) LUT6_1055 (
   .O(gates_800),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1001001001001100011001010111001100001110011101110000110011101010)  
) LUT6_1056 (
   .O(gates_462),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b0110000001000001101001000011101011000000001100010100000011101110)  
) LUT6_1057 (
   .O(gates_585),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1100010111111110101011100010110010011101110100011101110010001110)  
) LUT6_1058 (
   .O(gates_1054),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0101001100001010001100000001100011010101110001110010011110010110)  
) LUT6_1059 (
   .O(gates_653),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1011010100000011100110100011011110001100001110100001000111000000)  
) LUT6_1060 (
   .O(gates_869),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1111001000011000000110011101110011101110111010110000101110000001)  
) LUT6_1061 (
   .O(gates_989),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0010110000111000101111101100110100100110111101010110001001010000)  
) LUT6_1062 (
   .O(gates_1478),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0100110111011110001000000110011000101101000011100000001100001111)  
) LUT6_1063 (
   .O(gates_1331),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0100101010111111100000101000011000010010101111100110111111111110)  
) LUT6_1064 (
   .O(gates_842),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1111011100000100101111001100001000111111010100001001011100111111)  
) LUT6_1065 (
   .O(gates_650),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1000101100100110101110001011001000100111111111010010110001110001)  
) LUT6_1066 (
   .O(gates_645),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0010000100001010010010010111111001110100010111000010000001000011)  
) LUT6_1067 (
   .O(gates_1245),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0011010101100001001100000100010000110111111101000110100111011111)  
) LUT6_1068 (
   .O(gates_657),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1101110000000011010001000011001000010011011010010010000001111101)  
) LUT6_1069 (
   .O(gates_464),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b1101011010111110010011101100100101010011001101101111011000001011)  
) LUT6_1070 (
   .O(gates_167),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b1011110101111101001111110010011111100011101100101000001110101000)  
) LUT6_1071 (
   .O(gates_1386),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0111011111000011100011100110110111111110001010101101010011111111)  
) LUT6_1072 (
   .O(gates_678),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0101011100110011100000110001110110011110000000010000001111110101)  
) LUT6_1073 (
   .O(gates_1049),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0011001101000010011010011010011100011000101001101000101000101111)  
) LUT6_1074 (
   .O(gates_898),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0000101000110110110011010110000101110010101010001001011101001011)  
) LUT6_1075 (
   .O(gates_538),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0111010011001100100010111110111111011001110010010011001010001011)  
) LUT6_1076 (
   .O(gates_845),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b1000011000100000110001110100000010110001000010000000011010010101)  
) LUT6_1077 (
   .O(gates_652),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0010011100011011000011110110101010110011011011001000000010001011)  
) LUT6_1078 (
   .O(gates_387),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0000110000011011111100001011011110101000001011000110110000001010)  
) LUT6_1079 (
   .O(gates_1370),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0001100011110110001000010000001011110111011001100001010010110000)  
) LUT6_1080 (
   .O(gates_1022),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1111001000111110001000001111011001101101100000110001001101100110)  
) LUT6_1081 (
   .O(gates_864),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1000000100100010010100101101001101011101111110110111111011011011)  
) LUT6_1082 (
   .O(gates_1251),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b0011000101100101010010001101000010111000100000010010010111000111)  
) LUT6_1083 (
   .O(gates_1086),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1111000101110000111100111001100000100010111111110101101010100000)  
) LUT6_1084 (
   .O(gates_47),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b0110001100000111010010001011011101101101111111111110110101101000)  
) LUT6_1085 (
   .O(gates_1479),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1001010010110101110110001000010001111011100101101110010001000101)  
) LUT6_1086 (
   .O(gates_1273),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0110010011000101100101100101100111100111010000001111011110001110)  
) LUT6_1087 (
   .O(gates_685),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0111000100011000111000111110101110010101101100110011010111101101)  
) LUT6_1088 (
   .O(gates_741),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0101011010101101110100011111001000010110111110110110111101111000)  
) LUT6_1089 (
   .O(gates_430),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0101110000101010110000101011001111011010111001010110100100100101)  
) LUT6_1090 (
   .O(gates_761),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b0010010010001001101001010110001101100010111010011010001111011010)  
) LUT6_1091 (
   .O(gates_1162),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0010100101101101001001110101110000001110110010010000101111101100)  
) LUT6_1092 (
   .O(gates_1423),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1100011010001111011011010100000011101101100100100101111101001110)  
) LUT6_1093 (
   .O(gates_1067),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b0010110000000100101011000101010111000001001111011100100001101110)  
) LUT6_1094 (
   .O(gates_540),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1010110111110000111011111101010111101110010101100000001011100110)  
) LUT6_1095 (
   .O(gates_94),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1001101001111001111111100001011001100110001000111001001101001101)  
) LUT6_1096 (
   .O(gates_1297),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0110000001110101111001011111100011100111001001001100110101001011)  
) LUT6_1097 (
   .O(gates_334),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010111011001001011001100011101010000011100000101110001010111101)  
) LUT6_1098 (
   .O(gates_529),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b1011001010111100100101010011010011010101110001100001001001101011)  
) LUT6_1099 (
   .O(gates_794),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0010011010000101010110110101111010100111011011101110100110101111)  
) LUT6_1100 (
   .O(gates_590),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0010001000101110001011100001111111100110100010110110111100110011)  
) LUT6_1101 (
   .O(gates_1501),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0010001111011000010011100100111110010001101100011101110101000001)  
) LUT6_1102 (
   .O(gates_467),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0110010001000111010001011101111111101100000011110111101100100010)  
) LUT6_1103 (
   .O(gates_1184),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1001101001010011110100001111011000000010000101100001010101011001)  
) LUT6_1104 (
   .O(gates_403),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1110001001111010100101001111011000110000111110010011101111110011)  
) LUT6_1105 (
   .O(gates_1183),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0000101011100011011000110010110001011010111011101101101101100000)  
) LUT6_1106 (
   .O(gates_152),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1100010100100001011111100110100011100101101110101000010001101111)  
) LUT6_1107 (
   .O(gates_1257),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b1101000000010011110110001001101110001011100000100010010111100110)  
) LUT6_1108 (
   .O(gates_526),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1101000101011010100111011010100101010110010000110111110111110000)  
) LUT6_1109 (
   .O(gates_28),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1111110011101111010010011111010000011010001001000101011111010100)  
) LUT6_1110 (
   .O(gates_558),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1001010010000110010010010101111101000100000010011101111000101110)  
) LUT6_1111 (
   .O(gates_422),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b1100011110010101000010110000101011001100000001100111000011101101)  
) LUT6_1112 (
   .O(gates_1293),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1101111101010100010110100100100011100111011011111110111000001001)  
) LUT6_1113 (
   .O(gates_1043),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0100100101101110110001100111000010111000010111011110000101011001)  
) LUT6_1114 (
   .O(gates_146),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b0010011111100111000011111110100111010111111010100001110101001111)  
) LUT6_1115 (
   .O(gates_461),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b0110011110111001011010101100001011010100111010110110101110010000)  
) LUT6_1116 (
   .O(gates_834),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b1011010010001010011010001110010110110101010111111111001101100010)  
) LUT6_1117 (
   .O(gates_1029),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0101100000110110101011100010010010010011100111010010011010000011)  
) LUT6_1118 (
   .O(gates_1339),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0011011110100100000000111111010001101001110000011110001110010001)  
) LUT6_1119 (
   .O(gates_545),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0101010100101011010110010101111000101110100100101111010110100101)  
) LUT6_1120 (
   .O(gates_587),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b0000000000000011110101000011010010110010100101011111110010001110)  
) LUT6_1121 (
   .O(gates_918),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b0001010101101000011110001010001011111101101011011010001101000111)  
) LUT6_1122 (
   .O(gates_1356),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b1101000000111011110100100110110100110010100000000101000100010100)  
) LUT6_1123 (
   .O(gates_91),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b0010011101100011011001000000111001111000110101101010010001100101)  
) LUT6_1124 (
   .O(gates_231),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0100000011101110000011001111001111001011110010001000011011110111)  
) LUT6_1125 (
   .O(gates_14),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1111111101010011100111001110100110001001011111011000000111110101)  
) LUT6_1126 (
   .O(gates_1455),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000010000000010110000001010001011011000011001110111111000100110)  
) LUT6_1127 (
   .O(gates_1254),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0011101100111100100011001010011011100100000010010111111101000111)  
) LUT6_1128 (
   .O(gates_319),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0110100000110110100110011111011101100011111010010010110111111010)  
) LUT6_1129 (
   .O(gates_125),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1110110111010101000011000000101001001001001111001011111011001101)  
) LUT6_1130 (
   .O(gates_389),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1000110001001110100001011011101101111111100111011000101100001100)  
) LUT6_1131 (
   .O(gates_75),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1100111111110001100010001011001001000111011000110100000100010010)  
) LUT6_1132 (
   .O(gates_53),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b0101011011100010111011100111111000111000001000001101100011000000)  
) LUT6_1133 (
   .O(gates_1304),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b0101011001010010001010001111111000101011110010100011100001101011)  
) LUT6_1134 (
   .O(gates_248),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0000111100000100101001111100000100111100100111110100001011100001)  
) LUT6_1135 (
   .O(gates_511),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b0001110001000111100101000100011100000011011101010101101110100111)  
) LUT6_1136 (
   .O(gates_265),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b0011000011011101110011000011110101000011111001100000100111111111)  
) LUT6_1137 (
   .O(gates_77),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1110110000111110100110111000110010110011000101011011000101010100)  
) LUT6_1138 (
   .O(gates_1328),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0100101111101100011010111111010011010111101110010111111101011100)  
) LUT6_1139 (
   .O(gates_390),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b0011111111010011110000010101101010101101110101000011010010110011)  
) LUT6_1140 (
   .O(gates_1549),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b1110010100111101001011000011100101010010100111100000111111000010)  
) LUT6_1141 (
   .O(gates_124),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0001101000011001101111110100101111110001001111101011101100111101)  
) LUT6_1142 (
   .O(gates_1091),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b0000010011000110101001100001000001110000111010010100011100111100)  
) LUT6_1143 (
   .O(gates_123),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1111111110010110001101011010110111001000011101000101001100000011)  
) LUT6_1144 (
   .O(gates_50),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0110101100111010111011000101010010110010101101100011001010000100)  
) LUT6_1145 (
   .O(gates_424),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1010111011001011101110001011100110011010100100101001101011010011)  
) LUT6_1146 (
   .O(gates_742),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0110000010011111001000110010010111011110111000110011010010010110)  
) LUT6_1147 (
   .O(gates_347),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0001011101010100111000010000101100011001011001001100110001110001)  
) LUT6_1148 (
   .O(gates_1393),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1011100110001011101110001010011111000101011011001100011111000101)  
) LUT6_1149 (
   .O(gates_1153),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b1100010100010010000110101010011001001111101110100111011000010101)  
) LUT6_1150 (
   .O(gates_1312),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1100111101000111110000111110000100101100100101000000001111001111)  
) LUT6_1151 (
   .O(gates_571),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b0110100010111010100001010110011100011111100010100101111010101011)  
) LUT6_1152 (
   .O(gates_234),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b0010010010000000011010100101100110011100111001101000111101110010)  
) LUT6_1153 (
   .O(gates_607),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0100111010010100101100111000111100011010100110000100000010000000)  
) LUT6_1154 (
   .O(gates_606),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1101101111000010101011000101000000000111100101110011111111101110)  
) LUT6_1155 (
   .O(gates_878),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1001010110010010000110111101110010110010001010000011001011010010)  
) LUT6_1156 (
   .O(gates_209),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0010010101111000101010110010010010001011001000111111100001101011)  
) LUT6_1157 (
   .O(gates_1490),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b1110110101111000001011100110010010111100000001010100111011010110)  
) LUT6_1158 (
   .O(gates_182),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b0110111001000111110011111110110011101001110010001101011101011011)  
) LUT6_1159 (
   .O(gates_1306),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b1011101111011111010000001000101011010010110010000001001110000011)  
) LUT6_1160 (
   .O(gates_207),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0110010111000111100010110010111111110001101100101001000010100000)  
) LUT6_1161 (
   .O(gates_658),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b0110000101011011001000000110011000110100010001001111101010010111)  
) LUT6_1162 (
   .O(gates_582),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0111100110011010110000100100010011111101011010101010010000111101)  
) LUT6_1163 (
   .O(gates_1438),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0010100001110100011101011000110111001100110101000010100001001101)  
) LUT6_1164 (
   .O(gates_317),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1111101101101001001011011010101001001111111011010101010111011011)  
) LUT6_1165 (
   .O(gates_786),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b0101001110000001001110100101100011001011011101111110101100111111)  
) LUT6_1166 (
   .O(gates_1280),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0001100110000110110111110101101001111101001101100110100101110001)  
) LUT6_1167 (
   .O(gates_541),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b1001100001110011100010001111110000110100111011010101010011000111)  
) LUT6_1168 (
   .O(gates_1453),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0000010110111101111100010111001111100011101010111101010011110000)  
) LUT6_1169 (
   .O(gates_776),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1101011111100010010011000110001000010001011010000100000001110111)  
) LUT6_1170 (
   .O(gates_1209),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0101011110000100110000011001011110001001110010011011110010000110)  
) LUT6_1171 (
   .O(gates_627),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0010010100100011111010110001100110111101111111100100100110101000)  
) LUT6_1172 (
   .O(gates_367),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0111000000101010100001011001111100101001111001011110000000000010)  
) LUT6_1173 (
   .O(gates_176),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0011001010010011011111111011010010101110110101111111010101011111)  
) LUT6_1174 (
   .O(gates_398),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0101101011010000110110010100100100000010110011000011001010000101)  
) LUT6_1175 (
   .O(gates_5),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b1010110111000001100010110010000011111011001001111001100010110110)  
) LUT6_1176 (
   .O(gates_300),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b0001011111100010000011110101111001101011110111100000011111100100)  
) LUT6_1177 (
   .O(gates_224),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b1001101100000010010111100000101111000111100100111001011100100100)  
) LUT6_1178 (
   .O(gates_1109),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1101100100101111101001111111110010101010101011001001011000001011)  
) LUT6_1179 (
   .O(gates_902),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b1000101000111100101110100100010011100100101000110011100011110111)  
) LUT6_1180 (
   .O(gates_101),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1010110000000111100101001000001011010101110000101111111100111110)  
) LUT6_1181 (
   .O(gates_1314),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0110001110000000000101010111001101101000101100001011010110111110)  
) LUT6_1182 (
   .O(gates_1024),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1111000001101001100001010110100111110101001100100001111001110110)  
) LUT6_1183 (
   .O(gates_532),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1001111010111000100011011101011100010111110110001101101010100011)  
) LUT6_1184 (
   .O(gates_1072),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010000000101011000101111001111011111000100001001101111010000101)  
) LUT6_1185 (
   .O(gates_364),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b0100100110100111101110110111101011001100110110110111000000100100)  
) LUT6_1186 (
   .O(gates_212),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b1010111100010101000100010010100100010001001011011000011110001000)  
) LUT6_1187 (
   .O(gates_1216),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b0001101111101100111010101011000011000111000001110101111001010110)  
) LUT6_1188 (
   .O(gates_1291),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b1001000011111100101010100011001110111001000011011000100101100110)  
) LUT6_1189 (
   .O(gates_843),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b1111010011001100110010001010110100011100001000101100110101000111)  
) LUT6_1190 (
   .O(gates_586),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1001100101011001111001010000010101111111000010110010101110111000)  
) LUT6_1191 (
   .O(gates_122),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b0101100110001110100100000011010011011100110011110001101110001010)  
) LUT6_1192 (
   .O(gates_861),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1110010101101101001110010011010101101110100011011011010000110000)  
) LUT6_1193 (
   .O(gates_100),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1101000010110010100000111100000110011111101010111101011010000100)  
) LUT6_1194 (
   .O(gates_1237),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0110010111101001000101101100011010101011010110101011001001011110)  
) LUT6_1195 (
   .O(gates_596),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0001100000010101011001101100000011111110011011101001010000111101)  
) LUT6_1196 (
   .O(gates_956),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b1001011111110100001100111000111000000111011001100010011010101100)  
) LUT6_1197 (
   .O(gates_149),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b0110010100101111000001111011111010111010010010101110000100010000)  
) LUT6_1198 (
   .O(gates_856),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b1001001000100000110110001110100110110100110111011101100010011111)  
) LUT6_1199 (
   .O(gates_766),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1100111001010000101110101010110000111011101000011111100100011110)  
) LUT6_1200 (
   .O(gates_373),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1100011100100111101011001001110001100100111111111000100011001001)  
) LUT6_1201 (
   .O(gates_1421),
   .I0(InputBits[200]),
   .I1(InputBits[118]),
   .I2(InputBits[525]),
   .I3(InputBits[408]),
   .I4(InputBits[7]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0100100100111100011001101100010011100100111101101110010111001000)  
) LUT6_1202 (
   .O(gates_73),
   .I0(InputBits[433]),
   .I1(InputBits[76]),
   .I2(InputBits[386]),
   .I3(InputBits[92]),
   .I4(InputBits[477]),
   .I5(InputBits[360])
);
LUT6 #(
   .INIT(64'b1001111101111110001011001111110001101001010011110001101110000101)  
) LUT6_1203 (
   .O(gates_1156),
   .I0(InputBits[275]),
   .I1(InputBits[217]),
   .I2(InputBits[363]),
   .I3(InputBits[341]),
   .I4(InputBits[244]),
   .I5(InputBits[252])
);
LUT6 #(
   .INIT(64'b0001001000100110000100000010100101001011101010010011000011010110)  
) LUT6_1204 (
   .O(gates_943),
   .I0(InputBits[192]),
   .I1(InputBits[73]),
   .I2(InputBits[537]),
   .I3(InputBits[391]),
   .I4(InputBits[557]),
   .I5(InputBits[260])
);
LUT6 #(
   .INIT(64'b1110011111010010111101101111111001101101111100010111010001101001)  
) LUT6_1205 (
   .O(gates_1321),
   .I0(InputBits[403]),
   .I1(InputBits[320]),
   .I2(InputBits[115]),
   .I3(InputBits[145]),
   .I4(InputBits[8]),
   .I5(InputBits[276])
);
LUT6 #(
   .INIT(64'b1000100011010000110100010011111100000101100010100101100110100101)  
) LUT6_1206 (
   .O(gates_914),
   .I0(InputBits[68]),
   .I1(InputBits[307]),
   .I2(InputBits[132]),
   .I3(InputBits[328]),
   .I4(InputBits[72]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0101000010110010111011010010101111010100000001111110110010001010)  
) LUT6_1207 (
   .O(gates_921),
   .I0(InputBits[208]),
   .I1(InputBits[298]),
   .I2(InputBits[106]),
   .I3(InputBits[348]),
   .I4(InputBits[299]),
   .I5(InputBits[124])
);
LUT6 #(
   .INIT(64'b0101011110000101111101010000111001111010010000101011101110011001)  
) LUT6_1208 (
   .O(gates_491),
   .I0(InputBits[308]),
   .I1(InputBits[225]),
   .I2(InputBits[5]),
   .I3(InputBits[296]),
   .I4(InputBits[456]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b0010101111011011011010010110111001110110101000011000001001001011)  
) LUT6_1209 (
   .O(gates_156),
   .I0(InputBits[284]),
   .I1(InputBits[100]),
   .I2(InputBits[452]),
   .I3(InputBits[480]),
   .I4(InputBits[53]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0001001010001110101111111100011100101011011001110000010000001001)  
) LUT6_1210 (
   .O(gates_835),
   .I0(InputBits[249]),
   .I1(InputBits[550]),
   .I2(InputBits[450]),
   .I3(InputBits[130]),
   .I4(InputBits[3]),
   .I5(InputBits[30])
);
LUT6 #(
   .INIT(64'b1101110011101010000001010110110101100110100110100111100110110011)  
) LUT6_1211 (
   .O(gates_1132),
   .I0(InputBits[455]),
   .I1(InputBits[432]),
   .I2(InputBits[66]),
   .I3(InputBits[165]),
   .I4(InputBits[462]),
   .I5(InputBits[302])
);
LUT6 #(
   .INIT(64'b1000101101110000111111110011101101111001010000010110110111111001)  
) LUT6_1212 (
   .O(gates_132),
   .I0(InputBits[57]),
   .I1(InputBits[385]),
   .I2(InputBits[120]),
   .I3(InputBits[399]),
   .I4(InputBits[131]),
   .I5(InputBits[454])
);
LUT6 #(
   .INIT(64'b0101000111011111110001011100100000111001110111010010000110100100)  
) LUT6_1213 (
   .O(gates_595),
   .I0(InputBits[436]),
   .I1(InputBits[256]),
   .I2(InputBits[239]),
   .I3(InputBits[240]),
   .I4(InputBits[113]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0111110010001101100000111101011000011110100101000001110101011011)  
) LUT6_1214 (
   .O(gates_1468),
   .I0(InputBits[488]),
   .I1(InputBits[55]),
   .I2(InputBits[316]),
   .I3(InputBits[481]),
   .I4(InputBits[380]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1010101110011001110011011111100100101110000010100010011000101111)  
) LUT6_1215 (
   .O(gates_946),
   .I0(InputBits[558]),
   .I1(InputBits[335]),
   .I2(InputBits[84]),
   .I3(InputBits[410]),
   .I4(InputBits[379]),
   .I5(InputBits[446])
);
LUT6 #(
   .INIT(64'b0111001011001110000110010001001110011011011001001110000001111000)  
) LUT6_1216 (
   .O(gates_129),
   .I0(InputBits[78]),
   .I1(InputBits[114]),
   .I2(InputBits[63]),
   .I3(InputBits[21]),
   .I4(InputBits[474]),
   .I5(InputBits[313])
);
LUT6 #(
   .INIT(64'b1101011010010001001011000101011001110110111100100000100000011100)  
) LUT6_1217 (
   .O(gates_96),
   .I0(InputBits[64]),
   .I1(InputBits[435]),
   .I2(InputBits[143]),
   .I3(InputBits[133]),
   .I4(InputBits[285]),
   .I5(InputBits[219])
);
LUT6 #(
   .INIT(64'b1010011111111000110110011110101011101100100001110101111010111110)  
) LUT6_1218 (
   .O(gates_828),
   .I0(InputBits[332]),
   .I1(InputBits[262]),
   .I2(InputBits[147]),
   .I3(InputBits[184]),
   .I4(InputBits[368]),
   .I5(InputBits[354])
);
LUT6 #(
   .INIT(64'b0100001111111110100111101000100111110000111111010001100101110111)  
) LUT6_1219 (
   .O(gates_1235),
   .I0(InputBits[352]),
   .I1(InputBits[168]),
   .I2(InputBits[530]),
   .I3(InputBits[314]),
   .I4(InputBits[416]),
   .I5(InputBits[315])
);
LUT6 #(
   .INIT(64'b1001000100001100010101011110011010010111000111000011001010010100)  
) LUT6_1220 (
   .O(gates_1150),
   .I0(InputBits[236]),
   .I1(InputBits[559]),
   .I2(InputBits[31]),
   .I3(InputBits[524]),
   .I4(InputBits[282]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0111011100101101110001111111100101111010010000111011010111110111)  
) LUT6_1221 (
   .O(gates_610),
   .I0(InputBits[248]),
   .I1(InputBits[213]),
   .I2(InputBits[501]),
   .I3(InputBits[243]),
   .I4(InputBits[40]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1011110111001010101001010100011010101001111001101100100110100100)  
) LUT6_1222 (
   .O(gates_1429),
   .I0(InputBits[52]),
   .I1(InputBits[330]),
   .I2(InputBits[43]),
   .I3(InputBits[400]),
   .I4(InputBits[412]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1011001100111001100100100111011011001110110101000010110101101011)  
) LUT6_1223 (
   .O(gates_1426),
   .I0(InputBits[235]),
   .I1(InputBits[500]),
   .I2(InputBits[292]),
   .I3(InputBits[362]),
   .I4(InputBits[108]),
   .I5(InputBits[107])
);
LUT6 #(
   .INIT(64'b0101101100101010100111101011111111011000001111110000101111101001)  
) LUT6_1224 (
   .O(gates_225),
   .I0(InputBits[25]),
   .I1(InputBits[547]),
   .I2(InputBits[326]),
   .I3(InputBits[270]),
   .I4(InputBits[451]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0110100111110011101110000101100101011010111000111001101001011110)  
) LUT6_1225 (
   .O(gates_1498),
   .I0(InputBits[357]),
   .I1(InputBits[301]),
   .I2(InputBits[398]),
   .I3(InputBits[420]),
   .I4(InputBits[228]),
   .I5(InputBits[4])
);
LUT6 #(
   .INIT(64'b1001010101100001000001010001110101101110001001100100100001010000)  
) LUT6_1226 (
   .O(gates_40),
   .I0(InputBits[6]),
   .I1(InputBits[424]),
   .I2(InputBits[99]),
   .I3(InputBits[476]),
   .I4(InputBits[247]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001111000000001001100100011001001001000101110011101011100001010)  
) LUT6_1227 (
   .O(gates_277),
   .I0(InputBits[505]),
   .I1(InputBits[407]),
   .I2(InputBits[79]),
   .I3(InputBits[461]),
   .I4(InputBits[345]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0101011111101111110110010010010010100111101011000011000111100111)  
) LUT6_1228 (
   .O(gates_1294),
   .I0(InputBits[241]),
   .I1(InputBits[134]),
   .I2(InputBits[50]),
   .I3(InputBits[374]),
   .I4(InputBits[289]),
   .I5(InputBits[49])
);
LUT6 #(
   .INIT(64'b1001100011111000001100111000010110011010000111110111001010011111)  
) LUT6_1229 (
   .O(gates_1224),
   .I0(InputBits[81]),
   .I1(InputBits[404]),
   .I2(InputBits[526]),
   .I3(InputBits[553]),
   .I4(InputBits[163]),
   .I5(InputBits[506])
);
LUT6 #(
   .INIT(64'b1011001111011000111111010010000010010010011001100111000001100000)  
) LUT6_1230 (
   .O(gates_561),
   .I0(InputBits[365]),
   .I1(InputBits[51]),
   .I2(InputBits[469]),
   .I3(InputBits[569]),
   .I4(InputBits[375]),
   .I5(InputBits[12])
);
LUT6 #(
   .INIT(64'b0100000110110100101000100110101001110111011110100101111110101110)  
) LUT6_1231 (
   .O(gates_443),
   .I0(InputBits[261]),
   .I1(InputBits[512]),
   .I2(InputBits[103]),
   .I3(InputBits[264]),
   .I4(InputBits[572]),
   .I5(InputBits[287])
);
LUT6 #(
   .INIT(64'b1111101011010010001001100011101110011001100001100101011111101001)  
) LUT6_1232 (
   .O(gates_1551),
   .I0(InputBits[267]),
   .I1(InputBits[358]),
   .I2(InputBits[46]),
   .I3(InputBits[234]),
   .I4(InputBits[364]),
   .I5(InputBits[279])
);
LUT6 #(
   .INIT(64'b1010001000010010100100010100101100011100001101011001111010111001)  
) LUT6_1233 (
   .O(gates_676),
   .I0(InputBits[257]),
   .I1(InputBits[281]),
   .I2(InputBits[182]),
   .I3(InputBits[158]),
   .I4(InputBits[155]),
   .I5(InputBits[371])
);
LUT6 #(
   .INIT(64'b1111101001010101100000100001000010011111101010000110111111010100)  
) LUT6_1234 (
   .O(gates_255),
   .I0(InputBits[271]),
   .I1(InputBits[490]),
   .I2(InputBits[14]),
   .I3(InputBits[156]),
   .I4(InputBits[541]),
   .I5(InputBits[492])
);
LUT6 #(
   .INIT(64'b0001100000110111110001011101101110001000000101111010110000111100)  
) LUT6_1235 (
   .O(gates_552),
   .I0(InputBits[190]),
   .I1(InputBits[318]),
   .I2(InputBits[425]),
   .I3(InputBits[463]),
   .I4(InputBits[389]),
   .I5(InputBits[439])
);
LUT6 #(
   .INIT(64'b1110100001010111001101011101011001110101001110001100111111111000)  
) LUT6_1236 (
   .O(gates_1194),
   .I0(InputBits[369]),
   .I1(InputBits[430]),
   .I2(InputBits[567]),
   .I3(InputBits[510]),
   .I4(InputBits[449]),
   .I5(InputBits[70])
);
LUT6 #(
   .INIT(64'b0110111000010000111010100011011111010010111000110111111100101000)  
) LUT6_1237 (
   .O(gates_1268),
   .I0(InputBits[278]),
   .I1(InputBits[61]),
   .I2(InputBits[434]),
   .I3(InputBits[438]),
   .I4(InputBits[98]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1110110001101110010010101100101100111000001110001101010110100100)  
) LUT6_1238 (
   .O(gates_1398),
   .I0(InputBits[502]),
   .I1(InputBits[135]),
   .I2(InputBits[45]),
   .I3(InputBits[531]),
   .I4(InputBits[413]),
   .I5(InputBits[22])
);
LUT6 #(
   .INIT(64'b1111100001100111011110101101110101101110111101110100000110010100)  
) LUT6_1239 (
   .O(gates_107),
   .I0(InputBits[382]),
   .I1(InputBits[376]),
   .I2(InputBits[237]),
   .I3(InputBits[109]),
   .I4(InputBits[176]),
   .I5(InputBits[544])
);
LUT6 #(
   .INIT(64'b1100010011110110101000111111001001011001001001001111000001011100)  
) LUT6_1240 (
   .O(gates_1544),
   .I0(InputBits[204]),
   .I1(InputBits[518]),
   .I2(InputBits[90]),
   .I3(InputBits[126]),
   .I4(InputBits[29]),
   .I5(InputBits[390])
);
LUT6 #(
   .INIT(64'b0000110010101011111010111100010100110100111011001111001011001101)  
) LUT6_1241 (
   .O(gates_620),
   .I0(InputBits[136]),
   .I1(InputBits[334]),
   .I2(InputBits[402]),
   .I3(InputBits[312]),
   .I4(InputBits[294]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1010000011101001111110010101101010010100100111011000001011000001)  
) LUT6_1242 (
   .O(gates_829),
   .I0(InputBits[283]),
   .I1(InputBits[185]),
   .I2(InputBits[28]),
   .I3(InputBits[311]),
   .I4(InputBits[231]),
   .I5(InputBits[503])
);
LUT6 #(
   .INIT(64'b0010101101001110010110000110101111110100001000010001010100001001)  
) LUT6_1243 (
   .O(gates_120),
   .I0(InputBits[485]),
   .I1(InputBits[26]),
   .I2(InputBits[542]),
   .I3(InputBits[258]),
   .I4(InputBits[548]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1110110001101001001100001001100101000111100110110010011101010010)  
) LUT6_1244 (
   .O(gates_82),
   .I0(InputBits[27]),
   .I1(InputBits[198]),
   .I2(InputBits[297]),
   .I3(InputBits[336]),
   .I4(InputBits[138]),
   .I5(InputBits[191])
);
LUT6 #(
   .INIT(64'b1100011001000000111101010110100010110010110101100111100111111010)  
) LUT6_1245 (
   .O(gates_939),
   .I0(InputBits[286]),
   .I1(InputBits[36]),
   .I2(InputBits[419]),
   .I3(InputBits[161]),
   .I4(InputBits[9]),
   .I5(InputBits[353])
);
LUT6 #(
   .INIT(64'b0100101101011110010010110001111001101100011011110010000111100111)  
) LUT6_1246 (
   .O(gates_218),
   .I0(InputBits[277]),
   .I1(InputBits[346]),
   .I2(InputBits[127]),
   .I3(InputBits[268]),
   .I4(InputBits[370]),
   .I5(InputBits[459])
);
LUT6 #(
   .INIT(64'b1101111010111100000101100110010011000010110001011110100000011010)  
) LUT6_1247 (
   .O(gates_489),
   .I0(InputBits[414]),
   .I1(InputBits[229]),
   .I2(InputBits[169]),
   .I3(InputBits[331]),
   .I4(InputBits[201]),
   .I5(InputBits[423])
);
LUT6 #(
   .INIT(64'b1101111010101111010101110001000100111011100110010101011001000000)  
) LUT6_1248 (
   .O(gates_151),
   .I0(InputBits[245]),
   .I1(InputBits[196]),
   .I2(InputBits[150]),
   .I3(InputBits[495]),
   .I4(InputBits[180]),
   .I5(InputBits[377])
);
LUT6 #(
   .INIT(64'b1000000001000101000100101001101001011000111000000000001111101000)  
) LUT6_1249 (
   .O(gates_410),
   .I0(InputBits[274]),
   .I1(InputBits[445]),
   .I2(InputBits[227]),
   .I3(InputBits[508]),
   .I4(InputBits[69]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b1111111111110100011110110011101110011000110001001110100111111010)  
) LUT6_1250 (
   .O(gates_1042),
   .I0(InputBits[305]),
   .I1(InputBits[87]),
   .I2(InputBits[540]),
   .I3(InputBits[504]),
   .I4(InputBits[493]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0110100101001000101011011100110110010100000110001010011101100111)  
) LUT6_1251 (
   .O(gates_214),
   .I0(InputBits[361]),
   .I1(InputBits[266]),
   .I2(InputBits[197]),
   .I3(InputBits[82]),
   .I4(InputBits[426]),
   .I5(InputBits[112])
);
LUT6 #(
   .INIT(64'b1100010101010011010000100111101101101110010010011001011000010011)  
) LUT6_1252 (
   .O(gates_104),
   .I0(InputBits[177]),
   .I1(InputBits[67]),
   .I2(InputBits[202]),
   .I3(InputBits[556]),
   .I4(InputBits[300]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1000000101010111000111010001101010000011011000111011011101001000)  
) LUT6_1253 (
   .O(gates_257),
   .I0(InputBits[521]),
   .I1(InputBits[513]),
   .I2(InputBits[566]),
   .I3(InputBits[467]),
   .I4(InputBits[232]),
   .I5(InputBits[2])
);
LUT6 #(
   .INIT(64'b0110010001000011110110110110001110011011010000101110000010001100)  
) LUT6_1254 (
   .O(gates_58),
   .I0(InputBits[255]),
   .I1(InputBits[265]),
   .I2(InputBits[464]),
   .I3(InputBits[555]),
   .I4(InputBits[366]),
   .I5(InputBits[80])
);
LUT6 #(
   .INIT(64'b1110011010100101011001110101001101111000101110000110100000111001)  
) LUT6_1255 (
   .O(gates_1320),
   .I0(InputBits[440]),
   .I1(InputBits[458]),
   .I2(InputBits[441]),
   .I3(InputBits[102]),
   .I4(InputBits[457]),
   .I5(InputBits[397])
);
LUT6 #(
   .INIT(64'b0110000001101010001111101101000111101100000011110100100010000101)  
) LUT6_1256 (
   .O(gates_903),
   .I0(InputBits[162]),
   .I1(InputBits[562]),
   .I2(InputBits[499]),
   .I3(InputBits[105]),
   .I4(InputBits[409]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0111011111001000111000100110110001011011001101000110100100100001)  
) LUT6_1257 (
   .O(gates_140),
   .I0(InputBits[317]),
   .I1(InputBits[230]),
   .I2(InputBits[478]),
   .I3(InputBits[273]),
   .I4(InputBits[47]),
   .I5(InputBits[343])
);
LUT6 #(
   .INIT(64'b1000111000100010010100011101111110011100110011110100000001110100)  
) LUT6_1258 (
   .O(gates_1531),
   .I0(InputBits[373]),
   .I1(InputBits[573]),
   .I2(InputBits[269]),
   .I3(InputBits[473]),
   .I4(InputBits[203]),
   .I5(InputBits[405])
);
LUT6 #(
   .INIT(64'b0101101000010010010101000010010100010100100111000101001101101011)  
) LUT6_1259 (
   .O(gates_682),
   .I0(InputBits[254]),
   .I1(InputBits[211]),
   .I2(InputBits[507]),
   .I3(InputBits[381]),
   .I4(InputBits[442]),
   .I5(InputBits[337])
);
LUT6 #(
   .INIT(64'b0010000110101011000010000011111000001010100101101111010110110100)  
) LUT6_1260 (
   .O(gates_542),
   .I0(InputBits[212]),
   .I1(InputBits[323]),
   .I2(InputBits[415]),
   .I3(InputBits[533]),
   .I4(InputBits[329]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1011101011010000110001011100001011111011000010011010111111100111)  
) LUT6_1261 (
   .O(gates_314),
   .I0(InputBits[333]),
   .I1(InputBits[179]),
   .I2(InputBits[242]),
   .I3(InputBits[546]),
   .I4(InputBits[206]),
   .I5(InputBits[538])
);
LUT6 #(
   .INIT(64'b1101110101011111110000010110101101100010001001110001001100100100)  
) LUT6_1262 (
   .O(gates_1110),
   .I0(InputBits[528]),
   .I1(InputBits[173]),
   .I2(InputBits[93]),
   .I3(InputBits[37]),
   .I4(InputBits[293]),
   .I5(InputBits[71])
);
LUT6 #(
   .INIT(64'b0110010000101101000111101001001100100001101111100000000001100111)  
) LUT6_1263 (
   .O(gates_139),
   .I0(InputBits[166]),
   .I1(InputBits[561]),
   .I2(InputBits[448]),
   .I3(InputBits[199]),
   .I4(InputBits[119]),
   .I5(InputBits[83])
);
LUT6 #(
   .INIT(64'b0110110001110100010101101111101000001000100110110010001001101101)  
) LUT6_1264 (
   .O(gates_361),
   .I0(InputBits[444]),
   .I1(InputBits[122]),
   .I2(InputBits[13]),
   .I3(InputBits[194]),
   .I4(InputBits[178]),
   .I5(InputBits[575])
);
LUT6 #(
   .INIT(64'b0100010010101000000000011011011110110111011101100110101010110001)  
) LUT6_1265 (
   .O(gates_49),
   .I0(InputBits[1]),
   .I1(InputBits[170]),
   .I2(InputBits[460]),
   .I3(InputBits[195]),
   .I4(InputBits[218]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1001011001000100011000001100101100101010000000011111001011110100)  
) LUT6_1266 (
   .O(gates_42),
   .I0(InputBits[535]),
   .I1(InputBits[186]),
   .I2(InputBits[406]),
   .I3(InputBits[74]),
   .I4(InputBits[250]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1000100111000000111001000001110000100001111101100101001101010010)  
) LUT6_1267 (
   .O(gates_1508),
   .I0(InputBits[16]),
   .I1(InputBits[325]),
   .I2(InputBits[129]),
   .I3(InputBits[378]),
   .I4(InputBits[207]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0000100101011101011101101101100101101011011011111101010010110011)  
) LUT6_1268 (
   .O(gates_356),
   .I0(InputBits[523]),
   .I1(InputBits[189]),
   .I2(InputBits[56]),
   .I3(InputBits[520]),
   .I4(InputBits[142]),
   .I5(InputBits[489])
);
LUT6 #(
   .INIT(64'b0110000011111011011100111101110101101111010101001111000010110110)  
) LUT6_1269 (
   .O(gates_194),
   .I0(InputBits[388]),
   .I1(InputBits[251]),
   .I2(InputBits[384]),
   .I3(InputBits[466]),
   .I4(InputBits[157]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1101111000110100001001100011111000011101001101001111001011111100)  
) LUT6_1270 (
   .O(gates_153),
   .I0(InputBits[327]),
   .I1(InputBits[539]),
   .I2(InputBits[395]),
   .I3(InputBits[295]),
   .I4(InputBits[153]),
   .I5(InputBits[140])
);
LUT6 #(
   .INIT(64'b0011010000011001110010111110101000001110000011010101110010011110)  
) LUT6_1271 (
   .O(gates_232),
   .I0(InputBits[85]),
   .I1(InputBits[172]),
   .I2(InputBits[321]),
   .I3(InputBits[543]),
   .I4(InputBits[23]),
   .I5(InputBits[560])
);
LUT6 #(
   .INIT(64'b0000001100110110011100010110111111001011010001001101011111111110)  
) LUT6_1272 (
   .O(gates_1242),
   .I0(InputBits[65]),
   .I1(InputBits[209]),
   .I2(InputBits[339]),
   .I3(InputBits[89]),
   .I4(InputBits[470]),
   .I5(InputBits[221])
);
LUT6 #(
   .INIT(64'b1110011011110011010001101000001001001111001100111010010111011011)  
) LUT6_1273 (
   .O(gates_950),
   .I0(InputBits[342]),
   .I1(InputBits[351]),
   .I2(InputBits[291]),
   .I3(InputBits[280]),
   .I4(InputBits[574]),
   .I5(InputBits[259])
);
LUT6 #(
   .INIT(64'b0001011100011001110110111000101001110010011000010010111110001001)  
) LUT6_1274 (
   .O(gates_887),
   .I0(InputBits[565]),
   .I1(InputBits[401]),
   .I2(InputBits[527]),
   .I3(InputBits[19]),
   .I4(InputBits[11]),
   .I5(InputBits[536])
);
LUT6 #(
   .INIT(64'b1110100011111001000110001111101111100000001111101011101010000100)  
) LUT6_1275 (
   .O(gates_18),
   .I0(InputBits[137]),
   .I1(InputBits[246]),
   .I2(InputBits[220]),
   .I3(InputBits[42]),
   .I4(InputBits[171]),
   .I5(InputBits[17])
);
LUT6 #(
   .INIT(64'b0110001010000001101000111001100010111100001011001011111001100001)  
) LUT6_1276 (
   .O(gates_733),
   .I0(InputBits[139]),
   .I1(InputBits[272]),
   .I2(InputBits[91]),
   .I3(InputBits[128]),
   .I4(InputBits[383]),
   .I5(InputBits[496])
);
LUT6 #(
   .INIT(64'b1010000000111100001101010110010000111111101110110110110100101111)  
) LUT6_1277 (
   .O(gates_1333),
   .I0(InputBits[164]),
   .I1(InputBits[101]),
   .I2(InputBits[193]),
   .I3(InputBits[447]),
   .I4(InputBits[367]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000100001010001001111011110011011011000110101100100101011101111)  
) LUT6_1278 (
   .O(gates_1),
   .I0(InputBits[223]),
   .I1(InputBits[497]),
   .I2(InputBits[144]),
   .I3(InputBits[174]),
   .I4(InputBits[214]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0111111000000110100011000110101010010111100111110011111000111011)  
) LUT6_1279 (
   .O(gates_978),
   .I0(InputBits[554]),
   .I1(InputBits[411]),
   .I2(InputBits[529]),
   .I3(InputBits[570]),
   .I4(InputBits[304]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1011111101111000110100111111000100100100000100001011111101010110)  
) LUT6_1280 (
   .O(gates_563),
   .I0(InputBits[110]),
   .I1(InputBits[392]),
   .I2(InputBits[20]),
   .I3(InputBits[288]),
   .I4(InputBits[552]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1000001011010011111100110110100110101000101111011010101001010101)  
) LUT6_1281 (
   .O(gates_1500),
   .I0(InputBits[349]),
   .I1(InputBits[350]),
   .I2(InputBits[117]),
   .I3(InputBits[41]),
   .I4(InputBits[465]),
   .I5(InputBits[422])
);
LUT6 #(
   .INIT(64'b1111001101011011100010101100100001111010101111011000100100010110)  
) LUT6_1282 (
   .O(gates_1066),
   .I0(InputBits[355]),
   .I1(InputBits[417]),
   .I2(InputBits[479]),
   .I3(InputBits[222]),
   .I4(InputBits[515]),
   .I5(InputBits[428])
);
LUT6 #(
   .INIT(64'b1011111001011111011000001000110000010010111110111011001111100101)  
) LUT6_1283 (
   .O(gates_708),
   .I0(InputBits[181]),
   .I1(InputBits[148]),
   .I2(InputBits[482]),
   .I3(InputBits[205]),
   .I4(InputBits[226]),
   .I5(InputBits[58])
);
LUT6 #(
   .INIT(64'b1100110110111010110101110011001100001110101010010011000011110100)  
) LUT6_1284 (
   .O(gates_908),
   .I0(InputBits[319]),
   .I1(InputBits[429]),
   .I2(InputBits[431]),
   .I3(InputBits[290]),
   .I4(InputBits[487]),
   .I5(InputBits[549])
);
LUT6 #(
   .INIT(64'b0111101110001011111011000111010100111010100110000100000001111100)  
) LUT6_1285 (
   .O(gates_1295),
   .I0(InputBits[356]),
   .I1(InputBits[253]),
   .I2(InputBits[522]),
   .I3(InputBits[427]),
   .I4(InputBits[216]),
   .I5(InputBits[95])
);
LUT6 #(
   .INIT(64'b1110000010100000011011011011000110101010111100100001101101111101)  
) LUT6_1286 (
   .O(gates_500),
   .I0(InputBits[97]),
   .I1(InputBits[154]),
   .I2(InputBits[532]),
   .I3(InputBits[188]),
   .I4(InputBits[88]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1001011011111100001110000000001101011111001110001101111010011010)  
) LUT6_1287 (
   .O(gates_380),
   .I0(InputBits[54]),
   .I1(InputBits[387]),
   .I2(InputBits[152]),
   .I3(InputBits[568]),
   .I4(InputBits[344]),
   .I5(InputBits[44])
);
LUT6 #(
   .INIT(64'b1001001011111011111011100010111101100001100101011001010001100011)  
) LUT6_1288 (
   .O(gates_654),
   .I0(InputBits[514]),
   .I1(InputBits[303]),
   .I2(InputBits[123]),
   .I3(InputBits[175]),
   .I4(InputBits[310]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0000001001110011101011100110110011000111010110010000001111011111)  
) LUT6_1289 (
   .O(gates_243),
   .I0(InputBits[563]),
   .I1(InputBits[519]),
   .I2(InputBits[394]),
   .I3(InputBits[94]),
   .I4(InputBits[359]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0001110000010110100001110010010010101100111011010001110011010101)  
) LUT6_1290 (
   .O(gates_1210),
   .I0(InputBits[443]),
   .I1(InputBits[86]),
   .I2(InputBits[151]),
   .I3(InputBits[10]),
   .I4(InputBits[32]),
   .I5(InputBits[146])
);
LUT6 #(
   .INIT(64'b0101100111100101001111001010010100011101110000110010001001000000)  
) LUT6_1291 (
   .O(gates_900),
   .I0(InputBits[472]),
   .I1(InputBits[468]),
   .I2(InputBits[511]),
   .I3(InputBits[38]),
   .I4(InputBits[60]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1011011111111100111111110111101110111011111110111110010001100001)  
) LUT6_1292 (
   .O(gates_1155),
   .I0(InputBits[210]),
   .I1(InputBits[309]),
   .I2(InputBits[437]),
   .I3(InputBits[418]),
   .I4(InputBits[15]),
   .I5(InputBits[48])
);
LUT6 #(
   .INIT(64'b0110110111101000001111110100110000100010000111000011011011110000)  
) LUT6_1293 (
   .O(gates_700),
   .I0(InputBits[516]),
   .I1(InputBits[509]),
   .I2(InputBits[77]),
   .I3(InputBits[141]),
   .I4(InputBits[393]),
   .I5(InputBits[338])
);
LUT6 #(
   .INIT(64'b1001110011100110110001011000010000000000111011010001000101000001)  
) LUT6_1294 (
   .O(gates_362),
   .I0(InputBits[104]),
   .I1(InputBits[59]),
   .I2(InputBits[498]),
   .I3(InputBits[534]),
   .I4(InputBits[263]),
   .I5(InputBits[576])
);
LUT6 #(
   .INIT(64'b0111100001010101011111111000100101010011010001011101110010101011)  
) LUT6_1295 (
   .O(gates_1190),
   .I0(InputBits[564]),
   .I1(InputBits[160]),
   .I2(InputBits[322]),
   .I3(InputBits[545]),
   .I4(InputBits[159]),
   .I5(InputBits[551])
);
LUT6 #(
   .INIT(64'b1011010010000110000110001100000000001100010010010110011100010111)  
) LUT6_1296 (
   .O(gates_1056),
   .I0(InputBits[215]),
   .I1(InputBits[517]),
   .I2(InputBits[111]),
   .I3(InputBits[39]),
   .I4(InputBits[486]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0010110110010110111100100000001110000001000010111010101011110000)  
) LUT6_1297 (
   .O(gates_1211),
   .I0(gates_297),
   .I1(gates_307),
   .I2(gates_1528),
   .I3(gates_1179),
   .I4(gates_46),
   .I5(gates_819)
);
LUT6 #(
   .INIT(64'b1101101000001101011010111011101011011000011100100011100010100001)  
) LUT6_1298 (
   .O(gates_570),
   .I0(gates_619),
   .I1(gates_1144),
   .I2(gates_948),
   .I3(gates_106),
   .I4(gates_907),
   .I5(gates_1517)
);
LUT6 #(
   .INIT(64'b1101110010111100010101010111110100100010100011101110100010111010)  
) LUT6_1299 (
   .O(gates_128),
   .I0(gates_1470),
   .I1(gates_1415),
   .I2(gates_1397),
   .I3(gates_1378),
   .I4(gates_801),
   .I5(gates_1414)
);
LUT6 #(
   .INIT(64'b0011100101011000110000010001001000000111011010100110001110110001)  
) LUT6_1300 (
   .O(gates_470),
   .I0(gates_1428),
   .I1(gates_1367),
   .I2(gates_341),
   .I3(gates_1530),
   .I4(gates_1463),
   .I5(gates_740)
);
LUT6 #(
   .INIT(64'b1110010111001100011000001001010000001100111100010010110011101010)  
) LUT6_1301 (
   .O(gates_1296),
   .I0(gates_318),
   .I1(gates_960),
   .I2(gates_577),
   .I3(gates_1240),
   .I4(gates_998),
   .I5(gates_1408)
);
LUT6 #(
   .INIT(64'b0010111100111110101111001110010100101010101011111001100001101101)  
) LUT6_1302 (
   .O(gates_1201),
   .I0(gates_964),
   .I1(gates_327),
   .I2(gates_1262),
   .I3(gates_1088),
   .I4(gates_830),
   .I5(gates_449)
);
LUT6 #(
   .INIT(64'b0111100001001001110111111010100101011110110110010110001001110001)  
) LUT6_1303 (
   .O(gates_13),
   .I0(gates_188),
   .I1(gates_202),
   .I2(gates_175),
   .I3(gates_1555),
   .I4(gates_97),
   .I5(gates_1009)
);
LUT6 #(
   .INIT(64'b0110101011000000111001110001000001001110111011010000110101100011)  
) LUT6_1304 (
   .O(gates_820),
   .I0(gates_250),
   .I1(gates_868),
   .I2(gates_1098),
   .I3(gates_1329),
   .I4(gates_1315),
   .I5(gates_293)
);
LUT6 #(
   .INIT(64'b0110100000100111110111001001011011000100000010100100111001110101)  
) LUT6_1305 (
   .O(gates_838),
   .I0(gates_970),
   .I1(gates_817),
   .I2(gates_1418),
   .I3(gates_539),
   .I4(gates_1137),
   .I5(gates_378)
);
LUT6 #(
   .INIT(64'b0011010100000000010011111110011000001100010101111101101000001000)  
) LUT6_1306 (
   .O(gates_1141),
   .I0(gates_747),
   .I1(gates_1152),
   .I2(gates_1343),
   .I3(gates_683),
   .I4(gates_947),
   .I5(gates_637)
);
LUT6 #(
   .INIT(64'b0101101101100000110000100100100110101000001100100011101001000010)  
) LUT6_1307 (
   .O(gates_1079),
   .I0(gates_1545),
   .I1(gates_1158),
   .I2(gates_1122),
   .I3(gates_411),
   .I4(gates_1177),
   .I5(gates_275)
);
LUT6 #(
   .INIT(64'b1100010010011011100010100101111110110011101100100001111000110110)  
) LUT6_1308 (
   .O(gates_1015),
   .I0(gates_980),
   .I1(gates_911),
   .I2(gates_7),
   .I3(gates_593),
   .I4(gates_1146),
   .I5(gates_460)
);
LUT6 #(
   .INIT(64'b1110100010110011000001111100110001110000000111000001111110000111)  
) LUT6_1309 (
   .O(gates_1433),
   .I0(gates_312),
   .I1(gates_549),
   .I2(gates_1149),
   .I3(gates_548),
   .I4(gates_1033),
   .I5(gates_315)
);
LUT6 #(
   .INIT(64'b0111010010100101011001000010100111111101000001001011111000110110)  
) LUT6_1310 (
   .O(gates_753),
   .I0(gates_977),
   .I1(gates_1365),
   .I2(gates_601),
   .I3(gates_1446),
   .I4(gates_617),
   .I5(gates_771)
);
LUT6 #(
   .INIT(64'b1001101000001111101011001011111011000001011101000111101010011011)  
) LUT6_1311 (
   .O(gates_233),
   .I0(gates_1290),
   .I1(gates_30),
   .I2(gates_655),
   .I3(gates_141),
   .I4(gates_459),
   .I5(gates_64)
);
LUT6 #(
   .INIT(64'b0110000100111000000011111001101000111011010010001111001110000011)  
) LUT6_1312 (
   .O(gates_1161),
   .I0(gates_452),
   .I1(gates_57),
   .I2(gates_4),
   .I3(gates_353),
   .I4(gates_8),
   .I5(gates_1362)
);
LUT6 #(
   .INIT(64'b0101010000111010110101101100111100111101111110000001000110111100)  
) LUT6_1313 (
   .O(gates_337),
   .I0(gates_406),
   .I1(gates_1082),
   .I2(gates_1167),
   .I3(gates_567),
   .I4(gates_301),
   .I5(gates_1001)
);
LUT6 #(
   .INIT(64'b1000011101010010100101000011010111000110101011001110101010001111)  
) LUT6_1314 (
   .O(gates_899),
   .I0(gates_381),
   .I1(gates_1221),
   .I2(gates_335),
   .I3(gates_1048),
   .I4(gates_1204),
   .I5(gates_641)
);
LUT6 #(
   .INIT(64'b0101110001010110100010100110111111100010010110010100110111011101)  
) LUT6_1315 (
   .O(gates_1441),
   .I0(gates_1169),
   .I1(gates_1021),
   .I2(gates_1010),
   .I3(gates_69),
   .I4(gates_159),
   .I5(gates_935)
);
LUT6 #(
   .INIT(64'b0001010111011011010010001010101011100101110111110000101000011100)  
) LUT6_1316 (
   .O(gates_754),
   .I0(gates_1159),
   .I1(gates_1368),
   .I2(gates_992),
   .I3(gates_937),
   .I4(gates_1032),
   .I5(gates_455)
);
LUT6 #(
   .INIT(64'b1101010100001001111101011011100100011110111010001011110010001111)  
) LUT6_1317 (
   .O(gates_1030),
   .I0(gates_521),
   .I1(gates_527),
   .I2(gates_432),
   .I3(gates_514),
   .I4(gates_147),
   .I5(gates_922)
);
LUT6 #(
   .INIT(64'b1011101101011110011001010100001101000000011111110111001011110000)  
) LUT6_1318 (
   .O(gates_1263),
   .I0(gates_859),
   .I1(gates_909),
   .I2(gates_916),
   .I3(gates_1244),
   .I4(gates_768),
   .I5(gates_1278)
);
LUT6 #(
   .INIT(64'b0001101111110001001010000000010001011001001101110011110000000001)  
) LUT6_1319 (
   .O(gates_1053),
   .I0(gates_59),
   .I1(gates_725),
   .I2(gates_1350),
   .I3(gates_238),
   .I4(gates_1261),
   .I5(gates_242)
);
LUT6 #(
   .INIT(64'b0010011111111100001001000000110111111110001101000110001000101110)  
) LUT6_1320 (
   .O(gates_925),
   .I0(gates_1482),
   .I1(gates_930),
   .I2(gates_1134),
   .I3(gates_506),
   .I4(gates_79),
   .I5(gates_1464)
);
LUT6 #(
   .INIT(64'b0001100000010011011001110010101001100011001100110101001110011001)  
) LUT6_1321 (
   .O(gates_37),
   .I0(gates_1431),
   .I1(gates_656),
   .I2(gates_1197),
   .I3(gates_393),
   .I4(gates_498),
   .I5(gates_1385)
);
LUT6 #(
   .INIT(64'b1101011010100101010110101101000111000110101111101110111011011100)  
) LUT6_1322 (
   .O(gates_732),
   .I0(gates_444),
   .I1(gates_763),
   .I2(gates_778),
   .I3(gates_524),
   .I4(gates_1136),
   .I5(gates_580)
);
LUT6 #(
   .INIT(64'b0111100111000001001111001001010100000001101001010000110000111110)  
) LUT6_1323 (
   .O(gates_1347),
   .I0(gates_485),
   .I1(gates_636),
   .I2(gates_1388),
   .I3(gates_906),
   .I4(gates_181),
   .I5(gates_757)
);
LUT6 #(
   .INIT(64'b1101100110011101100000001110100011010101110011010010100010000111)  
) LUT6_1324 (
   .O(gates_330),
   .I0(gates_457),
   .I1(gates_1299),
   .I2(gates_1489),
   .I3(gates_1391),
   .I4(gates_1539),
   .I5(gates_581)
);
LUT6 #(
   .INIT(64'b1011110111000111010010000010001001101100111111000000111111101100)  
) LUT6_1325 (
   .O(gates_1148),
   .I0(gates_1436),
   .I1(gates_1379),
   .I2(gates_1027),
   .I3(gates_811),
   .I4(gates_1521),
   .I5(gates_407)
);
LUT6 #(
   .INIT(64'b1100101111000111100110000110110010111111111001010110100011010000)  
) LUT6_1326 (
   .O(gates_774),
   .I0(gates_261),
   .I1(gates_174),
   .I2(gates_1284),
   .I3(gates_1230),
   .I4(gates_1234),
   .I5(gates_372)
);
LUT6 #(
   .INIT(64'b0010000101101100011000010100100101001011101111010111010111010001)  
) LUT6_1327 (
   .O(gates_143),
   .I0(gates_446),
   .I1(gates_673),
   .I2(gates_793),
   .I3(gates_17),
   .I4(gates_1120),
   .I5(gates_788)
);
LUT6 #(
   .INIT(64'b1001001010001101100110100001110000011101011110011001011010001010)  
) LUT6_1328 (
   .O(gates_296),
   .I0(gates_1425),
   .I1(gates_837),
   .I2(gates_724),
   .I3(gates_1324),
   .I4(gates_1387),
   .I5(gates_433)
);
LUT6 #(
   .INIT(64'b0101001100111110100101111111000111011010011101101001100000110001)  
) LUT6_1329 (
   .O(gates_850),
   .I0(gates_928),
   .I1(gates_649),
   .I2(gates_163),
   .I3(gates_728),
   .I4(gates_1228),
   .I5(gates_1335)
);
LUT6 #(
   .INIT(64'b0011110010110001011100110100001000110101101010111100001110110100)  
) LUT6_1330 (
   .O(gates_993),
   .I0(gates_594),
   .I1(gates_183),
   .I2(gates_1044),
   .I3(gates_78),
   .I4(gates_1256),
   .I5(gates_1318)
);
LUT6 #(
   .INIT(64'b1101111010010100111001011001101110011001010001101000001111101111)  
) LUT6_1331 (
   .O(gates_1341),
   .I0(gates_1166),
   .I1(gates_565),
   .I2(gates_699),
   .I3(gates_1178),
   .I4(gates_775),
   .I5(gates_697)
);
LUT6 #(
   .INIT(64'b0111101011011110010010000001110010101011010101101111010010100011)  
) LUT6_1332 (
   .O(gates_591),
   .I0(gates_815),
   .I1(gates_764),
   .I2(gates_688),
   .I3(gates_1493),
   .I4(gates_629),
   .I5(gates_628)
);
LUT6 #(
   .INIT(64'b0110111101101011001001010111101110111000001100111100100100010101)  
) LUT6_1333 (
   .O(gates_386),
   .I0(gates_1481),
   .I1(gates_285),
   .I2(gates_394),
   .I3(gates_1116),
   .I4(gates_1352),
   .I5(gates_612)
);
LUT6 #(
   .INIT(64'b0111100000100111100010111011101110011111111010101111010001001101)  
) LUT6_1334 (
   .O(gates_217),
   .I0(gates_1449),
   .I1(gates_709),
   .I2(gates_1499),
   .I3(gates_1483),
   .I4(gates_831),
   .I5(gates_1488)
);
LUT6 #(
   .INIT(64'b0100110101010100101001001001111111100110011011101010101100010110)  
) LUT6_1335 (
   .O(gates_421),
   .I0(gates_1422),
   .I1(gates_858),
   .I2(gates_1163),
   .I3(gates_23),
   .I4(gates_1515),
   .I5(gates_929)
);
LUT6 #(
   .INIT(64'b0110111100001111110111111100000011011110000101000010100011110010)  
) LUT6_1336 (
   .O(gates_1090),
   .I0(gates_752),
   .I1(gates_475),
   .I2(gates_1496),
   .I3(gates_726),
   .I4(gates_43),
   .I5(gates_1147)
);
LUT6 #(
   .INIT(64'b0100000010001110011101001101000000000111111100100111000011010001)  
) LUT6_1337 (
   .O(gates_547),
   .I0(gates_185),
   .I1(gates_823),
   .I2(gates_1487),
   .I3(gates_468),
   .I4(gates_177),
   .I5(gates_1330)
);
LUT6 #(
   .INIT(64'b0101110111101100101001000001001000100010111101001011010100101101)  
) LUT6_1338 (
   .O(gates_1133),
   .I0(gates_1401),
   .I1(gates_1452),
   .I2(gates_1239),
   .I3(gates_1382),
   .I4(gates_70),
   .I5(gates_219)
);
LUT6 #(
   .INIT(64'b0011100011100011011100100100111110011111010010001001001111010001)  
) LUT6_1339 (
   .O(gates_1223),
   .I0(gates_642),
   .I1(gates_95),
   .I2(gates_1014),
   .I3(gates_533),
   .I4(gates_1506),
   .I5(gates_745)
);
LUT6 #(
   .INIT(64'b1010000001010101100110010100111010011010010001010101010110111110)  
) LUT6_1340 (
   .O(gates_694),
   .I0(gates_324),
   .I1(gates_166),
   .I2(gates_718),
   .I3(gates_1220),
   .I4(gates_1375),
   .I5(gates_543)
);
LUT6 #(
   .INIT(64'b1100000000111000011110011110010110101101011001000101101000000011)  
) LUT6_1341 (
   .O(gates_1435),
   .I0(gates_1316),
   .I1(gates_1052),
   .I2(gates_263),
   .I3(gates_537),
   .I4(gates_622),
   .I5(gates_158)
);
LUT6 #(
   .INIT(64'b1001010110000010110000000111000011001101010011110100001010000110)  
) LUT6_1342 (
   .O(gates_790),
   .I0(gates_927),
   .I1(gates_1064),
   .I2(gates_260),
   .I3(gates_1175),
   .I4(gates_150),
   .I5(gates_1351)
);
LUT6 #(
   .INIT(64'b1111010010111000010010110100100000110001111101110111110110011110)  
) LUT6_1343 (
   .O(gates_760),
   .I0(gates_555),
   .I1(gates_1236),
   .I2(gates_574),
   .I3(gates_1182),
   .I4(gates_963),
   .I5(gates_1491)
);
LUT6 #(
   .INIT(64'b1101101011001110101001010100100100100110011110101110100111100110)  
) LUT6_1344 (
   .O(gates_727),
   .I0(gates_1276),
   .I1(gates_520),
   .I2(gates_735),
   .I3(gates_503),
   .I4(gates_1008),
   .I5(gates_1522)
);
LUT6 #(
   .INIT(64'b0001110000110000110111100110100110001100100101101100111000100011)  
) LUT6_1345 (
   .O(gates_551),
   .I0(gates_891),
   .I1(gates_497),
   .I2(gates_679),
   .I3(gates_784),
   .I4(gates_447),
   .I5(gates_1012)
);
LUT6 #(
   .INIT(64'b0101000101010001001011100100101101101100011110000011100001100111)  
) LUT6_1346 (
   .O(gates_1051),
   .I0(gates_1461),
   .I1(gates_405),
   .I2(gates_1469),
   .I3(gates_779),
   .I4(gates_1125),
   .I5(gates_19)
);
LUT6 #(
   .INIT(64'b0110010101110001010111010001001110001111110101011101111101101000)  
) LUT6_1347 (
   .O(gates_229),
   .I0(gates_1484),
   .I1(gates_1550),
   .I2(gates_442),
   .I3(gates_1078),
   .I4(gates_780),
   .I5(gates_1281)
);
LUT6 #(
   .INIT(64'b0100011101000011110111111010011100001101111011101111110011010110)  
) LUT6_1348 (
   .O(gates_1016),
   .I0(gates_309),
   .I1(gates_923),
   .I2(gates_1536),
   .I3(gates_722),
   .I4(gates_1430),
   .I5(gates_988)
);
LUT6 #(
   .INIT(64'b0010010110100000110001101111010111110111001101001100001111010100)  
) LUT6_1349 (
   .O(gates_982),
   .I0(gates_695),
   .I1(gates_867),
   .I2(gates_995),
   .I3(gates_846),
   .I4(gates_1371),
   .I5(gates_401)
);
LUT6 #(
   .INIT(64'b1101011110000000010100101011010011110001111111000010101110111001)  
) LUT6_1350 (
   .O(gates_395),
   .I0(gates_999),
   .I1(gates_1187),
   .I2(gates_1059),
   .I3(gates_1003),
   .I4(gates_1113),
   .I5(gates_154)
);
LUT6 #(
   .INIT(64'b1010110110101111000000010110100111111110101000100100000011001001)  
) LUT6_1351 (
   .O(gates_487),
   .I0(gates_1444),
   .I1(gates_294),
   .I2(gates_1226),
   .I3(gates_1031),
   .I4(gates_711),
   .I5(gates_65)
);
LUT6 #(
   .INIT(64'b1001111111011100011101001110110001100101100001111101110001011101)  
) LUT6_1352 (
   .O(gates_419),
   .I0(gates_1176),
   .I1(gates_1202),
   .I2(gates_1344),
   .I3(gates_663),
   .I4(gates_1288),
   .I5(gates_873)
);
LUT6 #(
   .INIT(64'b1110100010011001111110010100111011110001011010111110001010100000)  
) LUT6_1353 (
   .O(gates_518),
   .I0(gates_1248),
   .I1(gates_93),
   .I2(gates_634),
   .I3(gates_344),
   .I4(gates_1447),
   .I5(gates_161)
);
LUT6 #(
   .INIT(64'b0001111000101001011000101010111110100011100100010010100001000001)  
) LUT6_1354 (
   .O(gates_795),
   .I0(gates_665),
   .I1(gates_368),
   .I2(gates_1277),
   .I3(gates_379),
   .I4(gates_501),
   .I5(gates_1513)
);
LUT6 #(
   .INIT(64'b1010001001110101110101110110000111000110010101011111011100000000)  
) LUT6_1355 (
   .O(gates_1264),
   .I0(gates_11),
   .I1(gates_208),
   .I2(gates_1337),
   .I3(gates_569),
   .I4(gates_1231),
   .I5(gates_621)
);
LUT6 #(
   .INIT(64'b0000110001001001011011011101000111110100001001111001110110101010)  
) LUT6_1356 (
   .O(gates_945),
   .I0(gates_813),
   .I1(gates_536),
   .I2(gates_616),
   .I3(gates_412),
   .I4(gates_1282),
   .I5(gates_1005)
);
LUT6 #(
   .INIT(64'b1000000100101111000001001000010111111111100010101011011011100100)  
) LUT6_1357 (
   .O(gates_239),
   .I0(gates_640),
   .I1(gates_857),
   .I2(gates_954),
   .I3(gates_1145),
   .I4(gates_1164),
   .I5(gates_72)
);
LUT6 #(
   .INIT(64'b0001000011101111110011001010011100011110101110111100011110101000)  
) LUT6_1358 (
   .O(gates_734),
   .I0(gates_1172),
   .I1(gates_959),
   .I2(gates_967),
   .I3(gates_1395),
   .I4(gates_1404),
   .I5(gates_262)
);
LUT6 #(
   .INIT(64'b1001111100100001111100011011110010110110111001110110111001111000)  
) LUT6_1359 (
   .O(gates_851),
   .I0(gates_860),
   .I1(gates_707),
   .I2(gates_463),
   .I3(gates_917),
   .I4(gates_1541),
   .I5(gates_919)
);
LUT6 #(
   .INIT(64'b1001101111010011000000000111110010001111100011111000111000000000)  
) LUT6_1360 (
   .O(gates_2),
   .I0(gates_1300),
   .I1(gates_1507),
   .I2(gates_291),
   .I3(gates_1336),
   .I4(gates_1523),
   .I5(gates_703)
);
LUT6 #(
   .INIT(64'b1110001000110101001000010111101001101100110000011101000100000011)  
) LUT6_1361 (
   .O(gates_1472),
   .I0(gates_320),
   .I1(gates_1265),
   .I2(gates_1127),
   .I3(gates_646),
   .I4(gates_1474),
   .I5(gates_886)
);
LUT6 #(
   .INIT(64'b0111001111110010111110011000101000010001010011001101000011000001)  
) LUT6_1362 (
   .O(gates_979),
   .I0(gates_1095),
   .I1(gates_3),
   .I2(gates_557),
   .I3(gates_739),
   .I4(gates_1527),
   .I5(gates_659)
);
LUT6 #(
   .INIT(64'b0111111111101101111110101011011001110110010110001011001000100011)  
) LUT6_1363 (
   .O(gates_1373),
   .I0(gates_329),
   .I1(gates_354),
   .I2(gates_1057),
   .I3(gates_897),
   .I4(gates_1062),
   .I5(gates_789)
);
LUT6 #(
   .INIT(64'b0001100001101010011101101010001000000101111111111001101110000111)  
) LUT6_1364 (
   .O(gates_377),
   .I0(gates_1466),
   .I1(gates_544),
   .I2(gates_633),
   .I3(gates_839),
   .I4(gates_560),
   .I5(gates_105)
);
LUT6 #(
   .INIT(64'b1101111010100111010000000001010010010011101001111011110100100110)  
) LUT6_1365 (
   .O(gates_1092),
   .I0(gates_1298),
   .I1(gates_670),
   .I2(gates_731),
   .I3(gates_357),
   .I4(gates_690),
   .I5(gates_102)
);
LUT6 #(
   .INIT(64'b0001100110110110011011110100111101011001010001001100011001011000)  
) LUT6_1366 (
   .O(gates_385),
   .I0(gates_84),
   .I1(gates_647),
   .I2(gates_483),
   .I3(gates_138),
   .I4(gates_1497),
   .I5(gates_441)
);
LUT6 #(
   .INIT(64'b0011001010010101001110011011000000100100101001000101101000110110)  
) LUT6_1367 (
   .O(gates_848),
   .I0(gates_267),
   .I1(gates_350),
   .I2(gates_797),
   .I3(gates_173),
   .I4(gates_568),
   .I5(gates_113)
);
LUT6 #(
   .INIT(64'b1110111000001000100100011010011011001111111001000000100110011101)  
) LUT6_1368 (
   .O(gates_598),
   .I0(gates_597),
   .I1(gates_871),
   .I2(gates_103),
   .I3(gates_6),
   .I4(gates_608),
   .I5(gates_1420)
);
LUT6 #(
   .INIT(64'b0000010100000110001101011011010101101110101100000101100100011110)  
) LUT6_1369 (
   .O(gates_348),
   .I0(gates_1504),
   .I1(gates_1104),
   .I2(gates_228),
   .I3(gates_806),
   .I4(gates_675),
   .I5(gates_599)
);
LUT6 #(
   .INIT(64'b1110000111011000100000001100000110100011101110110001010011000001)  
) LUT6_1370 (
   .O(gates_112),
   .I0(gates_142),
   .I1(gates_1473),
   .I2(gates_802),
   .I3(gates_799),
   .I4(gates_1100),
   .I5(gates_359)
);
LUT6 #(
   .INIT(64'b0100000100011100010110101101001000111110110010001000100100110110)  
) LUT6_1371 (
   .O(gates_1039),
   .I0(gates_426),
   .I1(gates_479),
   .I2(gates_336),
   .I3(gates_717),
   .I4(gates_1101),
   .I5(gates_1546)
);
LUT6 #(
   .INIT(64'b0011011100101000011001101111111011111110111001101000000111100101)  
) LUT6_1372 (
   .O(gates_1348),
   .I0(gates_272),
   .I1(gates_625),
   .I2(gates_1267),
   .I3(gates_721),
   .I4(gates_1069),
   .I5(gates_332)
);
LUT6 #(
   .INIT(64'b0110010110010000100100010000110100110000001101101110010011000011)  
) LUT6_1373 (
   .O(gates_941),
   .I0(gates_1097),
   .I1(gates_1325),
   .I2(gates_504),
   .I3(gates_1198),
   .I4(gates_805),
   .I5(gates_345)
);
LUT6 #(
   .INIT(64'b1011000101101011110110001000101010001010101110110111110100101010)  
) LUT6_1374 (
   .O(gates_117),
   .I0(gates_667),
   .I1(gates_316),
   .I2(gates_1448),
   .I3(gates_1406),
   .I4(gates_1170),
   .I5(gates_415)
);
LUT6 #(
   .INIT(64'b1101000101011000101110011001011110101001011111111110111111011101)  
) LUT6_1375 (
   .O(gates_1309),
   .I0(gates_1106),
   .I1(gates_264),
   .I2(gates_687),
   .I3(gates_614),
   .I4(gates_1355),
   .I5(gates_448)
);
LUT6 #(
   .INIT(64'b0000111010010001001100010011011110111001011111110110100011000100)  
) LUT6_1376 (
   .O(gates_1108),
   .I0(gates_326),
   .I1(gates_118),
   .I2(gates_306),
   .I3(gates_1389),
   .I4(gates_531),
   .I5(gates_638)
);
LUT6 #(
   .INIT(64'b1001110000110010001110111111001111011111011101111000101100111101)  
) LUT6_1377 (
   .O(gates_1512),
   .I0(gates_51),
   .I1(gates_1041),
   .I2(gates_1495),
   .I3(gates_237),
   .I4(gates_825),
   .I5(gates_877)
);
LUT6 #(
   .INIT(64'b1111011100100101111100101101010000101100110101001001010001010001)  
) LUT6_1378 (
   .O(gates_437),
   .I0(gates_912),
   .I1(gates_38),
   .I2(gates_197),
   .I3(gates_639),
   .I4(gates_666),
   .I5(gates_169)
);
LUT6 #(
   .INIT(64'b0011010011101101010101001010000011110011111110001010001101000100)  
) LUT6_1379 (
   .O(gates_1272),
   .I0(gates_1199),
   .I1(gates_592),
   .I2(gates_1372),
   .I3(gates_1099),
   .I4(gates_1255),
   .I5(gates_938)
);
LUT6 #(
   .INIT(64'b1011110101000110101000100000101101101110111101000000010010011011)  
) LUT6_1380 (
   .O(gates_1129),
   .I0(gates_210),
   .I1(gates_1357),
   .I2(gates_1227),
   .I3(gates_289),
   .I4(gates_681),
   .I5(gates_1215)
);
LUT6 #(
   .INIT(64'b0000101110001111010001110011010001000000010110101101111101100011)  
) LUT6_1381 (
   .O(gates_133),
   .I0(gates_477),
   .I1(gates_528),
   .I2(gates_865),
   .I3(gates_630),
   .I4(gates_895),
   .I5(gates_1128)
);
LUT6 #(
   .INIT(64'b1100010001111110000010001010110110010001000010000001101001000111)  
) LUT6_1382 (
   .O(gates_1416),
   .I0(gates_116),
   .I1(gates_1542),
   .I2(gates_1219),
   .I3(gates_400),
   .I4(gates_1364),
   .I5(gates_1055)
);
LUT6 #(
   .INIT(64'b1110101111001111111010100101110100101010101100001001101101100111)  
) LUT6_1383 (
   .O(gates_1400),
   .I0(gates_546),
   .I1(gates_60),
   .I2(gates_429),
   .I3(gates_1253),
   .I4(gates_1434),
   .I5(gates_976)
);
LUT6 #(
   .INIT(64'b1110100011111001111001001001100001111011110000110110100001011001)  
) LUT6_1384 (
   .O(gates_213),
   .I0(gates_677),
   .I1(gates_874),
   .I2(gates_29),
   .I3(gates_1023),
   .I4(gates_63),
   .I5(gates_767)
);
LUT6 #(
   .INIT(64'b1010110010111101011110010011110111011110001101010110111011100101)  
) LUT6_1385 (
   .O(gates_1459),
   .I0(gates_975),
   .I1(gates_456),
   .I2(gates_321),
   .I3(gates_126),
   .I4(gates_466),
   .I5(gates_1140)
);
LUT6 #(
   .INIT(64'b0000111110111111010111100111111100000000111001100011001001001001)  
) LUT6_1386 (
   .O(gates_196),
   .I0(gates_576),
   .I1(gates_61),
   .I2(gates_809),
   .I3(gates_254),
   .I4(gates_875),
   .I5(gates_1063)
);
LUT6 #(
   .INIT(64'b1010101001101100010100110111101001001001100011001100000101111011)  
) LUT6_1387 (
   .O(gates_15),
   .I0(gates_283),
   .I1(gates_1287),
   .I2(gates_710),
   .I3(gates_712),
   .I4(gates_894),
   .I5(gates_1510)
);
LUT6 #(
   .INIT(64'b1000000111000101110100100111001001010001011101011101000100101101)  
) LUT6_1388 (
   .O(gates_1168),
   .I0(gates_1065),
   .I1(gates_1486),
   .I2(gates_1117),
   .I3(gates_1074),
   .I4(gates_792),
   .I5(gates_785)
);
LUT6 #(
   .INIT(64'b1101100110100101001000001000100001100101110001110100000110011001)  
) LUT6_1389 (
   .O(gates_525),
   .I0(gates_340),
   .I1(gates_879),
   .I2(gates_1121),
   .I3(gates_1135),
   .I4(gates_402),
   .I5(gates_1292)
);
LUT6 #(
   .INIT(64'b1000000010000011000001001000011001111011100001100110110111010110)  
) LUT6_1390 (
   .O(gates_1327),
   .I0(gates_346),
   .I1(gates_200),
   .I2(gates_472),
   .I3(gates_417),
   .I4(gates_1080),
   .I5(gates_510)
);
LUT6 #(
   .INIT(64'b0001000011000100011010100101010100101010011110010111111110010111)  
) LUT6_1391 (
   .O(gates_952),
   .I0(gates_564),
   .I1(gates_1084),
   .I2(gates_686),
   .I3(gates_486),
   .I4(gates_1180),
   .I5(gates_553)
);
LUT6 #(
   .INIT(64'b0111100000110011001110100000010100010100100010001010111100010100)  
) LUT6_1392 (
   .O(gates_1307),
   .I0(gates_1537),
   .I1(gates_435),
   .I2(gates_1285),
   .I3(gates_1390),
   .I4(gates_632),
   .I5(gates_719)
);
LUT6 #(
   .INIT(64'b0101100001110000111111101111101001101000101110110001100100001011)  
) LUT6_1393 (
   .O(gates_969),
   .I0(gates_1529),
   .I1(gates_1413),
   .I2(gates_866),
   .I3(gates_824),
   .I4(gates_812),
   .I5(gates_80)
);
LUT6 #(
   .INIT(64'b1111010101100111001000101100001000111110101100101101001010011110)  
) LUT6_1394 (
   .O(gates_203),
   .I0(gates_1247),
   .I1(gates_266),
   .I2(gates_155),
   .I3(gates_74),
   .I4(gates_883),
   .I5(gates_221)
);
LUT6 #(
   .INIT(64'b1011011001110000000001010100111010100101011101010011011111010110)  
) LUT6_1395 (
   .O(gates_172),
   .I0(gates_1310),
   .I1(gates_278),
   .I2(gates_589),
   .I3(gates_1118),
   .I4(gates_782),
   .I5(gates_438)
);
LUT6 #(
   .INIT(64'b1010101111101001010111011000001101101001110001110110111010110110)  
) LUT6_1396 (
   .O(gates_473),
   .I0(gates_89),
   .I1(gates_25),
   .I2(gates_1131),
   .I3(gates_684),
   .I4(gates_985),
   .I5(gates_882)
);
LUT6 #(
   .INIT(64'b1000100000000100011000011000001001110110100000000000100010101100)  
) LUT6_1397 (
   .O(gates_66),
   .I0(gates_136),
   .I1(gates_295),
   .I2(gates_171),
   .I3(gates_465),
   .I4(gates_669),
   .I5(gates_199)
);
LUT6 #(
   .INIT(64'b0101111010101110010100011001011101111101011100100110100001011011)  
) LUT6_1398 (
   .O(gates_270),
   .I0(gates_840),
   .I1(gates_10),
   .I2(gates_204),
   .I3(gates_1369),
   .I4(gates_1000),
   .I5(gates_698)
);
LUT6 #(
   .INIT(64'b1010010110110000100110011001100111001100001000000011000101010111)  
) LUT6_1399 (
   .O(gates_720),
   .I0(gates_1139),
   .I1(gates_723),
   .I2(gates_781),
   .I3(gates_1323),
   .I4(gates_1342),
   .I5(gates_1002)
);
LUT6 #(
   .INIT(64'b0001000010000111011010011100001110001011101111101010010000010011)  
) LUT6_1400 (
   .O(gates_756),
   .I0(gates_370),
   .I1(gates_885),
   .I2(gates_814),
   .I3(gates_365),
   .I4(gates_1308),
   .I5(gates_578)
);
LUT6 #(
   .INIT(64'b1111010111000110100001111100110011011001010101010110100000010111)  
) LUT6_1401 (
   .O(gates_439),
   .I0(gates_157),
   .I1(gates_281),
   .I2(gates_855),
   .I3(gates_1188),
   .I4(gates_1260),
   .I5(gates_1076)
);
LUT6 #(
   .INIT(64'b0111100000011111101111001100000010001111001100001001111110001110)  
) LUT6_1402 (
   .O(gates_1534),
   .I0(gates_1458),
   .I1(gates_744),
   .I2(gates_436),
   .I3(gates_249),
   .I4(gates_144),
   .I5(gates_870)
);
LUT6 #(
   .INIT(64'b1110000010100010101010101011100001110111100100010110101010100001)  
) LUT6_1403 (
   .O(gates_1093),
   .I0(gates_822),
   .I1(gates_1360),
   .I2(gates_1028),
   .I3(gates_635),
   .I4(gates_268),
   .I5(gates_1543)
);
LUT6 #(
   .INIT(64'b0000000101000101001000111101001100001111100011100100000011000000)  
) LUT6_1404 (
   .O(gates_1233),
   .I0(gates_205),
   .I1(gates_360),
   .I2(gates_55),
   .I3(gates_273),
   .I4(gates_1303),
   .I5(gates_1006)
);
LUT6 #(
   .INIT(64'b0000110110111000011101110000101011101111011001010010101010010110)  
) LUT6_1405 (
   .O(gates_371),
   .I0(gates_1036),
   .I1(gates_1025),
   .I2(gates_1346),
   .I3(gates_1383),
   .I4(gates_997),
   .I5(gates_668)
);
LUT6 #(
   .INIT(64'b0100101110011000100011000010110001100000110100010110100101011100)  
) LUT6_1406 (
   .O(gates_1119),
   .I0(gates_349),
   .I1(gates_482),
   .I2(gates_494),
   .I3(gates_1142),
   .I4(gates_1271),
   .I5(gates_253)
);
LUT6 #(
   .INIT(64'b1000010011010100011111010100110101001110011000010010010101100110)  
) LUT6_1407 (
   .O(gates_1485),
   .I0(gates_821),
   .I1(gates_1061),
   .I2(gates_109),
   .I3(gates_206),
   .I4(gates_716),
   .I5(gates_1274)
);
LUT6 #(
   .INIT(64'b0111011100010100010100011101000111100110001010011110100001011010)  
) LUT6_1408 (
   .O(gates_958),
   .I0(gates_88),
   .I1(gates_696),
   .I2(gates_787),
   .I3(gates_1454),
   .I4(gates_1195),
   .I5(gates_383)
);
LUT6 #(
   .INIT(64'b0101101001110111011001100111000001111110100001001000100110111100)  
) LUT6_1409 (
   .O(gates_1381),
   .I0(gates_458),
   .I1(gates_111),
   .I2(gates_1011),
   .I3(gates_192),
   .I4(gates_994),
   .I5(gates_876)
);
LUT6 #(
   .INIT(64'b1000100111010001010100010001100110000100000000111001111111101001)  
) LUT6_1410 (
   .O(gates_507),
   .I0(gates_689),
   .I1(gates_990),
   .I2(gates_924),
   .I3(gates_1302),
   .I4(gates_445),
   .I5(gates_286)
);
LUT6 #(
   .INIT(64'b0101110111111100110111110111101001101000100000011000100101011110)  
) LUT6_1411 (
   .O(gates_962),
   .I0(gates_1174),
   .I1(gates_863),
   .I2(gates_1126),
   .I3(gates_404),
   .I4(gates_376),
   .I5(gates_1114)
);
LUT6 #(
   .INIT(64'b1111101101111001000000011001100101000010110001010111001001000010)  
) LUT6_1412 (
   .O(gates_816),
   .I0(gates_953),
   .I1(gates_905),
   .I2(gates_1519),
   .I3(gates_949),
   .I4(gates_852),
   .I5(gates_762)
);
LUT6 #(
   .INIT(64'b1000101111000001101111000001110111110011011010011110011100011110)  
) LUT6_1413 (
   .O(gates_1411),
   .I0(gates_333),
   .I1(gates_481),
   .I2(gates_572),
   .I3(gates_310),
   .I4(gates_508),
   .I5(gates_1229)
);
LUT6 #(
   .INIT(64'b1010100010010110010011000111111111001010010100111000100111100010)  
) LUT6_1414 (
   .O(gates_288),
   .I0(gates_478),
   .I1(gates_418),
   .I2(gates_186),
   .I3(gates_1394),
   .I4(gates_148),
   .I5(gates_1191)
);
LUT6 #(
   .INIT(64'b1110010111101000100010100110011101100111001000100111110111011110)  
) LUT6_1415 (
   .O(gates_428),
   .I0(gates_1419),
   .I1(gates_434),
   .I2(gates_1450),
   .I3(gates_991),
   .I4(gates_931),
   .I5(gates_1094)
);
LUT6 #(
   .INIT(64'b0000111001110101010111100001100011111011110101100111001100011010)  
) LUT6_1416 (
   .O(gates_1047),
   .I0(gates_1034),
   .I1(gates_187),
   .I2(gates_783),
   .I3(gates_127),
   .I4(gates_1465),
   .I5(gates_382)
);
LUT6 #(
   .INIT(64'b1001011100101101100111000100001100001010000000000001110011000111)  
) LUT6_1417 (
   .O(gates_1243),
   .I0(gates_339),
   .I1(gates_904),
   .I2(gates_1270),
   .I3(gates_416),
   .I4(gates_913),
   .I5(gates_36)
);
LUT6 #(
   .INIT(64'b0101110000010111011011111110000100001101100000000011000010110010)  
) LUT6_1418 (
   .O(gates_513),
   .I0(gates_692),
   .I1(gates_631),
   .I2(gates_1279),
   .I3(gates_881),
   .I4(gates_1123),
   .I5(gates_535)
);
LUT6 #(
   .INIT(64'b1011100111011001001101011000001001001110011000011010100011100000)  
) LUT6_1419 (
   .O(gates_179),
   .I0(gates_1250),
   .I1(gates_67),
   .I2(gates_1492),
   .I3(gates_550),
   .I4(gates_880),
   .I5(gates_1259)
);
LUT6 #(
   .INIT(64'b0000110000000101101111011100111010101110101011101111011010100000)  
) LUT6_1420 (
   .O(gates_201),
   .I0(gates_230),
   .I1(gates_623),
   .I2(gates_1338),
   .I3(gates_178),
   .I4(gates_108),
   .I5(gates_135)
);
LUT6 #(
   .INIT(64'b0001000000001001111111000101111001011000101101001010001010000110)  
) LUT6_1421 (
   .O(gates_1222),
   .I0(gates_220),
   .I1(gates_1019),
   .I2(gates_743),
   .I3(gates_1471),
   .I4(gates_604),
   .I5(gates_440)
);
LUT6 #(
   .INIT(64'b1100011000001100101100010110111111110111010101001110000001000110)  
) LUT6_1422 (
   .O(gates_983),
   .I0(gates_342),
   .I1(gates_749),
   .I2(gates_1509),
   .I3(gates_1212),
   .I4(gates_391),
   .I5(gates_484)
);
LUT6 #(
   .INIT(64'b0100111000101111010110000001110100001100110101011011001110000001)  
) LUT6_1423 (
   .O(gates_1060),
   .I0(gates_738),
   .I1(gates_45),
   .I2(gates_1045),
   .I3(gates_92),
   .I4(gates_189),
   .I5(gates_942)
);
LUT6 #(
   .INIT(64'b1111110111000111010010001100001101010110010101000011110010111010)  
) LUT6_1424 (
   .O(gates_1354),
   .I0(gates_955),
   .I1(gates_1112),
   .I2(gates_1200),
   .I3(gates_1046),
   .I4(gates_1181),
   .I5(gates_562)
);
LUT6 #(
   .INIT(64'b1010110100110010001001110110001010110100001110101000001111111100)  
) LUT6_1425 (
   .O(gates_1038),
   .I0(gates_245),
   .I1(gates_509),
   .I2(gates_556),
   .I3(gates_661),
   .I4(gates_369),
   .I5(gates_1102)
);
LUT6 #(
   .INIT(64'b0000011011111101011100100100101011110000101010010100000111100000)  
) LUT6_1426 (
   .O(gates_624),
   .I0(gates_375),
   .I1(gates_454),
   .I2(gates_137),
   .I3(gates_984),
   .I4(gates_311),
   .I5(gates_1505)
);
LUT6 #(
   .INIT(64'b1100111111100110111010000110011010000000001101010001000000100111)  
) LUT6_1427 (
   .O(gates_323),
   .I0(gates_76),
   .I1(gates_611),
   .I2(gates_1502),
   .I3(gates_1258),
   .I4(gates_1157),
   .I5(gates_1460)
);
LUT6 #(
   .INIT(64'b0110000111110111101101000100100100010011001011011101010101100010)  
) LUT6_1428 (
   .O(gates_292),
   .I0(gates_1358),
   .I1(gates_1073),
   .I2(gates_888),
   .I3(gates_1462),
   .I4(gates_1374),
   .I5(gates_715)
);
LUT6 #(
   .INIT(64'b1101000101111101110011101111100101011101100100011001000100101000)  
) LUT6_1429 (
   .O(gates_704),
   .I0(gates_32),
   .I1(gates_588),
   .I2(gates_1205),
   .I3(gates_1410),
   .I4(gates_119),
   .I5(gates_1218)
);
LUT6 #(
   .INIT(64'b0011101101100011011111011010010001001011111010111100011001010001)  
) LUT6_1430 (
   .O(gates_223),
   .I0(gates_672),
   .I1(gates_31),
   .I2(gates_773),
   .I3(gates_1232),
   .I4(gates_198),
   .I5(gates_796)
);
LUT6 #(
   .INIT(64'b1001000001111010101001101010010011010100111011100001001101010010)  
) LUT6_1431 (
   .O(gates_247),
   .I0(gates_1525),
   .I1(gates_1349),
   .I2(gates_833),
   .I3(gates_901),
   .I4(gates_844),
   .I5(gates_1111)
);
LUT6 #(
   .INIT(64'b0000011000110011100010010000000000011101010000110010001011111100)  
) LUT6_1432 (
   .O(gates_936),
   .I0(gates_854),
   .I1(gates_1442),
   .I2(gates_519),
   .I3(gates_644),
   .I4(gates_618),
   .I5(gates_363)
);
LUT6 #(
   .INIT(64'b0110011001011100100000011000101111001001011100101001100011011011)  
) LUT6_1433 (
   .O(gates_162),
   .I0(gates_241),
   .I1(gates_853),
   .I2(gates_769),
   .I3(gates_471),
   .I4(gates_1096),
   .I5(gates_44)
);
LUT6 #(
   .INIT(64'b1001100010010110011110010001011001100100010001011001110000011010)  
) LUT6_1434 (
   .O(gates_1154),
   .I0(gates_849),
   .I1(gates_1138),
   .I2(gates_603),
   .I3(gates_1007),
   .I4(gates_1313),
   .I5(gates_1185)
);
LUT6 #(
   .INIT(64'b0000101101110000010000001001010101110101010111011111010011001000)  
) LUT6_1435 (
   .O(gates_1289),
   .I0(gates_602),
   .I1(gates_934),
   .I2(gates_1035),
   .I3(gates_1514),
   .I4(gates_660),
   .I5(gates_280)
);
LUT6 #(
   .INIT(64'b0111010000000111000111000001101010001101100011001101111000100000)  
) LUT6_1436 (
   .O(gates_1018),
   .I0(gates_190),
   .I1(gates_164),
   .I2(gates_1475),
   .I3(gates_643),
   .I4(gates_298),
   .I5(gates_1377)
);
LUT6 #(
   .INIT(64'b0011111101110101000001001100101110111000101010100100010000011010)  
) LUT6_1437 (
   .O(gates_68),
   .I0(gates_579),
   .I1(gates_1249),
   .I2(gates_1203),
   .I3(gates_706),
   .I4(gates_605),
   .I5(gates_1467)
);
LUT6 #(
   .INIT(64'b0010100101010000110100010111111110011011000010001101010010001011)  
) LUT6_1438 (
   .O(gates_1050),
   .I0(gates_1451),
   .I1(gates_810),
   .I2(gates_21),
   .I3(gates_1380),
   .I4(gates_1058),
   .I5(gates_343)
);
LUT6 #(
   .INIT(64'b0110101110011111010101000011000101111110001010010001110110011000)  
) LUT6_1439 (
   .O(gates_512),
   .I0(gates_583),
   .I1(gates_1105),
   .I2(gates_986),
   .I3(gates_226),
   .I4(gates_575),
   .I5(gates_52)
);
LUT6 #(
   .INIT(64'b0110111001101100110111111010110010101010100110001001001000011001)  
) LUT6_1440 (
   .O(gates_755),
   .I0(gates_1087),
   .I1(gates_48),
   .I2(gates_258),
   .I3(gates_693),
   .I4(gates_1407),
   .I5(gates_98)
);
LUT6 #(
   .INIT(64'b0001000110101000000100001100110101111111011011011010001011000111)  
) LUT6_1441 (
   .O(gates_973),
   .I0(gates_211),
   .I1(gates_750),
   .I2(gates_322),
   .I3(gates_915),
   .I4(gates_20),
   .I5(gates_1345)
);
LUT6 #(
   .INIT(64'b1110101000000110010000110000001101100100010110101011111101101010)  
) LUT6_1442 (
   .O(gates_651),
   .I0(gates_502),
   .I1(gates_1083),
   .I2(gates_304),
   .I3(gates_276),
   .I4(gates_246),
   .I5(gates_1207)
);
LUT6 #(
   .INIT(64'b1100111100011101010101100110010001001110110110000011011101110111)  
) LUT6_1443 (
   .O(gates_1206),
   .I0(gates_170),
   .I1(gates_85),
   .I2(gates_1068),
   .I3(gates_290),
   .I4(gates_1213),
   .I5(gates_409)
);
LUT6 #(
   .INIT(64'b0010101100110110101011101101111000111011100011000011010011110010)  
) LUT6_1444 (
   .O(gates_450),
   .I0(gates_338),
   .I1(gates_981),
   .I2(gates_26),
   .I3(gates_86),
   .I4(gates_664),
   .I5(gates_1535)
);
LUT6 #(
   .INIT(64'b1110100110111100110000111100110110011111001000111101000001110000)  
) LUT6_1445 (
   .O(gates_1437),
   .I0(gates_1359),
   .I1(gates_1405),
   .I2(gates_1457),
   .I3(gates_1269),
   .I4(gates_22),
   .I5(gates_351)
);
LUT6 #(
   .INIT(64'b0110010100000111111001111100011111101101000100101000111100111101)  
) LUT6_1446 (
   .O(gates_1540),
   .I0(gates_1403),
   .I1(gates_1275),
   .I2(gates_974),
   .I3(gates_1165),
   .I4(gates_1266),
   .I5(gates_832)
);
LUT6 #(
   .INIT(64'b0101000010011111110011110111100000011111001100010110010101010111)  
) LUT6_1447 (
   .O(gates_847),
   .I0(gates_1402),
   .I1(gates_705),
   .I2(gates_702),
   .I3(gates_134),
   .I4(gates_81),
   .I5(gates_1538)
);
LUT6 #(
   .INIT(64'b1010000111100001011010100110100000101011101111110000010100111100)  
) LUT6_1448 (
   .O(gates_1214),
   .I0(gates_951),
   .I1(gates_554),
   .I2(gates_1017),
   .I3(gates_884),
   .I4(gates_384),
   .I5(gates_515)
);
LUT6 #(
   .INIT(64'b1001110000001010111101100001110110110011010110000101001111011111)  
) LUT6_1449 (
   .O(gates_1115),
   .I0(gates_24),
   .I1(gates_1071),
   .I2(gates_517),
   .I3(gates_573),
   .I4(gates_737),
   .I5(gates_1319)
);
LUT6 #(
   .INIT(64'b1011100110000011001010111000010101101111101000001100001100001101)  
) LUT6_1450 (
   .O(gates_62),
   .I0(gates_12),
   .I1(gates_1208),
   .I2(gates_244),
   .I3(gates_39),
   .I4(gates_671),
   .I5(gates_1376)
);
LUT6 #(
   .INIT(64'b1110100111100000000000111001110000101010100111011001101011000000)  
) LUT6_1451 (
   .O(gates_1417),
   .I0(gates_130),
   .I1(gates_83),
   .I2(gates_499),
   .I3(gates_759),
   .I4(gates_818),
   .I5(gates_1520)
);
LUT6 #(
   .INIT(64'b1000111011000010100110001001010010010010111100100010000001101000)  
) LUT6_1452 (
   .O(gates_932),
   .I0(gates_287),
   .I1(gates_505),
   .I2(gates_751),
   .I3(gates_1494),
   .I4(gates_496),
   .I5(gates_1524)
);
LUT6 #(
   .INIT(64'b1000101000111000110010001001111001000001010110011011011111000110)  
) LUT6_1453 (
   .O(gates_772),
   .I0(gates_1427),
   .I1(gates_305),
   .I2(gates_1189),
   .I3(gates_1477),
   .I4(gates_180),
   .I5(gates_662)
);
LUT6 #(
   .INIT(64'b1101111001010101101110010100111111000011110011100110001001000100)  
) LUT6_1454 (
   .O(gates_1353),
   .I0(gates_168),
   .I1(gates_1554),
   .I2(gates_282),
   .I3(gates_397),
   .I4(gates_325),
   .I5(gates_355)
);
LUT6 #(
   .INIT(64'b0000011111011101101100011110001111100110000101000101111011000011)  
) LUT6_1455 (
   .O(gates_713),
   .I0(gates_1480),
   .I1(gates_274),
   .I2(gates_1432),
   .I3(gates_940),
   .I4(gates_492),
   .I5(gates_1322)
);
LUT6 #(
   .INIT(64'b1100110100101010101100101110111101011011111101101111011110111101)  
) LUT6_1456 (
   .O(gates_1160),
   .I0(gates_957),
   .I1(gates_1238),
   .I2(gates_331),
   .I3(gates_758),
   .I4(gates_748),
   .I5(gates_889)
);
LUT6 #(
   .INIT(64'b1100111011100000101100011100100101110001100011001010011110000111)  
) LUT6_1457 (
   .O(gates_271),
   .I0(gates_191),
   .I1(gates_1334),
   .I2(gates_1085),
   .I3(gates_566),
   .I4(gates_872),
   .I5(gates_965)
);
LUT6 #(
   .INIT(64'b1001101001100001001101001010001101000111011110110000100100011100)  
) LUT6_1458 (
   .O(gates_392),
   .I0(gates_836),
   .I1(gates_1173),
   .I2(gates_626),
   .I3(gates_893),
   .I4(gates_1399),
   .I5(gates_1192)
);
LUT6 #(
   .INIT(64'b1100110101101010010100111010101001110111111101000001100100100000)  
) LUT6_1459 (
   .O(gates_279),
   .I0(gates_413),
   .I1(gates_399),
   .I2(gates_1532),
   .I3(gates_584),
   .I4(gates_896),
   .I5(gates_798)
);
LUT6 #(
   .INIT(64'b0001010010011110001001111100110111011111001110000001100001101010)  
) LUT6_1460 (
   .O(gates_35),
   .I0(gates_1366),
   .I1(gates_16),
   .I2(gates_1013),
   .I3(gates_613),
   .I4(gates_1081),
   .I5(gates_1443)
);
LUT6 #(
   .INIT(64'b0010101111111011010100001110101001000101100000001110101100101111)  
) LUT6_1461 (
   .O(gates_729),
   .I0(gates_890),
   .I1(gates_131),
   .I2(gates_691),
   .I3(gates_1476),
   .I4(gates_54),
   .I5(gates_862)
);
LUT6 #(
   .INIT(64'b1111010011000111000101000000100011001001111110000000101001100111)  
) LUT6_1462 (
   .O(gates_87),
   .I0(gates_777),
   .I1(gates_1547),
   .I2(gates_1241),
   .I3(gates_453),
   .I4(gates_944),
   .I5(gates_730)
);
LUT6 #(
   .INIT(64'b0010011100101111000000010010100011000011010101111011110000111011)  
) LUT6_1463 (
   .O(gates_251),
   .I0(gates_414),
   .I1(gates_523),
   .I2(gates_920),
   .I3(gates_1305),
   .I4(gates_1456),
   .I5(gates_1040)
);
LUT6 #(
   .INIT(64'b0001000011100010111000110000111011010011001010000111111110010111)  
) LUT6_1464 (
   .O(gates_1286),
   .I0(gates_1424),
   .I1(gates_474),
   .I2(gates_252),
   .I3(gates_1301),
   .I4(gates_1217),
   .I5(gates_145)
);
LUT6 #(
   .INIT(64'b1011110010101011001100100101000000110111111100101111101100110110)  
) LUT6_1465 (
   .O(gates_27),
   .I0(gates_235),
   .I1(gates_648),
   .I2(gates_609),
   .I3(gates_259),
   .I4(gates_1151),
   .I5(gates_534)
);
LUT6 #(
   .INIT(64'b1010011101110100011011010011110110110011111111111100100101101100)  
) LUT6_1466 (
   .O(gates_99),
   .I0(gates_1075),
   .I1(gates_966),
   .I2(gates_256),
   .I3(gates_490),
   .I4(gates_1439),
   .I5(gates_1143)
);
LUT6 #(
   .INIT(64'b0110100011011101000001100100101001101010000000011000111100000110)  
) LUT6_1467 (
   .O(gates_1548),
   .I0(gates_195),
   .I1(gates_431),
   .I2(gates_366),
   .I3(gates_308),
   .I4(gates_803),
   .I5(gates_358)
);
LUT6 #(
   .INIT(64'b0000011000111101000111111000001011110111110000110010011101100000)  
) LUT6_1468 (
   .O(gates_9),
   .I0(gates_1518),
   .I1(gates_222),
   .I2(gates_184),
   .I3(gates_114),
   .I4(gates_714),
   .I5(gates_425)
);
LUT6 #(
   .INIT(64'b0000110101000000001100001111110110011111001111000111101011001100)  
) LUT6_1469 (
   .O(gates_1340),
   .I0(gates_480),
   .I1(gates_827),
   .I2(gates_1225),
   .I3(gates_615),
   .I4(gates_90),
   .I5(gates_1026)
);
LUT6 #(
   .INIT(64'b0001100000101101001011111101110010010010011010111000101011101100)  
) LUT6_1470 (
   .O(gates_56),
   .I0(gates_971),
   .I1(gates_302),
   .I2(gates_115),
   .I3(gates_804),
   .I4(gates_1440),
   .I5(gates_469)
);
LUT6 #(
   .INIT(64'b0101111000101000111010001100111111010111011001001000100011100111)  
) LUT6_1471 (
   .O(gates_972),
   .I0(gates_284),
   .I1(gates_600),
   .I2(gates_530),
   .I3(gates_1363),
   .I4(gates_1246),
   .I5(gates_1511)
);
LUT6 #(
   .INIT(64'b1010111101001100011011111000010011100000011000011101011011100110)  
) LUT6_1472 (
   .O(gates_1503),
   .I0(gates_462),
   .I1(gates_800),
   .I2(gates_193),
   .I3(gates_165),
   .I4(gates_34),
   .I5(gates_770)
);
LUT6 #(
   .INIT(64'b0000101011111001000011010111011100111101010110010010101101000000)  
) LUT6_1473 (
   .O(gates_427),
   .I0(gates_1478),
   .I1(gates_989),
   .I2(gates_869),
   .I3(gates_653),
   .I4(gates_1054),
   .I5(gates_585)
);
LUT6 #(
   .INIT(64'b0110111111111011101100011111010110110100100100100111111111111100)  
) LUT6_1474 (
   .O(gates_71),
   .I0(gates_657),
   .I1(gates_1245),
   .I2(gates_645),
   .I3(gates_650),
   .I4(gates_842),
   .I5(gates_1331)
);
LUT6 #(
   .INIT(64'b0110101100101100000101111100101011111111011110011100011100111100)  
) LUT6_1475 (
   .O(gates_516),
   .I0(gates_898),
   .I1(gates_1049),
   .I2(gates_678),
   .I3(gates_1386),
   .I4(gates_167),
   .I5(gates_464)
);
LUT6 #(
   .INIT(64'b1100011111100100101011110100100110000100111000111101000000001110)  
) LUT6_1476 (
   .O(gates_968),
   .I0(gates_1022),
   .I1(gates_1370),
   .I2(gates_387),
   .I3(gates_652),
   .I4(gates_845),
   .I5(gates_538)
);
LUT6 #(
   .INIT(64'b1010001110001110011110011110100110001010100000000010000010001001)  
) LUT6_1477 (
   .O(gates_476),
   .I0(gates_1273),
   .I1(gates_1479),
   .I2(gates_47),
   .I3(gates_1086),
   .I4(gates_1251),
   .I5(gates_864)
);
LUT6 #(
   .INIT(64'b0101101110000111100110111111111001011110011110111100010011101111)  
) LUT6_1478 (
   .O(gates_33),
   .I0(gates_1423),
   .I1(gates_1162),
   .I2(gates_761),
   .I3(gates_430),
   .I4(gates_741),
   .I5(gates_685)
);
LUT6 #(
   .INIT(64'b1001000010111111011111010010001110001000110111100000001110010010)  
) LUT6_1479 (
   .O(gates_1037),
   .I0(gates_529),
   .I1(gates_334),
   .I2(gates_1297),
   .I3(gates_94),
   .I4(gates_540),
   .I5(gates_1067)
);
LUT6 #(
   .INIT(64'b0100011100011000000110100001010110100010001011100101010100111010)  
) LUT6_1480 (
   .O(gates_388),
   .I0(gates_403),
   .I1(gates_1184),
   .I2(gates_467),
   .I3(gates_1501),
   .I4(gates_590),
   .I5(gates_794)
);
LUT6 #(
   .INIT(64'b0110011110111110000101010111011101001111010000101011000101011100)  
) LUT6_1481 (
   .O(gates_1130),
   .I0(gates_558),
   .I1(gates_28),
   .I2(gates_526),
   .I3(gates_1257),
   .I4(gates_152),
   .I5(gates_1183)
);
LUT6 #(
   .INIT(64'b0010101111000100110010110010110001110010111101011111101101001111)  
) LUT6_1482 (
   .O(gates_1311),
   .I0(gates_834),
   .I1(gates_461),
   .I2(gates_146),
   .I3(gates_1043),
   .I4(gates_1293),
   .I5(gates_422)
);
LUT6 #(
   .INIT(64'b0110101001101100011010011110011010110111001101010001100111100110)  
) LUT6_1483 (
   .O(gates_996),
   .I0(gates_1356),
   .I1(gates_918),
   .I2(gates_587),
   .I3(gates_545),
   .I4(gates_1339),
   .I5(gates_1029)
);
LUT6 #(
   .INIT(64'b0101000000110010010010100010101110101110111101000100110100000000)  
) LUT6_1484 (
   .O(gates_1552),
   .I0(gates_319),
   .I1(gates_1254),
   .I2(gates_1455),
   .I3(gates_14),
   .I4(gates_231),
   .I5(gates_91)
);
LUT6 #(
   .INIT(64'b0101001000101110011011001011101101000010011000010100100111011100)  
) LUT6_1485 (
   .O(gates_1326),
   .I0(gates_248),
   .I1(gates_1304),
   .I2(gates_53),
   .I3(gates_75),
   .I4(gates_389),
   .I5(gates_125)
);
LUT6 #(
   .INIT(64'b1101110110000111110111011111110011011101011011101011010111101011)  
) LUT6_1486 (
   .O(gates_352),
   .I0(gates_1549),
   .I1(gates_390),
   .I2(gates_1328),
   .I3(gates_77),
   .I4(gates_265),
   .I5(gates_511)
);
LUT6 #(
   .INIT(64'b1110101111111111011011110000001010000000010101110000100101110100)  
) LUT6_1487 (
   .O(gates_701),
   .I0(gates_742),
   .I1(gates_424),
   .I2(gates_50),
   .I3(gates_123),
   .I4(gates_1091),
   .I5(gates_124)
);
LUT6 #(
   .INIT(64'b1011111000101111010000001011110010110010011001100011001110001101)  
) LUT6_1488 (
   .O(gates_674),
   .I0(gates_234),
   .I1(gates_571),
   .I2(gates_1312),
   .I3(gates_1153),
   .I4(gates_1393),
   .I5(gates_347)
);
LUT6 #(
   .INIT(64'b0010001101010111111101100001001001011111001100000001001100001111)  
) LUT6_1489 (
   .O(gates_240),
   .I0(gates_182),
   .I1(gates_1490),
   .I2(gates_209),
   .I3(gates_878),
   .I4(gates_606),
   .I5(gates_607)
);
LUT6 #(
   .INIT(64'b1000101101000101100001011000010011001011110000110011010001100110)  
) LUT6_1490 (
   .O(gates_987),
   .I0(gates_317),
   .I1(gates_1438),
   .I2(gates_582),
   .I3(gates_658),
   .I4(gates_207),
   .I5(gates_1306)
);
LUT6 #(
   .INIT(64'b1011101011110111011000000001001000010110110100010110100010110011)  
) LUT6_1491 (
   .O(gates_1020),
   .I0(gates_1209),
   .I1(gates_776),
   .I2(gates_1453),
   .I3(gates_541),
   .I4(gates_1280),
   .I5(gates_786)
);
LUT6 #(
   .INIT(64'b1000010011000001011001001001010101100100110001110100100100111011)  
) LUT6_1492 (
   .O(gates_396),
   .I0(gates_300),
   .I1(gates_5),
   .I2(gates_398),
   .I3(gates_176),
   .I4(gates_367),
   .I5(gates_627)
);
LUT6 #(
   .INIT(64'b1010001010001101001011110111111110100111001111111011001010010111)  
) LUT6_1493 (
   .O(gates_1193),
   .I0(gates_1024),
   .I1(gates_1314),
   .I2(gates_101),
   .I3(gates_902),
   .I4(gates_1109),
   .I5(gates_224)
);
LUT6 #(
   .INIT(64'b0001100100001111011011000110101000111101100010011100111000001001)  
) LUT6_1494 (
   .O(gates_559),
   .I0(gates_1291),
   .I1(gates_1216),
   .I2(gates_212),
   .I3(gates_364),
   .I4(gates_1072),
   .I5(gates_532)
);
LUT6 #(
   .INIT(64'b1000100101010000110011110001000000010010111010010011001101001011)  
) LUT6_1495 (
   .O(gates_303),
   .I0(gates_1237),
   .I1(gates_100),
   .I2(gates_861),
   .I3(gates_122),
   .I4(gates_586),
   .I5(gates_843)
);
LUT6 #(
   .INIT(64'b1100010010111111011110110111001010111010111000110100101001110001)  
) LUT6_1496 (
   .O(gates_1107),
   .I0(gates_373),
   .I1(gates_766),
   .I2(gates_856),
   .I3(gates_149),
   .I4(gates_956),
   .I5(gates_596)
);
LUT6 #(
   .INIT(64'b1100110110111000000111000000000000000011101010001010110111010111)  
) LUT6_1497 (
   .O(gates_299),
   .I0(gates_914),
   .I1(gates_1321),
   .I2(gates_943),
   .I3(gates_1156),
   .I4(gates_73),
   .I5(gates_1421)
);
LUT6 #(
   .INIT(64'b0010110100001100001011011010011011011000110000111011011101110110)  
) LUT6_1498 (
   .O(gates_933),
   .I0(gates_132),
   .I1(gates_1132),
   .I2(gates_835),
   .I3(gates_156),
   .I4(gates_491),
   .I5(gates_921)
);
LUT6 #(
   .INIT(64'b0101101111111010011011010000001010010001110110111000000111111011)  
) LUT6_1499 (
   .O(gates_1361),
   .I0(gates_828),
   .I1(gates_96),
   .I2(gates_129),
   .I3(gates_946),
   .I4(gates_1468),
   .I5(gates_595)
);
LUT6 #(
   .INIT(64'b1110000001011000101011100111110011001001001111010101101100110111)  
) LUT6_1500 (
   .O(gates_227),
   .I0(gates_225),
   .I1(gates_1426),
   .I2(gates_1429),
   .I3(gates_610),
   .I4(gates_1150),
   .I5(gates_1235)
);
LUT6 #(
   .INIT(64'b1111011000110000101001100001101111011111111101000101110001110110)  
) LUT6_1501 (
   .O(gates_1526),
   .I0(gates_561),
   .I1(gates_1224),
   .I2(gates_1294),
   .I3(gates_277),
   .I4(gates_40),
   .I5(gates_1498)
);
LUT6 #(
   .INIT(64'b0010100100010110000000001111100000101011110100111111001000110110)  
) LUT6_1502 (
   .O(gates_488),
   .I0(gates_1194),
   .I1(gates_552),
   .I2(gates_255),
   .I3(gates_676),
   .I4(gates_1551),
   .I5(gates_443)
);
LUT6 #(
   .INIT(64'b0101111111110011010010010001011000000111111100000111010001111100)  
) LUT6_1503 (
   .O(gates_41),
   .I0(gates_829),
   .I1(gates_620),
   .I2(gates_1544),
   .I3(gates_107),
   .I4(gates_1398),
   .I5(gates_1268)
);
LUT6 #(
   .INIT(64'b0110010101011100011011111101011001001110111100010000110000101000)  
) LUT6_1504 (
   .O(gates_420),
   .I0(gates_151),
   .I1(gates_489),
   .I2(gates_218),
   .I3(gates_939),
   .I4(gates_82),
   .I5(gates_120)
);
LUT6 #(
   .INIT(64'b1011010101100111101111111110111011110100101001110001010000100001)  
) LUT6_1505 (
   .O(gates_1533),
   .I0(gates_58),
   .I1(gates_257),
   .I2(gates_104),
   .I3(gates_214),
   .I4(gates_1042),
   .I5(gates_410)
);
LUT6 #(
   .INIT(64'b1101010000011101010100001111100111101010110111111000101001100110)  
) LUT6_1506 (
   .O(gates_236),
   .I0(gates_542),
   .I1(gates_682),
   .I2(gates_1531),
   .I3(gates_140),
   .I4(gates_903),
   .I5(gates_1320)
);
LUT6 #(
   .INIT(64'b0010101111101010010011100110101001110101000001011011000111101001)  
) LUT6_1507 (
   .O(gates_1103),
   .I0(gates_42),
   .I1(gates_49),
   .I2(gates_361),
   .I3(gates_139),
   .I4(gates_1110),
   .I5(gates_314)
);
LUT6 #(
   .INIT(64'b1011011101001110110011001011101100010111110010100101100000011011)  
) LUT6_1508 (
   .O(gates_791),
   .I0(gates_1242),
   .I1(gates_232),
   .I2(gates_153),
   .I3(gates_194),
   .I4(gates_356),
   .I5(gates_1508)
);
LUT6 #(
   .INIT(64'b1101001111010110110001101100111000101110111111110101010010111011)  
) LUT6_1509 (
   .O(gates_1186),
   .I0(gates_1),
   .I1(gates_1333),
   .I2(gates_733),
   .I3(gates_18),
   .I4(gates_887),
   .I5(gates_950)
);
LUT6 #(
   .INIT(64'b0010011011110000010011110011111010000000100011110011000101101001)  
) LUT6_1510 (
   .O(gates_269),
   .I0(gates_908),
   .I1(gates_708),
   .I2(gates_1066),
   .I3(gates_1500),
   .I4(gates_563),
   .I5(gates_978)
);
LUT6 #(
   .INIT(64'b0000110111000111011110100000000000000010110101110000010100101001)  
) LUT6_1511 (
   .O(gates_495),
   .I0(gates_1210),
   .I1(gates_243),
   .I2(gates_654),
   .I3(gates_380),
   .I4(gates_500),
   .I5(gates_1295)
);
LUT6 #(
   .INIT(64'b0001101010001001110011000001100111000001101101001011101000010010)  
) LUT6_1512 (
   .O(gates_160),
   .I0(gates_1056),
   .I1(gates_1190),
   .I2(gates_362),
   .I3(gates_700),
   .I4(gates_1155),
   .I5(gates_900)
);
LUT6 #(
   .INIT(64'b1100110000000101100011110110110100111110010010100011110011010101)  
) LUT6_1513 (
   .O(gates_807),
   .I0(gates_1201),
   .I1(gates_1296),
   .I2(gates_470),
   .I3(gates_128),
   .I4(gates_570),
   .I5(gates_1211)
);
LUT6 #(
   .INIT(64'b0100111101011100010111100011101111001100101011111101010110011101)  
) LUT6_1514 (
   .O(gates_892),
   .I0(gates_1015),
   .I1(gates_1079),
   .I2(gates_1141),
   .I3(gates_838),
   .I4(gates_820),
   .I5(gates_13)
);
LUT6 #(
   .INIT(64'b0101111010001101001100110001010100101010101110001010000101110011)  
) LUT6_1515 (
   .O(gates_746),
   .I0(gates_899),
   .I1(gates_337),
   .I2(gates_1161),
   .I3(gates_233),
   .I4(gates_753),
   .I5(gates_1433)
);
LUT6 #(
   .INIT(64'b1000100011010010110011011111011010110010100010001110011110000011)  
) LUT6_1516 (
   .O(gates_680),
   .I0(gates_925),
   .I1(gates_1053),
   .I2(gates_1263),
   .I3(gates_1030),
   .I4(gates_754),
   .I5(gates_1441)
);
LUT6 #(
   .INIT(64'b0001100000110011100101000100101111100110111100001001011000111011)  
) LUT6_1517 (
   .O(gates_1089),
   .I0(gates_774),
   .I1(gates_1148),
   .I2(gates_330),
   .I3(gates_1347),
   .I4(gates_732),
   .I5(gates_37)
);
LUT6 #(
   .INIT(64'b0101010111000011110101101101000110100011110010010010110011100100)  
) LUT6_1518 (
   .O(gates_1124),
   .I0(gates_591),
   .I1(gates_1341),
   .I2(gates_993),
   .I3(gates_850),
   .I4(gates_296),
   .I5(gates_143)
);
LUT6 #(
   .INIT(64'b0111111100101000110111011001100100010000111101010001011101000011)  
) LUT6_1519 (
   .O(gates_1317),
   .I0(gates_1133),
   .I1(gates_547),
   .I2(gates_1090),
   .I3(gates_421),
   .I4(gates_217),
   .I5(gates_386)
);
LUT6 #(
   .INIT(64'b1000100101000111011111101011101101110111001010011000010001001111)  
) LUT6_1520 (
   .O(gates_110),
   .I0(gates_727),
   .I1(gates_760),
   .I2(gates_790),
   .I3(gates_1435),
   .I4(gates_694),
   .I5(gates_1223)
);
LUT6 #(
   .INIT(64'b0010000111001000100100101011101010000000001101111110010101100001)  
) LUT6_1521 (
   .O(gates_1332),
   .I0(gates_395),
   .I1(gates_982),
   .I2(gates_1016),
   .I3(gates_229),
   .I4(gates_1051),
   .I5(gates_551)
);
LUT6 #(
   .INIT(64'b1100111100100010100010011000011010110010001001011000111100101010)  
) LUT6_1522 (
   .O(gates_1553),
   .I0(gates_945),
   .I1(gates_1264),
   .I2(gates_795),
   .I3(gates_518),
   .I4(gates_419),
   .I5(gates_487)
);
LUT6 #(
   .INIT(64'b0101100000111110110100010011000100010001111001100011101101101011)  
) LUT6_1523 (
   .O(gates_1516),
   .I0(gates_979),
   .I1(gates_1472),
   .I2(gates_2),
   .I3(gates_851),
   .I4(gates_734),
   .I5(gates_239)
);
LUT6 #(
   .INIT(64'b1111101100001001111010010010010001001111101001001100111010000100)  
) LUT6_1524 (
   .O(gates_451),
   .I0(gates_598),
   .I1(gates_848),
   .I2(gates_385),
   .I3(gates_1092),
   .I4(gates_377),
   .I5(gates_1373)
);
LUT6 #(
   .INIT(64'b1000110011100001011100100111011100011111000110110100000101110011)  
) LUT6_1525 (
   .O(gates_1384),
   .I0(gates_117),
   .I1(gates_941),
   .I2(gates_1348),
   .I3(gates_1039),
   .I4(gates_112),
   .I5(gates_348)
);
LUT6 #(
   .INIT(64'b0000111000001101111011011110000101101110100101111001101000000111)  
) LUT6_1526 (
   .O(gates_1004),
   .I0(gates_1129),
   .I1(gates_1272),
   .I2(gates_437),
   .I3(gates_1512),
   .I4(gates_1108),
   .I5(gates_1309)
);
LUT6 #(
   .INIT(64'b0010000000001101000110000110000100010111111100110110110011010111)  
) LUT6_1527 (
   .O(gates_423),
   .I0(gates_196),
   .I1(gates_1459),
   .I2(gates_213),
   .I3(gates_1400),
   .I4(gates_1416),
   .I5(gates_133)
);
LUT6 #(
   .INIT(64'b0110000000001010101110110110100110110110111001001011000010100101)  
) LUT6_1528 (
   .O(gates_1392),
   .I0(gates_1307),
   .I1(gates_952),
   .I2(gates_1327),
   .I3(gates_525),
   .I4(gates_1168),
   .I5(gates_15)
);
LUT6 #(
   .INIT(64'b0100101000000110011101110011100001110001000111111011001000000000)  
) LUT6_1529 (
   .O(gates_736),
   .I0(gates_270),
   .I1(gates_66),
   .I2(gates_473),
   .I3(gates_172),
   .I4(gates_203),
   .I5(gates_969)
);
LUT6 #(
   .INIT(64'b1100100010010001101000101001001100001010110111101110100001101110)  
) LUT6_1530 (
   .O(gates_522),
   .I0(gates_1233),
   .I1(gates_1093),
   .I2(gates_1534),
   .I3(gates_439),
   .I4(gates_756),
   .I5(gates_720)
);
LUT6 #(
   .INIT(64'b1010010001110010011000010101001010000010110010100001000011000010)  
) LUT6_1531 (
   .O(gates_1283),
   .I0(gates_507),
   .I1(gates_1381),
   .I2(gates_958),
   .I3(gates_1485),
   .I4(gates_1119),
   .I5(gates_371)
);
LUT6 #(
   .INIT(64'b1100000011100111101111010100101101010000000001101110000000001010)  
) LUT6_1532 (
   .O(gates_826),
   .I0(gates_1047),
   .I1(gates_428),
   .I2(gates_288),
   .I3(gates_1411),
   .I4(gates_816),
   .I5(gates_962)
);
LUT6 #(
   .INIT(64'b0100011000110011110110101110101110011011011101010100110101111101)  
) LUT6_1533 (
   .O(gates_1396),
   .I0(gates_983),
   .I1(gates_1222),
   .I2(gates_201),
   .I3(gates_179),
   .I4(gates_513),
   .I5(gates_1243)
);
LUT6 #(
   .INIT(64'b0111100001011001001000000110111001110011111001110011111101011001)  
) LUT6_1534 (
   .O(gates_1252),
   .I0(gates_292),
   .I1(gates_323),
   .I2(gates_624),
   .I3(gates_1038),
   .I4(gates_1354),
   .I5(gates_1060)
);
LUT6 #(
   .INIT(64'b0110100000100000000100011001011011100100000010000110001001000101)  
) LUT6_1535 (
   .O(gates_1409),
   .I0(gates_1154),
   .I1(gates_162),
   .I2(gates_936),
   .I3(gates_247),
   .I4(gates_223),
   .I5(gates_704)
);
LUT6 #(
   .INIT(64'b0100011011010001000101000100001011000100100111010000001100101100)  
) LUT6_1536 (
   .O(gates_215),
   .I0(gates_755),
   .I1(gates_512),
   .I2(gates_1050),
   .I3(gates_68),
   .I4(gates_1018),
   .I5(gates_1289)
);
LUT6 #(
   .INIT(64'b1010110000011010101110000010111101101101101010100101111110011011)  
) LUT6_1537 (
   .O(gates_926),
   .I0(gates_1540),
   .I1(gates_1437),
   .I2(gates_450),
   .I3(gates_1206),
   .I4(gates_651),
   .I5(gates_973)
);
LUT6 #(
   .INIT(64'b1111010010110101001010000110100010011000011000111011111000010100)  
) LUT6_1538 (
   .O(gates_374),
   .I0(gates_932),
   .I1(gates_1417),
   .I2(gates_62),
   .I3(gates_1115),
   .I4(gates_1214),
   .I5(gates_847)
);
LUT6 #(
   .INIT(64'b0010110010111111110101110111000110011110001000100000011110000111)  
) LUT6_1539 (
   .O(gates_1412),
   .I0(gates_392),
   .I1(gates_271),
   .I2(gates_1160),
   .I3(gates_713),
   .I4(gates_1353),
   .I5(gates_772)
);
LUT6 #(
   .INIT(64'b1111001010101001000001100101010101100001101100000011000010011000)  
) LUT6_1540 (
   .O(gates_808),
   .I0(gates_1286),
   .I1(gates_251),
   .I2(gates_87),
   .I3(gates_729),
   .I4(gates_35),
   .I5(gates_279)
);
LUT6 #(
   .INIT(64'b0100010111001000110000010101010111110010111000100001111111110011)  
) LUT6_1541 (
   .O(gates_121),
   .I0(gates_56),
   .I1(gates_1340),
   .I2(gates_9),
   .I3(gates_1548),
   .I4(gates_99),
   .I5(gates_27)
);
LUT6 #(
   .INIT(64'b1110101010010111011110100010011010010001100100111000001011011001)  
) LUT6_1542 (
   .O(gates_328),
   .I0(gates_968),
   .I1(gates_516),
   .I2(gates_71),
   .I3(gates_427),
   .I4(gates_1503),
   .I5(gates_972)
);
LUT6 #(
   .INIT(64'b0001110001010010010100001110000111010100100110000101100011001001)  
) LUT6_1543 (
   .O(gates_841),
   .I0(gates_1311),
   .I1(gates_1130),
   .I2(gates_388),
   .I3(gates_1037),
   .I4(gates_33),
   .I5(gates_476)
);
LUT6 #(
   .INIT(64'b0010011000001001011111011000001100011010001010101000000010111000)  
) LUT6_1544 (
   .O(gates_1077),
   .I0(gates_674),
   .I1(gates_701),
   .I2(gates_352),
   .I3(gates_1326),
   .I4(gates_1552),
   .I5(gates_996)
);
LUT6 #(
   .INIT(64'b0111100111001000101001011000100001010100111000010011100011100001)  
) LUT6_1545 (
   .O(gates_1171),
   .I0(gates_559),
   .I1(gates_1193),
   .I2(gates_396),
   .I3(gates_1020),
   .I4(gates_987),
   .I5(gates_240)
);
LUT6 #(
   .INIT(64'b0000100101001111100000101010011110011000001010111010000101101010)  
) LUT6_1546 (
   .O(gates_765),
   .I0(gates_227),
   .I1(gates_1361),
   .I2(gates_933),
   .I3(gates_299),
   .I4(gates_1107),
   .I5(gates_303)
);
LUT6 #(
   .INIT(64'b0001110100100000111010010101011111011001000000010001100000110110)  
) LUT6_1547 (
   .O(gates_1196),
   .I0(gates_236),
   .I1(gates_1533),
   .I2(gates_420),
   .I3(gates_41),
   .I4(gates_488),
   .I5(gates_1526)
);
LUT6 #(
   .INIT(64'b1101111110101010110001000010001000001001100110110000000000111111)  
) LUT6_1548 (
   .O(gates_493),
   .I0(gates_160),
   .I1(gates_495),
   .I2(gates_269),
   .I3(gates_1186),
   .I4(gates_791),
   .I5(gates_1103)
);
LUT6 #(
   .INIT(64'b1001010110010100100000101000100101100101110010011010101101011000)  
) LUT6_1549 (
   .O(gates_961),
   .I0(gates_1124),
   .I1(gates_1089),
   .I2(gates_680),
   .I3(gates_746),
   .I4(gates_892),
   .I5(gates_807)
);
LUT6 #(
   .INIT(64'b0100100000110111111100000101001101110111110001010101011001100100)  
) LUT6_1550 (
   .O(gates_1445),
   .I0(gates_451),
   .I1(gates_1516),
   .I2(gates_1553),
   .I3(gates_1332),
   .I4(gates_110),
   .I5(gates_1317)
);
LUT6 #(
   .INIT(64'b0101110100101110111110000100111001110101110000011000110001011011)  
) LUT6_1551 (
   .O(gates_313),
   .I0(gates_522),
   .I1(gates_736),
   .I2(gates_1392),
   .I3(gates_423),
   .I4(gates_1004),
   .I5(gates_1384)
);
LUT6 #(
   .INIT(64'b0011001001010111110111010010110111111111100100110010000100110011)  
) LUT6_1552 (
   .O(gates_216),
   .I0(gates_215),
   .I1(gates_1409),
   .I2(gates_1252),
   .I3(gates_1396),
   .I4(gates_826),
   .I5(gates_1283)
);
LUT6 #(
   .INIT(64'b0000100000001000001100111101111000000010011011100000100111101110)  
) LUT6_1553 (
   .O(gates_1070),
   .I0(gates_328),
   .I1(gates_121),
   .I2(gates_808),
   .I3(gates_1412),
   .I4(gates_374),
   .I5(gates_926)
);
LUT6 #(
   .INIT(64'b0001010100001010101000010000010000110110101001000110101000101001)  
) LUT6_1554 (
   .O(gates_910),
   .I0(gates_493),
   .I1(gates_1196),
   .I2(gates_765),
   .I3(gates_1171),
   .I4(gates_1077),
   .I5(gates_841)
);
LUT6 #(
   .INIT(64'b0110010010000010000001101010111110110110111110111001011011000011)  
) LUT6_1555 (
   .O(gates_408),
   .I0(gates_910),
   .I1(gates_1070),
   .I2(gates_216),
   .I3(gates_313),
   .I4(gates_1445),
   .I5(gates_961)
);



endmodule