module lut_5level_tree0(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [1728:0] data_in,
                       input       data_valid,
                       output      data_out     
                       );
wire    [1555:0] gates;
reg     [1555:0] gatesReg;
wire    [1728:0] InputBits;


assign gates[0] = 1'b0;

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    gatesReg <= 1556'b0;   
  else
    gatesReg <= gates;
end


assign  InputBits = data_in;
assign  data_out = data_valid & gates[807];

LUT6 #(
   .INIT(64'b0101100011011001101111111000110001011001000001001101100110000000)  
) LUT6_1 (
   .O(gates[127]),
   .I0(InputBits[1077]),
   .I1(InputBits[1123]),
   .I2(InputBits[246]),
   .I3(InputBits[93]),
   .I4(InputBits[1343]),
   .I5(InputBits[1519])
);
LUT6 #(
   .INIT(64'b0010101101010000010111111011011110101110001011101000001000100100)  
) LUT6_2 (
   .O(gates[1049]),
   .I0(InputBits[1372]),
   .I1(InputBits[1257]),
   .I2(InputBits[711]),
   .I3(InputBits[1608]),
   .I4(InputBits[1275]),
   .I5(InputBits[1360])
);
LUT6 #(
   .INIT(64'b0101011110010100110011000000010111001101111101001110100110010000)  
) LUT6_3 (
   .O(gates[71]),
   .I0(InputBits[1170]),
   .I1(InputBits[377]),
   .I2(InputBits[1387]),
   .I3(InputBits[961]),
   .I4(InputBits[1061]),
   .I5(InputBits[1079])
);
LUT6 #(
   .INIT(64'b1001110111110001010100111010000110101101101010011000101000110110)  
) LUT6_4 (
   .O(gates[1481]),
   .I0(InputBits[230]),
   .I1(InputBits[1584]),
   .I2(InputBits[983]),
   .I3(InputBits[893]),
   .I4(InputBits[1414]),
   .I5(InputBits[952])
);
LUT6 #(
   .INIT(64'b1011110111101001100000010111011111110111111111111111001000010010)  
) LUT6_5 (
   .O(gates[882]),
   .I0(InputBits[1166]),
   .I1(InputBits[1496]),
   .I2(InputBits[512]),
   .I3(InputBits[75]),
   .I4(InputBits[996]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0101011111011111010101000010111010101100110010011110100010111000)  
) LUT6_6 (
   .O(gates[1050]),
   .I0(InputBits[1554]),
   .I1(InputBits[1630]),
   .I2(InputBits[599]),
   .I3(InputBits[83]),
   .I4(InputBits[589]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0011011001110111101010011011101100000100001011110101110000010111)  
) LUT6_7 (
   .O(gates[1488]),
   .I0(InputBits[255]),
   .I1(InputBits[648]),
   .I2(InputBits[60]),
   .I3(InputBits[1582]),
   .I4(InputBits[1276]),
   .I5(InputBits[1510])
);
LUT6 #(
   .INIT(64'b0101001000101000001011111001010011101010011111110001000110010000)  
) LUT6_8 (
   .O(gates[560]),
   .I0(InputBits[1377]),
   .I1(InputBits[177]),
   .I2(InputBits[518]),
   .I3(InputBits[832]),
   .I4(InputBits[1199]),
   .I5(InputBits[851])
);
LUT6 #(
   .INIT(64'b1111001000101000100110110110000001001010000111111010001101000011)  
) LUT6_9 (
   .O(gates[1178]),
   .I0(InputBits[1617]),
   .I1(InputBits[1439]),
   .I2(InputBits[369]),
   .I3(InputBits[1701]),
   .I4(InputBits[1163]),
   .I5(InputBits[1487])
);
LUT6 #(
   .INIT(64'b1010101010111110101010110001011000100010100100010010110010100011)  
) LUT6_10 (
   .O(gates[898]),
   .I0(InputBits[1037]),
   .I1(InputBits[105]),
   .I2(InputBits[870]),
   .I3(InputBits[148]),
   .I4(InputBits[1652]),
   .I5(InputBits[735])
);
LUT6 #(
   .INIT(64'b1010101011011010010100100011101111111100100101001111001011010000)  
) LUT6_11 (
   .O(gates[798]),
   .I0(InputBits[759]),
   .I1(InputBits[531]),
   .I2(InputBits[661]),
   .I3(InputBits[261]),
   .I4(InputBits[905]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b0000111110101010011001111011100111111010110010101111110001111001)  
) LUT6_12 (
   .O(gates[1031]),
   .I0(InputBits[1288]),
   .I1(InputBits[955]),
   .I2(InputBits[1144]),
   .I3(InputBits[790]),
   .I4(InputBits[903]),
   .I5(InputBits[1032])
);
LUT6 #(
   .INIT(64'b0110011101000101110110001111000110011011100101010000010111111110)  
) LUT6_13 (
   .O(gates[1387]),
   .I0(InputBits[1569]),
   .I1(InputBits[53]),
   .I2(InputBits[773]),
   .I3(InputBits[1418]),
   .I4(InputBits[1012]),
   .I5(InputBits[1444])
);
LUT6 #(
   .INIT(64'b0000000001111011100000111010000011100111010010000111101101001100)  
) LUT6_14 (
   .O(gates[512]),
   .I0(InputBits[886]),
   .I1(InputBits[1421]),
   .I2(InputBits[919]),
   .I3(InputBits[1677]),
   .I4(InputBits[1334]),
   .I5(InputBits[859])
);
LUT6 #(
   .INIT(64'b1110101001010011000000100001110110011010111011000000010100001011)  
) LUT6_15 (
   .O(gates[463]),
   .I0(InputBits[1369]),
   .I1(InputBits[1683]),
   .I2(InputBits[348]),
   .I3(InputBits[719]),
   .I4(InputBits[639]),
   .I5(InputBits[730])
);
LUT6 #(
   .INIT(64'b1100100111000111001111101011011100010101011101110100101110101011)  
) LUT6_16 (
   .O(gates[1273]),
   .I0(InputBits[1603]),
   .I1(InputBits[1537]),
   .I2(InputBits[447]),
   .I3(InputBits[1309]),
   .I4(InputBits[1212]),
   .I5(InputBits[633])
);
LUT6 #(
   .INIT(64'b0111011010000001001000011100111100110110100000001110010111100111)  
) LUT6_17 (
   .O(gates[517]),
   .I0(InputBits[533]),
   .I1(InputBits[223]),
   .I2(InputBits[112]),
   .I3(InputBits[304]),
   .I4(InputBits[784]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b1011101111001011100111001000010011110101000110000000000101100000)  
) LUT6_18 (
   .O(gates[458]),
   .I0(InputBits[579]),
   .I1(InputBits[1561]),
   .I2(InputBits[1221]),
   .I3(InputBits[804]),
   .I4(InputBits[1684]),
   .I5(InputBits[1346])
);
LUT6 #(
   .INIT(64'b1010010110111011110011010101010100110010100111011011101001101101)  
) LUT6_19 (
   .O(gates[451]),
   .I0(InputBits[1556]),
   .I1(InputBits[879]),
   .I2(InputBits[490]),
   .I3(InputBits[1594]),
   .I4(InputBits[1027]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b1000011011010101110011111101110010011001001101111111110110101010)  
) LUT6_20 (
   .O(gates[454]),
   .I0(InputBits[478]),
   .I1(InputBits[499]),
   .I2(InputBits[173]),
   .I3(InputBits[1230]),
   .I4(InputBits[1669]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b1101110111100001000010101001000010010011101110110001111000111000)  
) LUT6_21 (
   .O(gates[1364]),
   .I0(InputBits[1121]),
   .I1(InputBits[1352]),
   .I2(InputBits[1315]),
   .I3(InputBits[30]),
   .I4(InputBits[322]),
   .I5(InputBits[1384])
);
LUT6 #(
   .INIT(64'b0101100011011011110110101011000110111101000001011100100000000101)  
) LUT6_22 (
   .O(gates[1408]),
   .I0(InputBits[1304]),
   .I1(InputBits[1150]),
   .I2(InputBits[1638]),
   .I3(InputBits[672]),
   .I4(InputBits[1686]),
   .I5(InputBits[1464])
);
LUT6 #(
   .INIT(64'b1110010101100011011010101001011100100111101000111011011010011000)  
) LUT6_23 (
   .O(gates[1250]),
   .I0(InputBits[614]),
   .I1(InputBits[1703]),
   .I2(InputBits[186]),
   .I3(InputBits[212]),
   .I4(InputBits[563]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b1101110001111101011100101010010100010010111001100011101111001110)  
) LUT6_24 (
   .O(gates[1363]),
   .I0(InputBits[682]),
   .I1(InputBits[133]),
   .I2(InputBits[839]),
   .I3(InputBits[1042]),
   .I4(InputBits[775]),
   .I5(InputBits[1294])
);
LUT6 #(
   .INIT(64'b1101110001100011010101000001111000110000100100110011001101100100)  
) LUT6_25 (
   .O(gates[722]),
   .I0(InputBits[316]),
   .I1(InputBits[1099]),
   .I2(InputBits[830]),
   .I3(InputBits[1403]),
   .I4(InputBits[277]),
   .I5(InputBits[1240])
);
LUT6 #(
   .INIT(64'b1010000000101001011111111111000010001110010001000011010011001010)  
) LUT6_26 (
   .O(gates[634]),
   .I0(InputBits[1149]),
   .I1(InputBits[1592]),
   .I2(InputBits[1621]),
   .I3(InputBits[1705]),
   .I4(InputBits[5]),
   .I5(InputBits[1645])
);
LUT6 #(
   .INIT(64'b1101001010011110010011001111101100000011010100000111110100100001)  
) LUT6_27 (
   .O(gates[1109]),
   .I0(InputBits[1481]),
   .I1(InputBits[207]),
   .I2(InputBits[613]),
   .I3(InputBits[1525]),
   .I4(InputBits[506]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0011001100011110001100110011011011101100010000101010001010111100)  
) LUT6_28 (
   .O(gates[578]),
   .I0(InputBits[1155]),
   .I1(InputBits[949]),
   .I2(InputBits[1243]),
   .I3(InputBits[1397]),
   .I4(InputBits[795]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b0010001011111010001110100101011111101110100001101001010111111010)  
) LUT6_29 (
   .O(gates[695]),
   .I0(InputBits[924]),
   .I1(InputBits[1066]),
   .I2(InputBits[1663]),
   .I3(InputBits[492]),
   .I4(InputBits[25]),
   .I5(InputBits[1719])
);
LUT6 #(
   .INIT(64'b1111101100101110010111100100100100011011101100000110100111101101)  
) LUT6_30 (
   .O(gates[978]),
   .I0(InputBits[1382]),
   .I1(InputBits[864]),
   .I2(InputBits[591]),
   .I3(InputBits[1602]),
   .I4(InputBits[1290]),
   .I5(InputBits[969])
);
LUT6 #(
   .INIT(64'b1000111100000101100101111011100101011011010010111110110011011001)  
) LUT6_31 (
   .O(gates[728]),
   .I0(InputBits[927]),
   .I1(InputBits[380]),
   .I2(InputBits[1164]),
   .I3(InputBits[1135]),
   .I4(InputBits[259]),
   .I5(InputBits[1172])
);
LUT6 #(
   .INIT(64'b1000101010111101010110000100100001010011001111111000110110101100)  
) LUT6_32 (
   .O(gates[1244]),
   .I0(InputBits[650]),
   .I1(InputBits[1411]),
   .I2(InputBits[658]),
   .I3(InputBits[1253]),
   .I4(InputBits[523]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b0011010110010100011110100011111100001000110001000111000001111011)  
) LUT6_33 (
   .O(gates[742]),
   .I0(InputBits[1470]),
   .I1(InputBits[1449]),
   .I2(InputBits[1385]),
   .I3(InputBits[1517]),
   .I4(InputBits[418]),
   .I5(InputBits[1355])
);
LUT6 #(
   .INIT(64'b0111000110111000011000010011001010010001111010110000100110101111)  
) LUT6_34 (
   .O(gates[325]),
   .I0(InputBits[436]),
   .I1(InputBits[1472]),
   .I2(InputBits[197]),
   .I3(InputBits[21]),
   .I4(InputBits[1658]),
   .I5(InputBits[1625])
);
LUT6 #(
   .INIT(64'b1010011110111001010001000101111111100110100001100011011001010011)  
) LUT6_35 (
   .O(gates[378]),
   .I0(InputBits[747]),
   .I1(InputBits[1319]),
   .I2(InputBits[1126]),
   .I3(InputBits[203]),
   .I4(InputBits[67]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b1110111001001011110000010001111110101101100100001011111100111011)  
) LUT6_36 (
   .O(gates[29]),
   .I0(InputBits[1190]),
   .I1(InputBits[1508]),
   .I2(InputBits[153]),
   .I3(InputBits[665]),
   .I4(InputBits[356]),
   .I5(InputBits[1301])
);
LUT6 #(
   .INIT(64'b0111100111111010001100010001111011011110001110001010111000011001)  
) LUT6_37 (
   .O(gates[889]),
   .I0(InputBits[973]),
   .I1(InputBits[36]),
   .I2(InputBits[122]),
   .I3(InputBits[1181]),
   .I4(InputBits[479]),
   .I5(InputBits[644])
);
LUT6 #(
   .INIT(64'b1110100100110100010010110000111010000000000101001101011000101001)  
) LUT6_38 (
   .O(gates[350]),
   .I0(InputBits[845]),
   .I1(InputBits[703]),
   .I2(InputBits[619]),
   .I3(InputBits[474]),
   .I4(InputBits[794]),
   .I5(InputBits[1447])
);
LUT6 #(
   .INIT(64'b1010101101111111111110111010100111110010010010110001010100011100)  
) LUT6_39 (
   .O(gates[1233]),
   .I0(InputBits[1197]),
   .I1(InputBits[1168]),
   .I2(InputBits[1558]),
   .I3(InputBits[438]),
   .I4(InputBits[338]),
   .I5(InputBits[91])
);
LUT6 #(
   .INIT(64'b1110100100001010001110100011000001100001011011110110000010010001)  
) LUT6_40 (
   .O(gates[540]),
   .I0(InputBits[788]),
   .I1(InputBits[1455]),
   .I2(InputBits[963]),
   .I3(InputBits[1489]),
   .I4(InputBits[553]),
   .I5(InputBits[821])
);
LUT6 #(
   .INIT(64'b0111100011010111111001001000100010001100111101011011011111011000)  
) LUT6_41 (
   .O(gates[58]),
   .I0(InputBits[428]),
   .I1(InputBits[1545]),
   .I2(InputBits[468]),
   .I3(InputBits[422]),
   .I4(InputBits[199]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b0111011001111110011100100011010100100110100010111111011011000111)  
) LUT6_42 (
   .O(gates[1162]),
   .I0(InputBits[270]),
   .I1(InputBits[114]),
   .I2(InputBits[397]),
   .I3(InputBits[538]),
   .I4(InputBits[1475]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1000100101000000100100011000010010111110000000100110001111111010)  
) LUT6_43 (
   .O(gates[153]),
   .I0(InputBits[1298]),
   .I1(InputBits[1040]),
   .I2(InputBits[59]),
   .I3(InputBits[663]),
   .I4(InputBits[761]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0110010000011011111111100101011011111100011100111001111010110000)  
) LUT6_44 (
   .O(gates[684]),
   .I0(InputBits[404]),
   .I1(InputBits[520]),
   .I2(InputBits[426]),
   .I3(InputBits[1696]),
   .I4(InputBits[990]),
   .I5(InputBits[1206])
);
LUT6 #(
   .INIT(64'b0001110111111100100100010110010110011011011000010011000110111111)  
) LUT6_45 (
   .O(gates[211]),
   .I0(InputBits[1441]),
   .I1(InputBits[319]),
   .I2(InputBits[1650]),
   .I3(InputBits[526]),
   .I4(InputBits[248]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b1110001100011101010010100010011100111100100010000110011111100001)  
) LUT6_46 (
   .O(gates[861]),
   .I0(InputBits[967]),
   .I1(InputBits[753]),
   .I2(InputBits[12]),
   .I3(InputBits[896]),
   .I4(InputBits[221]),
   .I5(InputBits[1010])
);
LUT6 #(
   .INIT(64'b0101100100110011111100000111001010001100101110001100110010010000)  
) LUT6_47 (
   .O(gates[337]),
   .I0(InputBits[603]),
   .I1(InputBits[1492]),
   .I2(InputBits[1021]),
   .I3(InputBits[637]),
   .I4(InputBits[1112]),
   .I5(InputBits[807])
);
LUT6 #(
   .INIT(64'b1010101000111001011010100111111111001111001110000101101101011001)  
) LUT6_48 (
   .O(gates[101]),
   .I0(InputBits[860]),
   .I1(InputBits[1028]),
   .I2(InputBits[1241]),
   .I3(InputBits[1034]),
   .I4(InputBits[440]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b0001011101011010000011101010000110001001110010010101110000101001)  
) LUT6_49 (
   .O(gates[1546]),
   .I0(InputBits[1259]),
   .I1(InputBits[801]),
   .I2(InputBits[101]),
   .I3(InputBits[279]),
   .I4(InputBits[587]),
   .I5(InputBits[655])
);
LUT6 #(
   .INIT(64'b1101111101011111011111011010110111000101110001010101101010011011)  
) LUT6_50 (
   .O(gates[340]),
   .I0(InputBits[109]),
   .I1(InputBits[1656]),
   .I2(InputBits[1103]),
   .I3(InputBits[1178]),
   .I4(InputBits[912]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b1110001111001111100111110001111011011010011110111101011100010111)  
) LUT6_51 (
   .O(gates[76]),
   .I0(InputBits[1225]),
   .I1(InputBits[771]),
   .I2(InputBits[626]),
   .I3(InputBits[389]),
   .I4(InputBits[1534]),
   .I5(InputBits[674])
);
LUT6 #(
   .INIT(64'b1101111000111000110000101001110110011100001111011110000110110110)  
) LUT6_52 (
   .O(gates[311]),
   .I0(InputBits[27]),
   .I1(InputBits[881]),
   .I2(InputBits[1287]),
   .I3(InputBits[44]),
   .I4(InputBits[1458]),
   .I5(InputBits[751])
);
LUT6 #(
   .INIT(64'b0010010101101000011100100110001101111011110011110101010101101111)  
) LUT6_53 (
   .O(gates[982]),
   .I0(InputBits[1345]),
   .I1(InputBits[1035]),
   .I2(InputBits[828]),
   .I3(InputBits[1559]),
   .I4(InputBits[1097]),
   .I5(InputBits[782])
);
LUT6 #(
   .INIT(64'b0000111010100110000111001000010011010000000100101100101010101011)  
) LUT6_54 (
   .O(gates[571]),
   .I0(InputBits[728]),
   .I1(InputBits[1048]),
   .I2(InputBits[688]),
   .I3(InputBits[1131]),
   .I4(InputBits[852]),
   .I5(InputBits[1327])
);
LUT6 #(
   .INIT(64'b1110011010111010101000111011100000001011110101010010011110001010)  
) LUT6_55 (
   .O(gates[1214]),
   .I0(InputBits[1679]),
   .I1(InputBits[107]),
   .I2(InputBits[544]),
   .I3(InputBits[1140]),
   .I4(InputBits[921]),
   .I5(InputBits[1433])
);
LUT6 #(
   .INIT(64'b0000110010000100000011101001000001001101001000100111001010110100)  
) LUT6_56 (
   .O(gates[1190]),
   .I0(InputBits[32]),
   .I1(InputBits[366]),
   .I2(InputBits[4]),
   .I3(InputBits[1311]),
   .I4(InputBits[1662]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1101101011001110111100010101010010100010011110000111000010110111)  
) LUT6_57 (
   .O(gates[825]),
   .I0(InputBits[146]),
   .I1(InputBits[305]),
   .I2(InputBits[561]),
   .I3(InputBits[888]),
   .I4(InputBits[695]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b1100110101010111010001110110101111110111001011101101010011010111)  
) LUT6_58 (
   .O(gates[389]),
   .I0(InputBits[346]),
   .I1(InputBits[382]),
   .I2(InputBits[675]),
   .I3(InputBits[330]),
   .I4(InputBits[1210]),
   .I5(InputBits[1350])
);
LUT6 #(
   .INIT(64'b1011011011010100101011000101010000100010111001001011100001101001)  
) LUT6_59 (
   .O(gates[917]),
   .I0(InputBits[262]),
   .I1(InputBits[744]),
   .I2(InputBits[1265]),
   .I3(InputBits[1053]),
   .I4(InputBits[1059]),
   .I5(InputBits[1152])
);
LUT6 #(
   .INIT(64'b0111001000110010000111110101100110101111110100110000010001001101)  
) LUT6_60 (
   .O(gates[495]),
   .I0(InputBits[1262]),
   .I1(InputBits[1499]),
   .I2(InputBits[1068]),
   .I3(InputBits[694]),
   .I4(InputBits[302]),
   .I5(InputBits[868])
);
LUT6 #(
   .INIT(64'b1111101111011100101111011100100111111111010100101001100001010010)  
) LUT6_61 (
   .O(gates[1345]),
   .I0(InputBits[50]),
   .I1(InputBits[352]),
   .I2(InputBits[876]),
   .I3(InputBits[1615]),
   .I4(InputBits[390]),
   .I5(InputBits[1605])
);
LUT6 #(
   .INIT(64'b0110100010111010110010000101110010000000010110000111100110100010)  
) LUT6_62 (
   .O(gates[1171]),
   .I0(InputBits[1565]),
   .I1(InputBits[1724]),
   .I2(InputBits[766]),
   .I3(InputBits[433]),
   .I4(InputBits[1580]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0000111010011010100001100100000010011111001111111101110110101000)  
) LUT6_63 (
   .O(gates[966]),
   .I0(InputBits[1527]),
   .I1(InputBits[1465]),
   .I2(InputBits[721]),
   .I3(InputBits[1707]),
   .I4(InputBits[19]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0000000110111011010001111101101010011101100100011010001001101010)  
) LUT6_64 (
   .O(gates[1123]),
   .I0(InputBits[1219]),
   .I1(InputBits[1479]),
   .I2(InputBits[1208]),
   .I3(InputBits[216]),
   .I4(InputBits[1416]),
   .I5(InputBits[1434])
);
LUT6 #(
   .INIT(64'b0101110001010000111010101001111110110100101011111101111001000000)  
) LUT6_65 (
   .O(gates[1322]),
   .I0(InputBits[1336]),
   .I1(InputBits[854]),
   .I2(InputBits[1278]),
   .I3(InputBits[169]),
   .I4(InputBits[1089]),
   .I5(InputBits[593])
);
LUT6 #(
   .INIT(64'b1111101101100010111010010000000100110011010011011011110000010001)  
) LUT6_66 (
   .O(gates[992]),
   .I0(InputBits[210]),
   .I1(InputBits[1408]),
   .I2(InputBits[1600]),
   .I3(InputBits[1389]),
   .I4(InputBits[1404]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0100010101100001111111011000010111110110011100100011111100010010)  
) LUT6_67 (
   .O(gates[758]),
   .I0(InputBits[1589]),
   .I1(InputBits[1095]),
   .I2(InputBits[288]),
   .I3(InputBits[1725]),
   .I4(InputBits[1370]),
   .I5(InputBits[1435])
);
LUT6 #(
   .INIT(64'b1011011110111010100100111110010001001100100110111001001111111010)  
) LUT6_68 (
   .O(gates[236]),
   .I0(InputBits[1071]),
   .I1(InputBits[358]),
   .I2(InputBits[684]),
   .I3(InputBits[1474]),
   .I4(InputBits[1157]),
   .I5(InputBits[837])
);
LUT6 #(
   .INIT(64'b1111100000010111111011101110000110101010000011000110100111100111)  
) LUT6_69 (
   .O(gates[706]),
   .I0(InputBits[7]),
   .I1(InputBits[324]),
   .I2(InputBits[269]),
   .I3(InputBits[645]),
   .I4(InputBits[726]),
   .I5(InputBits[1362])
);
LUT6 #(
   .INIT(64'b1010010111110101001111111000111000100100001000111100010111001111)  
) LUT6_70 (
   .O(gates[218]),
   .I0(InputBits[2]),
   .I1(InputBits[314]),
   .I2(InputBits[1635]),
   .I3(InputBits[1502]),
   .I4(InputBits[787]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b0110000011111000000010110100110000011010000111011101000001101101)  
) LUT6_71 (
   .O(gates[1172]),
   .I0(InputBits[749]),
   .I1(InputBits[1321]),
   .I2(InputBits[786]),
   .I3(InputBits[580]),
   .I4(InputBits[1249]),
   .I5(InputBits[1292])
);
LUT6 #(
   .INIT(64'b1111100001101100110010011011010100011100000011000101111110110110)  
) LUT6_72 (
   .O(gates[14]),
   .I0(InputBits[1678]),
   .I1(InputBits[1460]),
   .I2(InputBits[365]),
   .I3(InputBits[276]),
   .I4(InputBits[910]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1001011001100101100011110100001111011010111111111100000011101110)  
) LUT6_73 (
   .O(gates[1259]),
   .I0(InputBits[1310]),
   .I1(InputBits[143]),
   .I2(InputBits[1227]),
   .I3(InputBits[1437]),
   .I4(InputBits[482]),
   .I5(InputBits[1084])
);
LUT6 #(
   .INIT(64'b1111000111111011100011000001110011111000110000110010001010111011)  
) LUT6_74 (
   .O(gates[834]),
   .I0(InputBits[900]),
   .I1(InputBits[843]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[1087]),
   .I5(InputBits[799])
);
LUT6 #(
   .INIT(64'b0000011011110100100010010110110000001000101101111001000011100011)  
) LUT6_75 (
   .O(gates[285]),
   .I0(InputBits[70]),
   .I1(InputBits[281]),
   .I2(InputBits[1431]),
   .I3(InputBits[847]),
   .I4(InputBits[1176]),
   .I5(InputBits[1374])
);
LUT6 #(
   .INIT(64'b1000110011111101011011101000001101011110101001111011000100011011)  
) LUT6_76 (
   .O(gates[234]),
   .I0(InputBits[740]),
   .I1(InputBits[898]),
   .I2(InputBits[286]),
   .I3(InputBits[327]),
   .I4(InputBits[1272]),
   .I5(InputBits[1183])
);
LUT6 #(
   .INIT(64'b0110100000100100101111010110010010110101011101011100100001111111)  
) LUT6_77 (
   .O(gates[594]),
   .I0(InputBits[1466]),
   .I1(InputBits[1031]),
   .I2(InputBits[1203]),
   .I3(InputBits[1610]),
   .I4(InputBits[978]),
   .I5(InputBits[1215])
);
LUT6 #(
   .INIT(64'b0000001011000010001110000000010100011000110010000100001001101100)  
) LUT6_78 (
   .O(gates[1216]),
   .I0(InputBits[1086]),
   .I1(InputBits[1115]),
   .I2(InputBits[1532]),
   .I3(InputBits[1452]),
   .I4(InputBits[29]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b1011011010010011011010010011011011111110101011011110101100011000)  
) LUT6_79 (
   .O(gates[1438]),
   .I0(InputBits[22]),
   .I1(InputBits[601]),
   .I2(InputBits[17]),
   .I3(InputBits[1296]),
   .I4(InputBits[1417]),
   .I5(InputBits[1574])
);
LUT6 #(
   .INIT(64'b0100000100011011111101101101010101100101111001110111000101111100)  
) LUT6_80 (
   .O(gates[1135]),
   .I0(InputBits[595]),
   .I1(InputBits[451]),
   .I2(InputBits[690]),
   .I3(InputBits[1623]),
   .I4(InputBits[1280]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b0101110001001010010110000011001001100001110000101100011100110101)  
) LUT6_81 (
   .O(gates[1203]),
   .I0(InputBits[1314]),
   .I1(InputBits[575]),
   .I2(InputBits[353]),
   .I3(InputBits[170]),
   .I4(InputBits[34]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b1100100100001011010111100000110000110001010000001001001101001001)  
) LUT6_82 (
   .O(gates[96]),
   .I0(InputBits[995]),
   .I1(InputBits[1237]),
   .I2(InputBits[824]),
   .I3(InputBits[1128]),
   .I4(InputBits[1688]),
   .I5(InputBits[1448])
);
LUT6 #(
   .INIT(64'b0110111011000111101011010100000011111010101010101010001000111110)  
) LUT6_83 (
   .O(gates[1068]),
   .I0(InputBits[1064]),
   .I1(InputBits[464]),
   .I2(InputBits[115]),
   .I3(InputBits[455]),
   .I4(InputBits[1110]),
   .I5(InputBits[1279])
);
LUT6 #(
   .INIT(64'b0010111100010111000000111110011001111011000000100111110011111110)  
) LUT6_84 (
   .O(gates[486]),
   .I0(InputBits[57]),
   .I1(InputBits[913]),
   .I2(InputBits[1727]),
   .I3(InputBits[193]),
   .I4(InputBits[572]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0011000000011011111000010001010001101000111111101110010111111110)  
) LUT6_85 (
   .O(gates[1354]),
   .I0(InputBits[628]),
   .I1(InputBits[667]),
   .I2(InputBits[15]),
   .I3(InputBits[1118]),
   .I4(InputBits[345]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b1110011110010001101111111010011110010011101111001111110001110101)  
) LUT6_86 (
   .O(gates[160]),
   .I0(InputBits[1023]),
   .I1(InputBits[116]),
   .I2(InputBits[486]),
   .I3(InputBits[507]),
   .I4(InputBits[1338]),
   .I5(InputBits[1596])
);
LUT6 #(
   .INIT(64'b1000000010101101110101000001110100001001101000000100111011100010)  
) LUT6_87 (
   .O(gates[569]),
   .I0(InputBits[1506]),
   .I1(InputBits[1246]),
   .I2(InputBits[8]),
   .I3(InputBits[1536]),
   .I4(InputBits[611]),
   .I5(InputBits[1331])
);
LUT6 #(
   .INIT(64'b1111110111111100110000100011011001111110001100000011100101110100)  
) LUT6_88 (
   .O(gates[8]),
   .I0(InputBits[988]),
   .I1(InputBits[245]),
   .I2(InputBits[1266]),
   .I3(InputBits[546]),
   .I4(InputBits[162]),
   .I5(InputBits[1507])
);
LUT6 #(
   .INIT(64'b0100111101100110100101000011001101000110010010100000110011010011)  
) LUT6_89 (
   .O(gates[98]),
   .I0(InputBits[1002]),
   .I1(InputBits[1160]),
   .I2(InputBits[550]),
   .I3(InputBits[79]),
   .I4(InputBits[1139]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0000010000100110010100100100010011111110011100100110111001001100)  
) LUT6_90 (
   .O(gates[1278]),
   .I0(InputBits[293]),
   .I1(InputBits[621]),
   .I2(InputBits[1236]),
   .I3(InputBits[1159]),
   .I4(InputBits[1102]),
   .I5(InputBits[755])
);
LUT6 #(
   .INIT(64'b0001000101111010101000100111111010111110000100000010111100011101)  
) LUT6_91 (
   .O(gates[1048]),
   .I0(InputBits[312]),
   .I1(InputBits[940]),
   .I2(InputBits[931]),
   .I3(InputBits[1497]),
   .I4(InputBits[767]),
   .I5(InputBits[883])
);
LUT6 #(
   .INIT(64'b1100000101111010010001001101011011101011001011100101011111101101)  
) LUT6_92 (
   .O(gates[1000]),
   .I0(InputBits[762]),
   .I1(InputBits[1722]),
   .I2(InputBits[68]),
   .I3(InputBits[1691]),
   .I4(InputBits[950]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b1001011001011100001100110111110101000001011001110101011011000101)  
) LUT6_93 (
   .O(gates[1381]),
   .I0(InputBits[1381]),
   .I1(InputBits[654]),
   .I2(InputBits[371]),
   .I3(InputBits[469]),
   .I4(InputBits[819]),
   .I5(InputBits[970])
);
LUT6 #(
   .INIT(64'b0100111011110011101100011111010101101001011111000010110011110000)  
) LUT6_94 (
   .O(gates[1061]),
   .I0(InputBits[495]),
   .I1(InputBits[139]),
   .I2(InputBits[343]),
   .I3(InputBits[764]),
   .I4(InputBits[1186]),
   .I5(InputBits[1073])
);
LUT6 #(
   .INIT(64'b1000110010100001101100100100111000101001000111110100101001110000)  
) LUT6_95 (
   .O(gates[43]),
   .I0(InputBits[915]),
   .I1(InputBits[232]),
   .I2(InputBits[1217]),
   .I3(InputBits[196]),
   .I4(InputBits[696]),
   .I5(InputBits[582])
);
LUT6 #(
   .INIT(64'b0110011101000111000010011110001000000010110110001111101001101011)  
) LUT6_96 (
   .O(gates[686]),
   .I0(InputBits[1628]),
   .I1(InputBits[1260]),
   .I2(InputBits[1524]),
   .I3(InputBits[1239]),
   .I4(InputBits[566]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1011011100011110011101010100110100101000110101000101111110011100)  
) LUT6_97 (
   .O(gates[1396]),
   .I0(InputBits[1515]),
   .I1(InputBits[1153]),
   .I2(InputBits[1007]),
   .I3(InputBits[95]),
   .I4(InputBits[1196]),
   .I5(InputBits[1539])
);
LUT6 #(
   .INIT(64'b1011010101101000100010110010110110010000111111000100001101101000)  
) LUT6_98 (
   .O(gates[391]),
   .I0(InputBits[1234]),
   .I1(InputBits[519]),
   .I2(InputBits[984]),
   .I3(InputBits[1295]),
   .I4(InputBits[992]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0100111000101010000000001101001010010100000001100011111010010010)  
) LUT6_99 (
   .O(gates[193]),
   .I0(InputBits[1224]),
   .I1(InputBits[1693]),
   .I2(InputBits[1364]),
   .I3(InputBits[1398]),
   .I4(InputBits[584]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0001110111010001110111011011000111101110110110010001111101010111)  
) LUT6_100 (
   .O(gates[943]),
   .I0(InputBits[228]),
   .I1(InputBits[373]),
   .I2(InputBits[201]),
   .I3(InputBits[700]),
   .I4(InputBits[81]),
   .I5(InputBits[936])
);
LUT6 #(
   .INIT(64'b0110000111111010100001100001101110111010000100100100110000001100)  
) LUT6_101 (
   .O(gates[288]),
   .I0(InputBits[504]),
   .I1(InputBits[272]),
   .I2(InputBits[959]),
   .I3(InputBits[811]),
   .I4(InputBits[946]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b1011011010010001011001111000110111011101110011001010011101111010)  
) LUT6_102 (
   .O(gates[1555]),
   .I0(InputBits[1550]),
   .I1(InputBits[441]),
   .I2(InputBits[1356]),
   .I3(InputBits[715]),
   .I4(InputBits[220]),
   .I5(InputBits[863])
);
LUT6 #(
   .INIT(64'b0000010011010000011001001110011110101101110011011000001011001000)  
) LUT6_103 (
   .O(gates[119]),
   .I0(InputBits[1577]),
   .I1(InputBits[779]),
   .I2(InputBits[975]),
   .I3(InputBits[510]),
   .I4(InputBits[1401]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b0010101111101000110010100101000011111011101100110001111100000100)  
) LUT6_104 (
   .O(gates[586]),
   .I0(InputBits[1698]),
   .I1(InputBits[834]),
   .I2(InputBits[1009]),
   .I3(InputBits[1690]),
   .I4(InputBits[827]),
   .I5(InputBits[1391])
);
LUT6 #(
   .INIT(64'b1000010000100010101000010110100001101001101001001100100001011111)  
) LUT6_105 (
   .O(gates[180]),
   .I0(InputBits[1093]),
   .I1(InputBits[1080]),
   .I2(InputBits[175]),
   .I3(InputBits[722]),
   .I4(InputBits[798]),
   .I5(InputBits[296])
);
LUT6 #(
   .INIT(64'b0001000000100001010001111011110011110000001111011010110000001101)  
) LUT6_106 (
   .O(gates[1375]),
   .I0(InputBits[1643]),
   .I1(InputBits[1660]),
   .I2(InputBits[1075]),
   .I3(InputBits[604]),
   .I4(InputBits[1504]),
   .I5(InputBits[818])
);
LUT6 #(
   .INIT(64'b0110011111000001110101111101110111010110101101110000110001001010)  
) LUT6_107 (
   .O(gates[410]),
   .I0(InputBits[708]),
   .I1(InputBits[100]),
   .I2(InputBits[388]),
   .I3(InputBits[1708]),
   .I4(InputBits[1318]),
   .I5(InputBits[236])
);
LUT6 #(
   .INIT(64'b1011011100101000001000000101110000000100101000101100111000101111)  
) LUT6_108 (
   .O(gates[246]),
   .I0(InputBits[87]),
   .I1(InputBits[94]),
   .I2(InputBits[671]),
   .I3(InputBits[1323]),
   .I4(InputBits[625]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b1010011000111010111011011111101011001111100010010010001100000110)  
) LUT6_109 (
   .O(gates[690]),
   .I0(InputBits[1214]),
   .I1(InputBits[1193]),
   .I2(InputBits[243]),
   .I3(InputBits[980]),
   .I4(InputBits[77]),
   .I5(InputBits[857])
);
LUT6 #(
   .INIT(64'b1101011111111111001110010010011001110001001100010101001101000010)  
) LUT6_110 (
   .O(gates[999]),
   .I0(InputBits[132]),
   .I1(InputBits[597]),
   .I2(InputBits[724]),
   .I3(InputBits[278]),
   .I4(InputBits[1587]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0110110001110001100011101011101000110000100111010100001110111001)  
) LUT6_111 (
   .O(gates[61]),
   .I0(InputBits[1251]),
   .I1(InputBits[1564]),
   .I2(InputBits[1307]),
   .I3(InputBits[9]),
   .I4(InputBits[234]),
   .I5(InputBits[1477])
);
LUT6 #(
   .INIT(64'b1100011001101001111111111110001111100001101011110001000001101000)  
) LUT6_112 (
   .O(gates[1168]),
   .I0(InputBits[685]),
   .I1(InputBits[462]),
   .I2(InputBits[1108]),
   .I3(InputBits[1637]),
   .I4(InputBits[521]),
   .I5(InputBits[1468])
);
LUT6 #(
   .INIT(64'b1100011101111111110110111010111101110011101100110001011111011000)  
) LUT6_113 (
   .O(gates[1180]),
   .I0(InputBits[1329]),
   .I1(InputBits[1106]),
   .I2(InputBits[283]),
   .I3(InputBits[218]),
   .I4(InputBits[1611]),
   .I5(InputBits[1018])
);
LUT6 #(
   .INIT(64'b0010001111111111110001110011011100000110100000101000110110010110)  
) LUT6_114 (
   .O(gates[1185]),
   .I0(InputBits[1429]),
   .I1(InputBits[1522]),
   .I2(InputBits[1379]),
   .I3(InputBits[1305]),
   .I4(InputBits[102]),
   .I5(InputBits[1586])
);
LUT6 #(
   .INIT(64'b0010010110110000100100111010000001001110101101101001110010000000)  
) LUT6_115 (
   .O(gates[430]),
   .I0(InputBits[835]),
   .I1(InputBits[1454]),
   .I2(InputBits[630]),
   .I3(InputBits[1162]),
   .I4(InputBits[1025]),
   .I5(InputBits[1572])
);
LUT6 #(
   .INIT(64'b1010111111110001100000111110000110110110110000010001000001000100)  
) LUT6_116 (
   .O(gates[447]),
   .I0(InputBits[796]),
   .I1(InputBits[564]),
   .I2(InputBits[198]),
   .I3(InputBits[1632]),
   .I4(InputBits[570]),
   .I5(InputBits[1133])
);
LUT6 #(
   .INIT(64'b1111000011001001010000001101000010111000100000001110001011100001)  
) LUT6_117 (
   .O(gates[1446]),
   .I0(InputBits[292]),
   .I1(InputBits[998]),
   .I2(InputBits[242]),
   .I3(InputBits[1424]),
   .I4(InputBits[359]),
   .I5(InputBits[1715])
);
LUT6 #(
   .INIT(64'b1000100001001010110001000000110110001110000000001010111001100001)  
) LUT6_118 (
   .O(gates[536]),
   .I0(InputBits[891]),
   .I1(InputBits[1484]),
   .I2(InputBits[1014]),
   .I3(InputBits[1406]),
   .I4(InputBits[364]),
   .I5(InputBits[1201])
);
LUT6 #(
   .INIT(64'b1111110101100111010000001111100001110111010000111000100000100001)  
) LUT6_119 (
   .O(gates[1130]),
   .I0(InputBits[150]),
   .I1(InputBits[383]),
   .I2(InputBits[1445]),
   .I3(InputBits[540]),
   .I4(InputBits[1672]),
   .I5(InputBits[1046])
);
LUT6 #(
   .INIT(64'b1110000010001010000000000100101110111100100001111110110100101000)  
) LUT6_120 (
   .O(gates[1315]),
   .I0(InputBits[1044]),
   .I1(InputBits[1405]),
   .I2(InputBits[1552]),
   .I3(InputBits[1423]),
   .I4(InputBits[31]),
   .I5(InputBits[1016])
);
LUT6 #(
   .INIT(64'b0010010101111101011110000000000010101001101000110011001000101111)  
) LUT6_121 (
   .O(gates[415]),
   .I0(InputBits[431]),
   .I1(InputBits[1302]),
   .I2(InputBits[1051]),
   .I3(InputBits[367]),
   .I4(InputBits[1493]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0010110000001110000010110111000011011010011000101111010100010001)  
) LUT6_122 (
   .O(gates[1266]),
   .I0(InputBits[258]),
   .I1(InputBits[1393]),
   .I2(InputBits[842]),
   .I3(InputBits[505]),
   .I4(InputBits[1074]),
   .I5(InputBits[113])
);
LUT6 #(
   .INIT(64'b1101100010110001000101110100001111101010101000001001001111111111)  
) LUT6_123 (
   .O(gates[189]),
   .I0(InputBits[160]),
   .I1(InputBits[742]),
   .I2(InputBits[608]),
   .I3(InputBits[659]),
   .I4(InputBits[58]),
   .I5(InputBits[1349])
);
LUT6 #(
   .INIT(64'b0101111001110001100001111001111011110100010010010001100010101100)  
) LUT6_124 (
   .O(gates[1292]),
   .I0(InputBits[548]),
   .I1(InputBits[1394]),
   .I2(InputBits[791]),
   .I3(InputBits[155]),
   .I4(InputBits[640]),
   .I5(InputBits[669])
);
LUT6 #(
   .INIT(64'b1111001011110001100010010110110000001101111110000010011110000010)  
) LUT6_125 (
   .O(gates[1356]),
   .I0(InputBits[557]),
   .I1(InputBits[866]),
   .I2(InputBits[350]),
   .I3(InputBits[666]),
   .I4(InputBits[1282]),
   .I5(InputBits[1000])
);
LUT6 #(
   .INIT(64'b0011001010110000110100111110001100101101000110110110100100011011)  
) LUT6_126 (
   .O(gates[480]),
   .I0(InputBits[1648]),
   .I1(InputBits[1427]),
   .I2(InputBits[20]),
   .I3(InputBits[257]),
   .I4(InputBits[1681]),
   .I5(InputBits[873])
);
LUT6 #(
   .INIT(64'b0001111111011100110011000001001111110000111010101100101010010110)  
) LUT6_127 (
   .O(gates[438]),
   .I0(InputBits[386]),
   .I1(InputBits[214]),
   .I2(InputBits[1271]),
   .I3(InputBits[652]),
   .I4(InputBits[920]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b1111011001001001001000011101001011000000111111000011110110011100)  
) LUT6_128 (
   .O(gates[1153]),
   .I0(InputBits[917]),
   .I1(InputBits[118]),
   .I2(InputBits[577]),
   .I3(InputBits[977]),
   .I4(InputBits[1626]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0010001100010001001110011100001111101110001110011010110100000111)  
) LUT6_129 (
   .O(gates[107]),
   .I0(InputBits[1057]),
   .I1(InputBits[166]),
   .I2(InputBits[942]),
   .I3(InputBits[624]),
   .I4(InputBits[617]),
   .I5(InputBits[476])
);
LUT6 #(
   .INIT(64'b0010011010000100100111011011010000101000111100111010011111011010)  
) LUT6_130 (
   .O(gates[87]),
   .I0(InputBits[1495]),
   .I1(InputBits[717]),
   .I2(InputBits[334]),
   .I3(InputBits[1137]),
   .I4(InputBits[698]),
   .I5(InputBits[1091])
);
LUT6 #(
   .INIT(64'b1111000011011011101011001010000001110000101011111011100001011000)  
) LUT6_131 (
   .O(gates[1022]),
   .I0(InputBits[878]),
   .I1(InputBits[41]),
   .I2(InputBits[1232]),
   .I3(InputBits[250]),
   .I4(InputBits[1671]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b1011000110100111101100101111011100010100000100000110101110011100)  
) LUT6_132 (
   .O(gates[1458]),
   .I0(InputBits[172]),
   .I1(InputBits[1367]),
   .I2(InputBits[542]),
   .I3(InputBits[1142]),
   .I4(InputBits[1269]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0110001100101101100011010100011000101111101001100001101001010110)  
) LUT6_133 (
   .O(gates[444]),
   .I0(InputBits[1184]),
   .I1(InputBits[181]),
   .I2(InputBits[14]),
   .I3(InputBits[623]),
   .I4(InputBits[460]),
   .I5(InputBits[1354])
);
LUT6 #(
   .INIT(64'b0100001001101100110010011011000101011100010100001110000100001110)  
) LUT6_134 (
   .O(gates[508]),
   .I0(InputBits[1653]),
   .I1(InputBits[987]),
   .I2(InputBits[423]),
   .I3(InputBits[568]),
   .I4(InputBits[809]),
   .I5(InputBits[734])
);
LUT6 #(
   .INIT(64'b1011001101100101101001001000000000001110101110101010101001101010)  
) LUT6_135 (
   .O(gates[953]),
   .I0(InputBits[1005]),
   .I1(InputBits[85]),
   .I2(InputBits[1728]),
   .I3(InputBits[757]),
   .I4(InputBits[1154]),
   .I5(InputBits[1512])
);
LUT6 #(
   .INIT(64'b1010011000100000011010110111111001011110001000011111010000110111)  
) LUT6_136 (
   .O(gates[1336]),
   .I0(InputBits[1541]),
   .I1(InputBits[1120]),
   .I2(InputBits[1147]),
   .I3(InputBits[1175]),
   .I4(InputBits[1700]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0111001010110111110100011011100111010010010001001100011011111001)  
) LUT6_137 (
   .O(gates[221]),
   .I0(InputBits[1038]),
   .I1(InputBits[1641]),
   .I2(InputBits[1575]),
   .I3(InputBits[466]),
   .I4(InputBits[805]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1100101110100111001111011001111110011010011011110001110101110000)  
) LUT6_138 (
   .O(gates[39]),
   .I0(InputBits[1365]),
   .I1(InputBits[141]),
   .I2(InputBits[1613]),
   .I3(InputBits[848]),
   .I4(InputBits[483]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b1001011111010010100001101001001111100110001000101010010011010000)  
) LUT6_139 (
   .O(gates[1424]),
   .I0(InputBits[1568]),
   .I1(InputBits[706]),
   .I2(InputBits[493]),
   .I3(InputBits[1555]),
   .I4(InputBits[536]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b0000000001011001100010001100111111011110010101000111110100100011)  
) LUT6_140 (
   .O(gates[1089]),
   .I0(InputBits[777]),
   .I1(InputBits[416]),
   .I2(InputBits[1375]),
   .I3(InputBits[803]),
   .I4(InputBits[943]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b1000100001010100110010001101101111111101101110100000010000110000)  
) LUT6_141 (
   .O(gates[558]),
   .I0(InputBits[189]),
   .I1(InputBits[692]),
   .I2(InputBits[1619]),
   .I3(InputBits[1562]),
   .I4(InputBits[1312]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0111101110010011110101111010001011111000110100100011010001001000)  
) LUT6_142 (
   .O(gates[417]),
   .I0(InputBits[1316]),
   .I1(InputBits[308]),
   .I2(InputBits[1720]),
   .I3(InputBits[1358]),
   .I4(InputBits[908]),
   .I5(InputBits[745])
);
LUT6 #(
   .INIT(64'b1101110011000111010011011011000001101010000010011011011101111111)  
) LUT6_143 (
   .O(gates[12]),
   .I0(InputBits[925]),
   .I1(InputBits[938]),
   .I2(InputBits[92]),
   .I3(InputBits[341]),
   .I4(InputBits[1340]),
   .I5(InputBits[825])
);
LUT6 #(
   .INIT(64'b1111000110101001000111101000000001000010010010101010010011000010)  
) LUT6_144 (
   .O(gates[1554]),
   .I0(InputBits[813]),
   .I1(InputBits[131]),
   .I2(InputBits[400]),
   .I3(InputBits[1710]),
   .I4(InputBits[1222]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0101000001100110111110100111001110000100001111100110010111101011)  
) LUT6_145 (
   .O(gates[784]),
   .I0(InputBits[1229]),
   .I1(InputBits[119]),
   .I2(InputBits[1639]),
   .I3(InputBits[679]),
   .I4(InputBits[104]),
   .I5(InputBits[1191])
);
LUT6 #(
   .INIT(64'b0110100100001101000111110000010111100101100000110101100001010101)  
) LUT6_146 (
   .O(gates[260]),
   .I0(InputBits[240]),
   .I1(InputBits[1482]),
   .I2(InputBits[673]),
   .I3(InputBits[515]),
   .I4(InputBits[1245]),
   .I5(InputBits[618])
);
LUT6 #(
   .INIT(64'b0111100100010110010100010101101111010110000001000011010011000011)  
) LUT6_147 (
   .O(gates[573]),
   .I0(InputBits[213]),
   .I1(InputBits[1194]),
   .I2(InputBits[968]),
   .I3(InputBits[1718]),
   .I4(InputBits[840]),
   .I5(InputBits[810])
);
LUT6 #(
   .INIT(64'b1001001001100111001001110001010110001100011011001111011100100011)  
) LUT6_148 (
   .O(gates[1084]),
   .I0(InputBits[134]),
   .I1(InputBits[306]),
   .I2(InputBits[752]),
   .I3(InputBits[434]),
   .I4(InputBits[1270]),
   .I5(InputBits[1151])
);
LUT6 #(
   .INIT(64'b0111110010001001100110000010010000100111000101111011101101011001)  
) LUT6_149 (
   .O(gates[1530]),
   .I0(InputBits[606]),
   .I1(InputBits[1342]),
   .I2(InputBits[605]),
   .I3(InputBits[578]),
   .I4(InputBits[99]),
   .I5(InputBits[895])
);
LUT6 #(
   .INIT(64'b1010111001000011100100100000110110110101101111001001010001011111)  
) LUT6_150 (
   .O(gates[762]),
   .I0(InputBits[1713]),
   .I1(InputBits[1461]),
   .I2(InputBits[315]),
   .I3(InputBits[994]),
   .I4(InputBits[681]),
   .I5(InputBits[1674])
);
LUT6 #(
   .INIT(64'b1110000001010110000100111000110110011000111101111011100000000011)  
) LUT6_151 (
   .O(gates[1144]),
   .I0(InputBits[1291]),
   .I1(InputBits[911]),
   .I2(InputBits[1591]),
   .I3(InputBits[1300]),
   .I4(InputBits[1188]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0100011000010010101000000110111101001111001111011000101100001001)  
) LUT6_152 (
   .O(gates[638]),
   .I0(InputBits[1721]),
   .I1(InputBits[1453]),
   .I2(InputBits[465]),
   .I3(InputBits[590]),
   .I4(InputBits[1020]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0010010011010111010001110000010011101101101010101101101001101100)  
) LUT6_153 (
   .O(gates[734]),
   .I0(InputBits[649]),
   .I1(InputBits[1067]),
   .I2(InputBits[1469]),
   .I3(InputBits[1244]),
   .I4(InputBits[237]),
   .I5(InputBits[1335])
);
LUT6 #(
   .INIT(64'b1101110110111101101101001111010111111111100111101001000000111101)  
) LUT6_154 (
   .O(gates[875]),
   .I0(InputBits[217]),
   .I1(InputBits[769]),
   .I2(InputBits[662]),
   .I3(InputBits[778]),
   .I4(InputBits[1119]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1011001101110101100001001101101111011000110101101000101110011100)  
) LUT6_155 (
   .O(gates[1522]),
   .I0(InputBits[1601]),
   .I1(InputBits[1173]),
   .I2(InputBits[497]),
   .I3(InputBits[321]),
   .I4(InputBits[1313]),
   .I5(InputBits[1412])
);
LUT6 #(
   .INIT(64'b1101000110001011011101001100110101010000001110101010111100001001)  
) LUT6_156 (
   .O(gates[1]),
   .I0(InputBits[204]),
   .I1(InputBits[562]),
   .I2(InputBits[419]),
   .I3(InputBits[477]),
   .I4(InputBits[379]),
   .I5(InputBits[981])
);
LUT6 #(
   .INIT(64'b0101000001010001011001001101111111111011110010110110110000010111)  
) LUT6_157 (
   .O(gates[506]),
   .I0(InputBits[948]),
   .I1(InputBits[646]),
   .I2(InputBits[361]),
   .I3(InputBits[928]),
   .I4(InputBits[1471]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1011111001000110011110101110111110001001010010011100000001101000)  
) LUT6_158 (
   .O(gates[136]),
   .I0(InputBits[1252]),
   .I1(InputBits[748]),
   .I2(InputBits[1514]),
   .I3(InputBits[137]),
   .I4(InputBits[1125]),
   .I5(InputBits[704])
);
LUT6 #(
   .INIT(64'b0100010000000001100001011011111110000110010110000010001010001100)  
) LUT6_159 (
   .O(gates[116]),
   .I0(InputBits[1122]),
   .I1(InputBits[1402]),
   .I2(InputBits[290]),
   .I3(InputBits[123]),
   .I4(InputBits[1509]),
   .I5(InputBits[657])
);
LUT6 #(
   .INIT(64'b1110100110010111101101010001110101111000100001000011100101100111)  
) LUT6_160 (
   .O(gates[1197]),
   .I0(InputBits[331]),
   .I1(InputBits[1528]),
   .I2(InputBits[266]),
   .I3(InputBits[417]),
   .I4(InputBits[437]),
   .I5(InputBits[1518])
);
LUT6 #(
   .INIT(64'b0110011011010011101110011011101001100110000110001011110100010001)  
) LUT6_161 (
   .O(gates[144]),
   .I0(InputBits[923]),
   .I1(InputBits[287]),
   .I2(InputBits[785]),
   .I3(InputBits[588]),
   .I4(InputBits[710]),
   .I5(InputBits[822])
);
LUT6 #(
   .INIT(64'b0101101000001101100111101101101011010101110100101101011101111001)  
) LUT6_162 (
   .O(gates[661]),
   .I0(InputBits[894]),
   .I1(InputBits[90]),
   .I2(InputBits[574]),
   .I3(InputBits[945]),
   .I4(InputBits[1607]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b1100110110010001101011010100010111011110110111011100100001111010)  
) LUT6_163 (
   .O(gates[1440]),
   .I0(InputBits[1665]),
   .I1(InputBits[1283]),
   .I2(InputBits[200]),
   .I3(InputBits[1256]),
   .I4(InputBits[299]),
   .I5(InputBits[1371])
);
LUT6 #(
   .INIT(64'b0010011011011100111001010101000110110011100010001110111110010100)  
) LUT6_164 (
   .O(gates[381]),
   .I0(InputBits[1124]),
   .I1(InputBits[1344]),
   .I2(InputBits[1386]),
   .I3(InputBits[1490]),
   .I4(InputBits[627]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b1001011000000111100110110000100001110101100101000110010010011011)  
) LUT6_165 (
   .O(gates[1471]),
   .I0(InputBits[84]),
   .I1(InputBits[636]),
   .I2(InputBits[1062]),
   .I3(InputBits[1376]),
   .I4(InputBits[339]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b0100100000101111011101000011000111101011000011000111101001010001)  
) LUT6_166 (
   .O(gates[581]),
   .I0(InputBits[1583]),
   .I1(InputBits[1581]),
   .I2(InputBits[1328]),
   .I3(InputBits[634]),
   .I4(InputBits[732]),
   .I5(InputBits[985])
);
LUT6 #(
   .INIT(64'b1001101110000010001001010011110010000001001110011001111001000000)  
) LUT6_167 (
   .O(gates[308]),
   .I0(InputBits[705]),
   .I1(InputBits[1553]),
   .I2(InputBits[729]),
   .I3(InputBits[1440]),
   .I4(InputBits[157]),
   .I5(InputBits[789])
);
LUT6 #(
   .INIT(64'b1110100110100110101101010111001111110100010101000111101011100101)  
) LUT6_168 (
   .O(gates[906]),
   .I0(InputBits[1198]),
   .I1(InputBits[997]),
   .I2(InputBits[966]),
   .I3(InputBits[73]),
   .I4(InputBits[906]),
   .I5(InputBits[1631])
);
LUT6 #(
   .INIT(64'b0101110111110011100100100000110101110001100010010011101011111110)  
) LUT6_169 (
   .O(gates[1349]),
   .I0(InputBits[1664]),
   .I1(InputBits[880]),
   .I2(InputBits[1029]),
   .I3(InputBits[408]),
   .I4(InputBits[1167]),
   .I5(InputBits[816])
);
LUT6 #(
   .INIT(64'b0010001010111010111100000001101100011010111100100010111011100101)  
) LUT6_170 (
   .O(gates[177]),
   .I0(InputBits[179]),
   .I1(InputBits[964]),
   .I2(InputBits[530]),
   .I3(InputBits[1368]),
   .I4(InputBits[1055]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0010011000100101101101011000011100100010010100011101010001101000)  
) LUT6_171 (
   .O(gates[678]),
   .I0(InputBits[1675]),
   .I1(InputBits[1395]),
   .I2(InputBits[558]),
   .I3(InputBits[1560]),
   .I4(InputBits[1657]),
   .I5(InputBits[598])
);
LUT6 #(
   .INIT(64'b0000111001111101100101001010011100111101001011101101000110001101)  
) LUT6_172 (
   .O(gates[1517]),
   .I0(InputBits[1651]),
   .I1(InputBits[1419]),
   .I2(InputBits[524]),
   .I3(InputBits[850]),
   .I4(InputBits[1013]),
   .I5(InputBits[871])
);
LUT6 #(
   .INIT(64'b1000101101000110011001011110011001011011001011010001010101100011)  
) LUT6_173 (
   .O(gates[373]),
   .I0(InputBits[677]),
   .I1(InputBits[831]),
   .I2(InputBits[758]),
   .I3(InputBits[1286]),
   .I4(InputBits[1570]),
   .I5(InputBits[877])
);
LUT6 #(
   .INIT(64'b1101100100001011101010011000000000111000110100011101000001000100)  
) LUT6_174 (
   .O(gates[773]),
   .I0(InputBits[687]),
   .I1(InputBits[1274]),
   .I2(InputBits[887]),
   .I3(InputBits[699]),
   .I4(InputBits[432]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0010101010100101111101111101110101011100100010110011111111001010)  
) LUT6_175 (
   .O(gates[1247]),
   .I0(InputBits[1432]),
   .I1(InputBits[13]),
   .I2(InputBits[1026]),
   .I3(InputBits[252]),
   .I4(InputBits[144]),
   .I5(InputBits[1347])
);
LUT6 #(
   .INIT(64'b0010011011110001101000111001011110111010001000000001001111001001)  
) LUT6_176 (
   .O(gates[205]),
   .I0(InputBits[459]),
   .I1(InputBits[1047]),
   .I2(InputBits[922]),
   .I3(InputBits[265]),
   .I4(InputBits[1538]),
   .I5(InputBits[953])
);
LUT6 #(
   .INIT(64'b0001110100110000001100011000111100001011111111111110110010000000)  
) LUT6_177 (
   .O(gates[22]),
   .I0(InputBits[741]),
   .I1(InputBits[736]),
   .I2(InputBits[632]),
   .I3(InputBits[376]),
   .I4(InputBits[1036]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1010110111011011100111110101111101001111110111010101100000110011)  
) LUT6_178 (
   .O(gates[927]),
   .I0(InputBits[555]),
   .I1(InputBits[1289]),
   .I2(InputBits[902]),
   .I3(InputBits[247]),
   .I4(InputBits[413]),
   .I5(InputBits[1220])
);
LUT6 #(
   .INIT(64'b1101011011001111111011101011000010110010000000110011000000000101)  
) LUT6_179 (
   .O(gates[1309]),
   .I0(InputBits[1476]),
   .I1(InputBits[1456]),
   .I2(InputBits[689]),
   .I3(InputBits[1308]),
   .I4(InputBits[1593]),
   .I5(InputBits[1113])
);
LUT6 #(
   .INIT(64'b1100101100101110010111011001001110011110110001110111101100011011)  
) LUT6_180 (
   .O(gates[301]),
   .I0(InputBits[1543]),
   .I1(InputBits[1604]),
   .I2(InputBits[1695]),
   .I3(InputBits[718]),
   .I4(InputBits[856]),
   .I5(InputBits[1557])
);
LUT6 #(
   .INIT(64'b0000110001110101000001110100110000110000111001001010100011100111)  
) LUT6_181 (
   .O(gates[51]),
   .I0(InputBits[1614]),
   .I1(InputBits[145]),
   .I2(InputBits[1293]),
   .I3(InputBits[676]),
   .I4(InputBits[1054]),
   .I5(InputBits[406])
);
LUT6 #(
   .INIT(64'b1101110100010111101110111001110110010000101010000111100001011000)  
) LUT6_182 (
   .O(gates[1260]),
   .I0(InputBits[1540]),
   .I1(InputBits[1676]),
   .I2(InputBits[488]),
   .I3(InputBits[1706]),
   .I4(InputBits[576]),
   .I5(InputBits[1132])
);
LUT6 #(
   .INIT(64'b0111001001101110001100011001111110100000010001100110100011110000)  
) LUT6_183 (
   .O(gates[456]),
   .I0(InputBits[783]),
   .I1(InputBits[457]),
   .I2(InputBits[66]),
   .I3(InputBits[1415]),
   .I4(InputBits[347]),
   .I5(InputBits[776])
);
LUT6 #(
   .INIT(64'b0011101111101101000110111011000000000000001010010110110111000100)  
) LUT6_184 (
   .O(gates[652]),
   .I0(InputBits[6]),
   .I1(InputBits[1646]),
   .I2(InputBits[1702]),
   .I3(InputBits[311]),
   .I4(InputBits[329]),
   .I5(InputBits[565])
);
LUT6 #(
   .INIT(64'b1100011101001101100010110101101101001010010011100011111000000000)  
) LUT6_185 (
   .O(gates[874]),
   .I0(InputBits[446]),
   .I1(InputBits[1661]),
   .I2(InputBits[560]),
   .I3(InputBits[303]),
   .I4(InputBits[763]),
   .I5(InputBits[592])
);
LUT6 #(
   .INIT(64'b1001001010010100101110011011001010001111000000001001001111001001)  
) LUT6_186 (
   .O(gates[975]),
   .I0(InputBits[26]),
   .I1(InputBits[1096]),
   .I2(InputBits[49]),
   .I3(InputBits[1171]),
   .I4(InputBits[1480]),
   .I5(InputBits[1209])
);
LUT6 #(
   .INIT(64'b0010000000011010110100001110010001001100001101010010101101110111)  
) LUT6_187 (
   .O(gates[493]),
   .I0(InputBits[1242]),
   .I1(InputBits[1]),
   .I2(InputBits[254]),
   .I3(InputBits[480]),
   .I4(InputBits[1189]),
   .I5(InputBits[653])
);
LUT6 #(
   .INIT(64'b0111010001001011000001001110101100110010000011010011011101011110)  
) LUT6_188 (
   .O(gates[1033]),
   .I0(InputBits[176]),
   .I1(InputBits[1004]),
   .I2(InputBits[1644]),
   .I3(InputBits[211]),
   .I4(InputBits[191]),
   .I5(InputBits[1060])
);
LUT6 #(
   .INIT(64'b0110111010000011000000111010001001000011001101001110001011111000)  
) LUT6_189 (
   .O(gates[1436]),
   .I0(InputBits[612]),
   .I1(InputBits[425]),
   .I2(InputBits[581]),
   .I3(InputBits[720]),
   .I4(InputBits[1130]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1111011000100111010011100011101111101101100010101000101011000011)  
) LUT6_190 (
   .O(gates[1539]),
   .I0(InputBits[1598]),
   .I1(InputBits[1579]),
   .I2(InputBits[1530]),
   .I3(InputBits[1473]),
   .I4(InputBits[1616]),
   .I5(InputBits[1277])
);
LUT6 #(
   .INIT(64'b0110000110001011011100011000100001010010101010111011011001001001)  
) LUT6_191 (
   .O(gates[1320]),
   .I0(InputBits[517]),
   .I1(InputBits[1726]),
   .I2(InputBits[1694]),
   .I3(InputBits[1566]),
   .I4(InputBits[647]),
   .I5(InputBits[1716])
);
LUT6 #(
   .INIT(64'b1000000110011000010000111001100011100101011011111011100000010001)  
) LUT6_192 (
   .O(gates[796]),
   .I0(InputBits[683]),
   .I1(InputBits[313]),
   .I2(InputBits[1599]),
   .I3(InputBits[1069]),
   .I4(InputBits[208]),
   .I5(InputBits[1410])
);
LUT6 #(
   .INIT(64'b1010101011011100100010001101010001111110111101011011010001000010)  
) LUT6_193 (
   .O(gates[1026]),
   .I0(InputBits[355]),
   .I1(InputBits[235]),
   .I2(InputBits[323]),
   .I3(InputBits[1207]),
   .I4(InputBits[1521]),
   .I5(InputBits[833])
);
LUT6 #(
   .INIT(64'b0101000101100000110101011101111000110000101100111111010100101011)  
) LUT6_194 (
   .O(gates[366]),
   .I0(InputBits[1383]),
   .I1(InputBits[709]),
   .I2(InputBits[135]),
   .I3(InputBits[1409]),
   .I4(InputBits[1709]),
   .I5(InputBits[1156])
);
LUT6 #(
   .INIT(64'b0010000010000010110100011010110101101110011010010010000011010011)  
) LUT6_195 (
   .O(gates[844]),
   .I0(InputBits[545]),
   .I1(InputBits[427]),
   .I2(InputBits[947]),
   .I3(InputBits[1363]),
   .I4(InputBits[838]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1101101101001110000101000011110110100011000001000011001001110100)  
) LUT6_196 (
   .O(gates[1541]),
   .I0(InputBits[1248]),
   .I1(InputBits[1320]),
   .I2(InputBits[1667]),
   .I3(InputBits[1450]),
   .I4(InputBits[285]),
   .I5(InputBits[853])
);
LUT6 #(
   .INIT(64'b1000110001101000110001101100111100110000010010000100000111000000)  
) LUT6_197 (
   .O(gates[1390]),
   .I0(InputBits[514]),
   .I1(InputBits[1590]),
   .I2(InputBits[268]),
   .I3(InputBits[500]),
   .I4(InputBits[712]),
   .I5(InputBits[982])
);
LUT6 #(
   .INIT(64'b0010100110001011110001000011001110111110101010101010101010010011)  
) LUT6_198 (
   .O(gates[272]),
   .I0(InputBits[1396]),
   .I1(InputBits[1255]),
   .I2(InputBits[1649]),
   .I3(InputBits[473]),
   .I4(InputBits[106]),
   .I5(InputBits[1520])
);
LUT6 #(
   .INIT(64'b1010000100001100111000001111100111111100011010111110001011010000)  
) LUT6_199 (
   .O(gates[775]),
   .I0(InputBits[750]),
   .I1(InputBits[1486]),
   .I2(InputBits[51]),
   .I3(InputBits[509]),
   .I4(InputBits[37]),
   .I5(InputBits[378])
);
LUT6 #(
   .INIT(64'b0101101000010100100000010011101000101111100110001000110001111100)  
) LUT6_200 (
   .O(gates[1469]),
   .I0(InputBits[202]),
   .I1(InputBits[467]),
   .I2(InputBits[127]),
   .I3(InputBits[525]),
   .I4(InputBits[1226]),
   .I5(InputBits[1442])
);
LUT6 #(
   .INIT(64'b1101110101000100101110110001110110000111010010111111101000111010)  
) LUT6_201 (
   .O(gates[1499]),
   .I0(InputBits[861]),
   .I1(InputBits[552]),
   .I2(InputBits[142]),
   .I3(InputBits[43]),
   .I4(InputBits[656]),
   .I5(InputBits[727])
);
LUT6 #(
   .INIT(64'b1111010010111010100101101100011000111101010111011011010100010110)  
) LUT6_202 (
   .O(gates[746]),
   .I0(InputBits[215]),
   .I1(InputBits[1205]),
   .I2(InputBits[301]),
   .I3(InputBits[974]),
   .I4(InputBits[1180]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b1100110000110100101110011000101100111010110000001110000011110100)  
) LUT6_203 (
   .O(gates[400]),
   .I0(InputBits[760]),
   .I1(InputBits[802]),
   .I2(InputBits[929]),
   .I3(InputBits[702]),
   .I4(InputBits[889]),
   .I5(InputBits[1104])
);
LUT6 #(
   .INIT(64'b0110010100101010111100011011010110011011110010110100011011100000)  
) LUT6_204 (
   .O(gates[534]),
   .I0(InputBits[1430]),
   .I1(InputBits[793]),
   .I2(InputBits[691]),
   .I3(InputBits[1090]),
   .I4(InputBits[439]),
   .I5(InputBits[1697])
);
LUT6 #(
   .INIT(64'b1000101111011011110010110111100000010101110101001101111011100111)  
) LUT6_205 (
   .O(gates[919]),
   .I0(InputBits[1078]),
   .I1(InputBits[1655]),
   .I2(InputBits[71]),
   .I3(InputBits[1618]),
   .I4(InputBits[664]),
   .I5(InputBits[586])
);
LUT6 #(
   .INIT(64'b0011100001111101000101010110010001101001001001010101100110111100)  
) LUT6_206 (
   .O(gates[744]),
   .I0(InputBits[904]),
   .I1(InputBits[909]),
   .I2(InputBits[642]),
   .I3(InputBits[161]),
   .I4(InputBits[1299]),
   .I5(InputBits[226])
);
LUT6 #(
   .INIT(64'b0000010010000001110100100110100000000101111110111001111100011010)  
) LUT6_207 (
   .O(gates[1268]),
   .I0(InputBits[108]),
   .I1(InputBits[1333]),
   .I2(InputBits[128]),
   .I3(InputBits[602]),
   .I4(InputBits[56]),
   .I5(InputBits[858])
);
LUT6 #(
   .INIT(64'b0000010100010001100001110101011001111100100010101011111111100000)  
) LUT6_208 (
   .O(gates[20]),
   .I0(InputBits[1011]),
   .I1(InputBits[1491]),
   .I2(InputBits[280]),
   .I3(InputBits[11]),
   .I4(InputBits[829]),
   .I5(InputBits[1326])
);
LUT6 #(
   .INIT(64'b0111011111001011110001111111100011100101000100001001010001010101)  
) LUT6_209 (
   .O(gates[888]),
   .I0(InputBits[260]),
   .I1(InputBits[1082]),
   .I2(InputBits[534]),
   .I3(InputBits[532]),
   .I4(InputBits[1546]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1001000011101010100111111101111010111111111111111101110101110010)  
) LUT6_210 (
   .O(gates[633]),
   .I0(InputBits[629]),
   .I1(InputBits[743]),
   .I2(InputBits[1606]),
   .I3(InputBits[1463]),
   .I4(InputBits[808]),
   .I5(InputBits[781])
);
LUT6 #(
   .INIT(64'b1001011001101010011100010110100001010010100100011110000011000000)  
) LUT6_211 (
   .O(gates[1372]),
   .I0(InputBits[1353]),
   .I1(InputBits[738]),
   .I2(InputBits[152]),
   .I3(InputBits[956]),
   .I4(InputBits[1548]),
   .I5(InputBits[1049])
);
LUT6 #(
   .INIT(64'b0101110101101100111111010110110100010000010111101000111010011101)  
) LUT6_212 (
   .O(gates[1011]),
   .I0(InputBits[1533]),
   .I1(InputBits[337]),
   .I2(InputBits[635]),
   .I3(InputBits[222]),
   .I4(InputBits[489]),
   .I5(InputBits[991])
);
LUT6 #(
   .INIT(64'b0011010010000100100001111001100110110011000110000011011011010101)  
) LUT6_213 (
   .O(gates[151]),
   .I0(InputBits[1258]),
   .I1(InputBits[939]),
   .I2(InputBits[1169]),
   .I3(InputBits[962]),
   .I4(InputBits[1022]),
   .I5(InputBits[1111])
);
LUT6 #(
   .INIT(64'b1111011111101101101100010101100111010101100000101010101101001011)  
) LUT6_214 (
   .O(gates[468]),
   .I0(InputBits[1457]),
   .I1(InputBits[774]),
   .I2(InputBits[1179]),
   .I3(InputBits[410]),
   .I4(InputBits[45]),
   .I5(InputBits[1685])
);
LUT6 #(
   .INIT(64'b0001100111000110000010101100101111011001111101000011010001001110)  
) LUT6_215 (
   .O(gates[1161]),
   .I0(InputBits[185]),
   .I1(InputBits[1425]),
   .I2(InputBits[1098]),
   .I3(InputBits[1195]),
   .I4(InputBits[1101]),
   .I5(InputBits[972])
);
LUT6 #(
   .INIT(64'b0100001111011010111101000011000100000000000011001110011101100110)  
) LUT6_216 (
   .O(gates[1285]),
   .I0(InputBits[993]),
   .I1(InputBits[527]),
   .I2(InputBits[295]),
   .I3(InputBits[1501]),
   .I4(InputBits[1058]),
   .I5(InputBits[1138])
);
LUT6 #(
   .INIT(64'b1100100100000101110011010100110111011011110000011010101110100001)  
) LUT6_217 (
   .O(gates[1019]),
   .I0(InputBits[409]),
   .I1(InputBits[1547]),
   .I2(InputBits[1692]),
   .I3(InputBits[1070]),
   .I4(InputBits[1158]),
   .I5(InputBits[1263])
);
LUT6 #(
   .INIT(64'b1011110011100101010110111011010001101101010001010000110001001111)  
) LUT6_218 (
   .O(gates[700]),
   .I0(InputBits[869]),
   .I1(InputBits[916]),
   .I2(InputBits[64]),
   .I3(InputBits[1711]),
   .I4(InputBits[551]),
   .I5(InputBits[1141])
);
LUT6 #(
   .INIT(64'b1010011001010010011011110010100010100001010001000110001110100100)  
) LUT6_219 (
   .O(gates[287]),
   .I0(InputBits[1325]),
   .I1(InputBits[756]),
   .I2(InputBits[1523]),
   .I3(InputBits[643]),
   .I4(InputBits[138]),
   .I5(InputBits[1001])
);
LUT6 #(
   .INIT(64'b1001111111000010011011101101001111010011011010001101100100111010)  
) LUT6_220 (
   .O(gates[78]),
   .I0(InputBits[1392]),
   .I1(InputBits[251]),
   .I2(InputBits[733]),
   .I3(InputBits[183]),
   .I4(InputBits[231]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b1011100010100001001100011010101001111001011001010101101100011110)  
) LUT6_221 (
   .O(gates[475]),
   .I0(InputBits[294]),
   .I1(InputBits[1399]),
   .I2(InputBits[765]),
   .I3(InputBits[1094]),
   .I4(InputBits[1185]),
   .I5(InputBits[885])
);
LUT6 #(
   .INIT(64'b0000110111001011101100110011111101011101010001110111101000010010)  
) LUT6_222 (
   .O(gates[1380]),
   .I0(InputBits[585]),
   .I1(InputBits[1233]),
   .I2(InputBits[716]),
   .I3(InputBits[1670]),
   .I4(InputBits[812]),
   .I5(InputBits[1218])
);
LUT6 #(
   .INIT(64'b0010011000010101111101101010101100010011010110101100001001110000)  
) LUT6_223 (
   .O(gates[413]),
   .I0(InputBits[1500]),
   .I1(InputBits[1704]),
   .I2(InputBits[445]),
   .I3(InputBits[882]),
   .I4(InputBits[976]),
   .I5(InputBits[890])
);
LUT6 #(
   .INIT(64'b0100000011000100111010001101100111000011100011110110100011001111)  
) LUT6_224 (
   .O(gates[990]),
   .I0(InputBits[1576]),
   .I1(InputBits[1134]),
   .I2(InputBits[1485]),
   .I3(InputBits[874]),
   .I4(InputBits[1516]),
   .I5(InputBits[1235])
);
LUT6 #(
   .INIT(64'b1110001010011101011110010010101110001000010101101111110011110100)  
) LUT6_225 (
   .O(gates[294]),
   .I0(InputBits[1717]),
   .I1(InputBits[384]),
   .I2(InputBits[855]),
   .I3(InputBits[424]),
   .I4(InputBits[1542]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b1110010110001111000100100111001110111000101110100111110110101100)  
) LUT6_226 (
   .O(gates[349]),
   .I0(InputBits[1511]),
   .I1(InputBits[374]),
   .I2(InputBits[930]),
   .I3(InputBits[182]),
   .I4(InputBits[393]),
   .I5(InputBits[1588])
);
LUT6 #(
   .INIT(64'b1100001011101100110000010010100011111100001110111100010011110101)  
) LUT6_227 (
   .O(gates[932]),
   .I0(InputBits[403]),
   .I1(InputBits[407]),
   .I2(InputBits[1578]),
   .I3(InputBits[1006]),
   .I4(InputBits[54]),
   .I5(InputBits[415])
);
LUT6 #(
   .INIT(64'b0001001010010000001110111001100101011100101011111110110110010110)  
) LUT6_228 (
   .O(gates[1442]),
   .I0(InputBits[836]),
   .I1(InputBits[225]),
   .I2(InputBits[1668]),
   .I3(InputBits[1689]),
   .I4(InputBits[567]),
   .I5(InputBits[1264])
);
LUT6 #(
   .INIT(64'b0111011010110001010000011110101110100100011110000000011110100111)  
) LUT6_229 (
   .O(gates[764]),
   .I0(InputBits[309]),
   .I1(InputBits[725]),
   .I2(InputBits[1659]),
   .I3(InputBits[48]),
   .I4(InputBits[875]),
   .I5(InputBits[678])
);
LUT6 #(
   .INIT(64'b0101101111101100001100010111000100000000111100001110110101011111)  
) LUT6_230 (
   .O(gates[1549]),
   .I0(InputBits[1388]),
   .I1(InputBits[326]),
   .I2(InputBits[1041]),
   .I3(InputBits[826]),
   .I4(InputBits[707]),
   .I5(InputBits[1216])
);
LUT6 #(
   .INIT(64'b0101000101011001001111011000011100001010110100100101111011011011)  
) LUT6_231 (
   .O(gates[1525]),
   .I0(InputBits[820]),
   .I1(InputBits[381]),
   .I2(InputBits[701]),
   .I3(InputBits[1204]),
   .I4(InputBits[494]),
   .I5(InputBits[103])
);
LUT6 #(
   .INIT(64'b0100000000011111101001011110001101011001000011000100111100101000)  
) LUT6_232 (
   .O(gates[515]),
   .I0(InputBits[1357]),
   .I1(InputBits[1642]),
   .I2(InputBits[88]),
   .I3(InputBits[957]),
   .I4(InputBits[10]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0111101001100111001101001001001111101010111001010011011110101110)  
) LUT6_233 (
   .O(gates[1242]),
   .I0(InputBits[502]),
   .I1(InputBits[241]),
   .I2(InputBits[80]),
   .I3(InputBits[806]),
   .I4(InputBits[1443]),
   .I5(InputBits[620])
);
LUT6 #(
   .INIT(64'b0110001000100100100111110111000010101001000010001001101000000011)  
) LUT6_234 (
   .O(gates[1107]),
   .I0(InputBits[1083]),
   .I1(InputBits[317]),
   .I2(InputBits[935]),
   .I3(InputBits[1008]),
   .I4(InputBits[503]),
   .I5(InputBits[1531])
);
LUT6 #(
   .INIT(64'b0001100010101100010110001010000000001100100000001110010000010000)  
) LUT6_235 (
   .O(gates[1208]),
   .I0(InputBits[78]),
   .I1(InputBits[1088]),
   .I2(InputBits[1322]),
   .I3(InputBits[1380]),
   .I4(InputBits[387]),
   .I5(InputBits[958])
);
LUT6 #(
   .INIT(64'b1001011100010000110101000010101100100111100110111011010001110001)  
) LUT6_236 (
   .O(gates[138]),
   .I0(InputBits[487]),
   .I1(InputBits[450]),
   .I2(InputBits[151]),
   .I3(InputBits[284]),
   .I4(InputBits[1273]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1101001001100110011101100000010101101011001001010110000001100110)  
) LUT6_237 (
   .O(gates[606]),
   .I0(InputBits[631]),
   .I1(InputBits[1285]),
   .I2(InputBits[47]),
   .I3(InputBits[452]),
   .I4(InputBits[405]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b0100000101110101100001101110010111100101101001001101111100000011)  
) LUT6_238 (
   .O(gates[1383]),
   .I0(InputBits[800]),
   .I1(InputBits[1228]),
   .I2(InputBits[357]),
   .I3(InputBits[609]),
   .I4(InputBits[737]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b1011011011100000100100000101010100100010001010111101101100000000)  
) LUT6_239 (
   .O(gates[137]),
   .I0(InputBits[1467]),
   .I1(InputBits[125]),
   .I2(InputBits[398]),
   .I3(InputBits[1324]),
   .I4(InputBits[1202]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1011010000000101111000101101011110011100011110100011011001011111)  
) LUT6_240 (
   .O(gates[1414]),
   .I0(InputBits[899]),
   .I1(InputBits[522]),
   .I2(InputBits[481]),
   .I3(InputBits[484]),
   .I4(InputBits[192]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1000111011010111010010111000101100000111110111101111010110010111)  
) LUT6_241 (
   .O(gates[724]),
   .I0(InputBits[1573]),
   .I1(InputBits[1030]),
   .I2(InputBits[69]),
   .I3(InputBits[244]),
   .I4(InputBits[1337]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0011110010111010110001110011111001110011010101101110010110101100)  
) LUT6_242 (
   .O(gates[1201]),
   .I0(InputBits[140]),
   .I1(InputBits[979]),
   .I2(InputBits[823]),
   .I3(InputBits[1428]),
   .I4(InputBits[149]),
   .I5(InputBits[1459])
);
LUT6 #(
   .INIT(64'b0011010101010100100000001100111101100101011000000011100110010110)  
) LUT6_243 (
   .O(gates[432]),
   .I0(InputBits[1529]),
   .I1(InputBits[1332]),
   .I2(InputBits[194]),
   .I3(InputBits[897]),
   .I4(InputBits[573]),
   .I5(InputBits[668])
);
LUT6 #(
   .INIT(64'b0101010000001011110110110110000111111010000100010000100110000110)  
) LUT6_244 (
   .O(gates[666]),
   .I0(InputBits[1146]),
   .I1(InputBits[1129]),
   .I2(InputBits[1597]),
   .I3(InputBits[1015]),
   .I4(InputBits[385]),
   .I5(InputBits[754])
);
LUT6 #(
   .INIT(64'b0011101111110010111000110010011111110001110010010110010000001111)  
) LUT6_245 (
   .O(gates[519]),
   .I0(InputBits[86]),
   .I1(InputBits[360]),
   .I2(InputBits[1407]),
   .I3(InputBits[1109]),
   .I4(InputBits[1182]),
   .I5(InputBits[1629])
);
LUT6 #(
   .INIT(64'b0001111110110010110001110111001000101100111111000101100011101010)  
) LUT6_246 (
   .O(gates[1074]),
   .I0(InputBits[513]),
   .I1(InputBits[171]),
   .I2(InputBits[1003]),
   .I3(InputBits[1348]),
   .I4(InputBits[1117]),
   .I5(InputBits[610])
);
LUT6 #(
   .INIT(64'b0100011101011101100111001000111100001010110111001010110000110101)  
) LUT6_247 (
   .O(gates[860]),
   .I0(InputBits[263]),
   .I1(InputBits[792]),
   .I2(InputBits[539]),
   .I3(InputBits[282]),
   .I4(InputBits[159]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b1011001100000111100100010110100100010111001100101101110110110011)  
) LUT6_248 (
   .O(gates[1195]),
   .I0(InputBits[351]),
   .I1(InputBits[1231]),
   .I2(InputBits[1535]),
   .I3(InputBits[117]),
   .I4(InputBits[1422]),
   .I5(InputBits[1680])
);
LUT6 #(
   .INIT(64'b0001011010111000011100100101100101110000100000110000000111111111)  
) LUT6_249 (
   .O(gates[1063]),
   .I0(InputBits[768]),
   .I1(InputBits[770]),
   .I2(InputBits[130]),
   .I3(InputBits[456]),
   .I4(InputBits[336]),
   .I5(InputBits[1494])
);
LUT6 #(
   .INIT(64'b0011101101101101000010010100000110100100111110110001001110111010)  
) LUT6_250 (
   .O(gates[17]),
   .I0(InputBits[1267]),
   .I1(InputBits[1213]),
   .I2(InputBits[713]),
   .I3(InputBits[1478]),
   .I4(InputBits[772]),
   .I5(InputBits[714])
);
LUT6 #(
   .INIT(64'b0111101001011100000001011000000111100000100111001011011000111011)  
) LUT6_251 (
   .O(gates[1327]),
   .I0(InputBits[1624]),
   .I1(InputBits[1634]),
   .I2(InputBits[1359]),
   .I3(InputBits[989]),
   .I4(InputBits[1351]),
   .I5(InputBits[986])
);
LUT6 #(
   .INIT(64'b0010011111111010110011001111111010100011101110010001010110111010)  
) LUT6_252 (
   .O(gates[1274]),
   .I0(InputBits[1666]),
   .I1(InputBits[1177]),
   .I2(InputBits[1297]),
   .I3(InputBits[600]),
   .I4(InputBits[38]),
   .I5(InputBits[844])
);
LUT6 #(
   .INIT(64'b1101100111101001010011000110010011011101100111000110000100110010)  
) LUT6_253 (
   .O(gates[708]),
   .I0(InputBits[156]),
   .I1(InputBits[1436]),
   .I2(InputBits[1052]),
   .I3(InputBits[1281]),
   .I4(InputBits[547]),
   .I5(InputBits[1024])
);
LUT6 #(
   .INIT(64'b1111110010001001100110010110111010100110101101011101101000011010)  
) LUT6_254 (
   .O(gates[110]),
   .I0(InputBits[1687]),
   .I1(InputBits[461]),
   .I2(InputBits[1627]),
   .I3(InputBits[1513]),
   .I4(InputBits[165]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0001111010001111010101110001111010100111001100100010011101011011)  
) LUT6_255 (
   .O(gates[333]),
   .I0(InputBits[1498]),
   .I1(InputBits[651]),
   .I2(InputBits[622]),
   .I3(InputBits[333]),
   .I4(InputBits[941]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0110000000001101010001100000110110100100011001010100010110011001)  
) LUT6_256 (
   .O(gates[710]),
   .I0(InputBits[1712]),
   .I1(InputBits[731]),
   .I2(InputBits[814]),
   .I3(InputBits[375]),
   .I4(InputBits[1092]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b1001101110011111001101010100110101001111000110111110111110001001)  
) LUT6_257 (
   .O(gates[323]),
   .I0(InputBits[1261]),
   .I1(InputBits[195]),
   .I2(InputBits[253]),
   .I3(InputBits[184]),
   .I4(InputBits[1247]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b1100011101000111101000000010111000110001010110011011000010101111)  
) LUT6_258 (
   .O(gates[856]),
   .I0(InputBits[496]),
   .I1(InputBits[1127]),
   .I2(InputBits[1268]),
   .I3(InputBits[1446]),
   .I4(InputBits[934]),
   .I5(InputBits[849])
);
LUT6 #(
   .INIT(64'b1101100101001100110000111110011010010110111110010010001111111110)  
) LUT6_259 (
   .O(gates[112]),
   .I0(InputBits[1100]),
   .I1(InputBits[1622]),
   .I2(InputBits[954]),
   .I3(InputBits[1148]),
   .I4(InputBits[1400]),
   .I5(InputBits[616])
);
LUT6 #(
   .INIT(64'b1011001100001101100101110011011101101101111100111101100011110000)  
) LUT6_260 (
   .O(gates[545]),
   .I0(InputBits[1056]),
   .I1(InputBits[411]),
   .I2(InputBits[454]),
   .I3(InputBits[110]),
   .I4(InputBits[354]),
   .I5(InputBits[1072])
);
LUT6 #(
   .INIT(64'b1101000111011101010000100000101001101000100000101111000100110111)  
) LUT6_261 (
   .O(gates[191]),
   .I0(InputBits[227]),
   .I1(InputBits[884]),
   .I2(InputBits[1143]),
   .I3(InputBits[697]),
   .I4(InputBits[1187]),
   .I5(InputBits[951])
);
LUT6 #(
   .INIT(64'b0010001001111010011111100100010011101000000010101100110010110111)  
) LUT6_262 (
   .O(gates[187]),
   .I0(InputBits[529]),
   .I1(InputBits[918]),
   .I2(InputBits[1043]),
   .I3(InputBits[1654]),
   .I4(InputBits[1567]),
   .I5(InputBits[615])
);
LUT6 #(
   .INIT(64'b0011011101111000000000010100011001101101100000100110010111101001)  
) LUT6_263 (
   .O(gates[588]),
   .I0(InputBits[1341]),
   .I1(InputBits[780]),
   .I2(InputBits[867]),
   .I3(InputBits[1366]),
   .I4(InputBits[435]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1000101100011111010011011011111110111001010100101100000111100001)  
) LUT6_264 (
   .O(gates[646]),
   .I0(InputBits[1699]),
   .I1(InputBits[97]),
   .I2(InputBits[846]),
   .I3(InputBits[1640]),
   .I4(InputBits[937]),
   .I5(InputBits[907])
);
LUT6 #(
   .INIT(64'b0010110111010000111001001010000101001100100000101000100011001100)  
) LUT6_265 (
   .O(gates[756]),
   .I0(InputBits[498]),
   .I1(InputBits[1378]),
   .I2(InputBits[554]),
   .I3(InputBits[154]),
   .I4(InputBits[746]),
   .I5(InputBits[472])
);
LUT6 #(
   .INIT(64'b1010100000101010010010101010001111010001000101010100010010111111)  
) LUT6_266 (
   .O(gates[446]),
   .I0(InputBits[926]),
   .I1(InputBits[914]),
   .I2(InputBits[1317]),
   .I3(InputBits[190]),
   .I4(InputBits[1039]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b0001111110111100011000001100101100000001001110001000100110001110)  
) LUT6_267 (
   .O(gates[262]),
   .I0(InputBits[535]),
   .I1(InputBits[307]),
   .I2(InputBits[797]),
   .I3(InputBits[569]),
   .I4(InputBits[342]),
   .I5(InputBits[1105])
);
LUT6 #(
   .INIT(64'b1010010111110100010111010101110001001110000011100010110010011100)  
) LUT6_268 (
   .O(gates[1283]),
   .I0(InputBits[297]),
   .I1(InputBits[1136]),
   .I2(InputBits[817]),
   .I3(InputBits[1503]),
   .I4(InputBits[401]),
   .I5(InputBits[1390])
);
LUT6 #(
   .INIT(64'b0001111111100101111100000010000100111010011111100111101011100111)  
) LUT6_269 (
   .O(gates[1220]),
   .I0(InputBits[693]),
   .I1(InputBits[1223]),
   .I2(InputBits[680]),
   .I3(InputBits[1620]),
   .I4(InputBits[1526]),
   .I5(InputBits[1254])
);
LUT6 #(
   .INIT(64'b1001100110101011011101011000100010111011011000010100001111111010)  
) LUT6_270 (
   .O(gates[212]),
   .I0(InputBits[1544]),
   .I1(InputBits[1723]),
   .I2(InputBits[1076]),
   .I3(InputBits[723]),
   .I4(InputBits[872]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b1010000000001111111100000100100011100111011100111000001001011010)  
) LUT6_271 (
   .O(gates[1331]),
   .I0(InputBits[82]),
   .I1(InputBits[1211]),
   .I2(InputBits[1373]),
   .I3(InputBits[239]),
   .I4(InputBits[638]),
   .I5(InputBits[1081])
);
LUT6 #(
   .INIT(64'b0111110011010010000011000001111000011010110101111000011001110000)  
) LUT6_272 (
   .O(gates[1149]),
   .I0(InputBits[537]),
   .I1(InputBits[1413]),
   .I2(InputBits[944]),
   .I3(InputBits[901]),
   .I4(InputBits[1636]),
   .I5(InputBits[1250])
);
LUT6 #(
   .INIT(64'b1011010101000010001000010101111101011101100010100111011001000001)  
) LUT6_273 (
   .O(gates[542]),
   .I0(InputBits[541]),
   .I1(InputBits[229]),
   .I2(InputBits[1284]),
   .I3(InputBits[124]),
   .I4(InputBits[594]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b1001010110101000001111101001110110110111100100000001010010001010)  
) LUT6_274 (
   .O(gates[1305]),
   .I0(InputBits[1462]),
   .I1(InputBits[1085]),
   .I2(InputBits[65]),
   .I3(InputBits[1145]),
   .I4(InputBits[686]),
   .I5(InputBits[1549])
);
LUT6 #(
   .INIT(64'b0100110011000111010010110011110100011111111111111011111111110010)  
) LUT6_275 (
   .O(gates[961]),
   .I0(InputBits[1420]),
   .I1(InputBits[1505]),
   .I2(InputBits[1612]),
   .I3(InputBits[1192]),
   .I4(InputBits[328]),
   .I5(InputBits[607])
);
LUT6 #(
   .INIT(64'b1001001001100001101111101101100010100001010111001010110010100111)  
) LUT6_276 (
   .O(gates[1288]),
   .I0(InputBits[815]),
   .I1(InputBits[291]),
   .I2(InputBits[660]),
   .I3(InputBits[1116]),
   .I4(InputBits[370]),
   .I5(InputBits[999])
);
LUT6 #(
   .INIT(64'b0000000001010011011001110101001000101011101100101000111010001010)  
) LUT6_277 (
   .O(gates[1087]),
   .I0(InputBits[1019]),
   .I1(InputBits[1361]),
   .I2(InputBits[1571]),
   .I3(InputBits[1045]),
   .I4(InputBits[960]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b1011100011101000011100110011010100111000111001101010110101111001)  
) LUT6_278 (
   .O(gates[810]),
   .I0(InputBits[28]),
   .I1(InputBits[862]),
   .I2(InputBits[76]),
   .I3(InputBits[273]),
   .I4(InputBits[1050]),
   .I5(InputBits[1065])
);
LUT6 #(
   .INIT(64'b0011001110001011110100111110100110100100101011101100011111111111)  
) LUT6_279 (
   .O(gates[574]),
   .I0(InputBits[739]),
   .I1(InputBits[1451]),
   .I2(InputBits[583]),
   .I3(InputBits[965]),
   .I4(InputBits[892]),
   .I5(InputBits[670])
);
LUT6 #(
   .INIT(64'b1011001010000001101000111000100000001111111001000100111000010111)  
) LUT6_280 (
   .O(gates[1238]),
   .I0(InputBits[23]),
   .I1(InputBits[1673]),
   .I2(InputBits[1585]),
   .I3(InputBits[1488]),
   .I4(InputBits[1063]),
   .I5(InputBits[1426])
);
LUT6 #(
   .INIT(64'b0110001011010011011001101111101010000111111111111101110101001100)  
) LUT6_281 (
   .O(gates[170]),
   .I0(InputBits[1483]),
   .I1(InputBits[596]),
   .I2(InputBits[1238]),
   .I3(InputBits[274]),
   .I4(InputBits[362]),
   .I5(InputBits[1033])
);
LUT6 #(
   .INIT(64'b0100101101111001101101010110000010001010111011011011010101010110)  
) LUT6_282 (
   .O(gates[33]),
   .I0(InputBits[1438]),
   .I1(InputBits[349]),
   .I2(InputBits[206]),
   .I3(InputBits[74]),
   .I4(InputBits[363]),
   .I5(InputBits[1200])
);
LUT6 #(
   .INIT(64'b1110111001110101011001111100000011110001010011011101110001000001)  
) LUT6_283 (
   .O(gates[660]),
   .I0(InputBits[641]),
   .I1(InputBits[147]),
   .I2(InputBits[1682]),
   .I3(InputBits[1563]),
   .I4(InputBits[158]),
   .I5(InputBits[1595])
);
LUT6 #(
   .INIT(64'b1010001011110001011011000010010010011111010010110010011101010000)  
) LUT6_284 (
   .O(gates[7]),
   .I0(InputBits[1107]),
   .I1(InputBits[865]),
   .I2(InputBits[1174]),
   .I3(InputBits[549]),
   .I4(InputBits[1609]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1010111111101101000000100110111010001011101011110101011101100010)  
) LUT6_285 (
   .O(gates[227]),
   .I0(InputBits[1339]),
   .I1(InputBits[1303]),
   .I2(InputBits[174]),
   .I3(InputBits[971]),
   .I4(InputBits[1330]),
   .I5(InputBits[1306])
);
LUT6 #(
   .INIT(64'b0010101100011111100011000100000111100110111100001111000010011110)  
) LUT6_286 (
   .O(gates[26]),
   .I0(InputBits[933]),
   .I1(InputBits[1551]),
   .I2(InputBits[1017]),
   .I3(InputBits[219]),
   .I4(InputBits[932]),
   .I5(InputBits[1633])
);
LUT6 #(
   .INIT(64'b1110010011011111101000000001010000001100010000110110111010100011)  
) LUT6_287 (
   .O(gates[977]),
   .I0(InputBits[1647]),
   .I1(InputBits[841]),
   .I2(InputBits[164]),
   .I3(InputBits[1165]),
   .I4(InputBits[1161]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b1010101001100110100100110110010011011011011001101100010110010110)  
) LUT6_288 (
   .O(gates[566]),
   .I0(InputBits[508]),
   .I1(InputBits[1114]),
   .I2(InputBits[136]),
   .I3(InputBits[448]),
   .I4(InputBits[1714]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0001011101010100000100110001100011000010000011111110011000111100)  
) LUT6_289 (
   .O(gates[526]),
   .I0(InputBits[1077]),
   .I1(InputBits[1123]),
   .I2(InputBits[246]),
   .I3(InputBits[93]),
   .I4(InputBits[1343]),
   .I5(InputBits[1519])
);
LUT6 #(
   .INIT(64'b0010111010001110011000111100010111001001110000001101010111001000)  
) LUT6_290 (
   .O(gates[806]),
   .I0(InputBits[1372]),
   .I1(InputBits[1257]),
   .I2(InputBits[711]),
   .I3(InputBits[1608]),
   .I4(InputBits[1275]),
   .I5(InputBits[1360])
);
LUT6 #(
   .INIT(64'b0110011110010000010000100110000001001100000001010101001001101011)  
) LUT6_291 (
   .O(gates[264]),
   .I0(InputBits[1170]),
   .I1(InputBits[377]),
   .I2(InputBits[1387]),
   .I3(InputBits[961]),
   .I4(InputBits[1061]),
   .I5(InputBits[1079])
);
LUT6 #(
   .INIT(64'b1111010101100011000001000010011010000010110111000100111100100001)  
) LUT6_292 (
   .O(gates[255]),
   .I0(InputBits[230]),
   .I1(InputBits[1584]),
   .I2(InputBits[983]),
   .I3(InputBits[893]),
   .I4(InputBits[1414]),
   .I5(InputBits[952])
);
LUT6 #(
   .INIT(64'b1000000101110100101100011000010110101111100100110110111101110001)  
) LUT6_293 (
   .O(gates[359]),
   .I0(InputBits[1166]),
   .I1(InputBits[1496]),
   .I2(InputBits[512]),
   .I3(InputBits[75]),
   .I4(InputBits[996]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1000110010011010000001101010000111100010011001100001011111001000)  
) LUT6_294 (
   .O(gates[182]),
   .I0(InputBits[1554]),
   .I1(InputBits[1630]),
   .I2(InputBits[599]),
   .I3(InputBits[83]),
   .I4(InputBits[589]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b1101100100111110000000010010101001010110110000011010010001000000)  
) LUT6_295 (
   .O(gates[1229]),
   .I0(InputBits[255]),
   .I1(InputBits[648]),
   .I2(InputBits[60]),
   .I3(InputBits[1582]),
   .I4(InputBits[1276]),
   .I5(InputBits[1510])
);
LUT6 #(
   .INIT(64'b0000011101110111100111101100011010010000000000001101011001011100)  
) LUT6_296 (
   .O(gates[108]),
   .I0(InputBits[1377]),
   .I1(InputBits[177]),
   .I2(InputBits[518]),
   .I3(InputBits[832]),
   .I4(InputBits[1199]),
   .I5(InputBits[851])
);
LUT6 #(
   .INIT(64'b1100011101011001011100011001100011001100101111100011000100111001)  
) LUT6_297 (
   .O(gates[604]),
   .I0(InputBits[1617]),
   .I1(InputBits[1439]),
   .I2(InputBits[369]),
   .I3(InputBits[1701]),
   .I4(InputBits[1163]),
   .I5(InputBits[1487])
);
LUT6 #(
   .INIT(64'b0010100010111000001010010100001010110101011001010111001000001011)  
) LUT6_298 (
   .O(gates[1001]),
   .I0(InputBits[1037]),
   .I1(InputBits[105]),
   .I2(InputBits[870]),
   .I3(InputBits[148]),
   .I4(InputBits[1652]),
   .I5(InputBits[735])
);
LUT6 #(
   .INIT(64'b0101011101100111100011111001101001101111011010100101101001101011)  
) LUT6_299 (
   .O(gates[556]),
   .I0(InputBits[759]),
   .I1(InputBits[531]),
   .I2(InputBits[661]),
   .I3(InputBits[261]),
   .I4(InputBits[905]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b0000100000100001111000001100011100110110110011010110111110101111)  
) LUT6_300 (
   .O(gates[717]),
   .I0(InputBits[1288]),
   .I1(InputBits[955]),
   .I2(InputBits[1144]),
   .I3(InputBits[790]),
   .I4(InputBits[903]),
   .I5(InputBits[1032])
);
LUT6 #(
   .INIT(64'b0010101100011010010111001111100100100000010011010000100011000111)  
) LUT6_301 (
   .O(gates[232]),
   .I0(InputBits[1569]),
   .I1(InputBits[53]),
   .I2(InputBits[773]),
   .I3(InputBits[1418]),
   .I4(InputBits[1012]),
   .I5(InputBits[1444])
);
LUT6 #(
   .INIT(64'b1011110011011001111110101110111110101010000101111001000000001011)  
) LUT6_302 (
   .O(gates[477]),
   .I0(InputBits[886]),
   .I1(InputBits[1421]),
   .I2(InputBits[919]),
   .I3(InputBits[1677]),
   .I4(InputBits[1334]),
   .I5(InputBits[859])
);
LUT6 #(
   .INIT(64'b1001000111001000101001110101001001110100000100011000100110000011)  
) LUT6_303 (
   .O(gates[815]),
   .I0(InputBits[1369]),
   .I1(InputBits[1683]),
   .I2(InputBits[348]),
   .I3(InputBits[719]),
   .I4(InputBits[639]),
   .I5(InputBits[730])
);
LUT6 #(
   .INIT(64'b0101100111111011001110001110111000100100111101101001001110001110)  
) LUT6_304 (
   .O(gates[671]),
   .I0(InputBits[1603]),
   .I1(InputBits[1537]),
   .I2(InputBits[447]),
   .I3(InputBits[1309]),
   .I4(InputBits[1212]),
   .I5(InputBits[633])
);
LUT6 #(
   .INIT(64'b0001001101111101011001110000011111010100101011100000011111000001)  
) LUT6_305 (
   .O(gates[1338]),
   .I0(InputBits[533]),
   .I1(InputBits[223]),
   .I2(InputBits[112]),
   .I3(InputBits[304]),
   .I4(InputBits[784]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b1111011011011011000111001111101000111000011110000011010101001011)  
) LUT6_306 (
   .O(gates[1511]),
   .I0(InputBits[579]),
   .I1(InputBits[1561]),
   .I2(InputBits[1221]),
   .I3(InputBits[804]),
   .I4(InputBits[1684]),
   .I5(InputBits[1346])
);
LUT6 #(
   .INIT(64'b0100001001001100011111011011101001001101000111011011001010100010)  
) LUT6_307 (
   .O(gates[1182]),
   .I0(InputBits[1556]),
   .I1(InputBits[879]),
   .I2(InputBits[490]),
   .I3(InputBits[1594]),
   .I4(InputBits[1027]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b0110001010000001111001010100101000011110010000001011111100111111)  
) LUT6_308 (
   .O(gates[225]),
   .I0(InputBits[478]),
   .I1(InputBits[499]),
   .I2(InputBits[173]),
   .I3(InputBits[1230]),
   .I4(InputBits[1669]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b0100101100100110010111101101011111111100100010000001000011101001)  
) LUT6_309 (
   .O(gates[330]),
   .I0(InputBits[1121]),
   .I1(InputBits[1352]),
   .I2(InputBits[1315]),
   .I3(InputBits[30]),
   .I4(InputBits[322]),
   .I5(InputBits[1384])
);
LUT6 #(
   .INIT(64'b0000111011000001111100001110111010010111001011011110011101111011)  
) LUT6_310 (
   .O(gates[142]),
   .I0(InputBits[1304]),
   .I1(InputBits[1150]),
   .I2(InputBits[1638]),
   .I3(InputBits[672]),
   .I4(InputBits[1686]),
   .I5(InputBits[1464])
);
LUT6 #(
   .INIT(64'b0011010001000010011101000000111000101011011110100001101000110111)  
) LUT6_311 (
   .O(gates[1447]),
   .I0(InputBits[614]),
   .I1(InputBits[1703]),
   .I2(InputBits[186]),
   .I3(InputBits[212]),
   .I4(InputBits[563]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b0000111011011100110111001111011001100001110111000010000110000101)  
) LUT6_312 (
   .O(gates[207]),
   .I0(InputBits[682]),
   .I1(InputBits[133]),
   .I2(InputBits[839]),
   .I3(InputBits[1042]),
   .I4(InputBits[775]),
   .I5(InputBits[1294])
);
LUT6 #(
   .INIT(64'b0010001001101100101001010000110111010001111110101100000011111100)  
) LUT6_313 (
   .O(gates[1510]),
   .I0(InputBits[316]),
   .I1(InputBits[1099]),
   .I2(InputBits[830]),
   .I3(InputBits[1403]),
   .I4(InputBits[277]),
   .I5(InputBits[1240])
);
LUT6 #(
   .INIT(64'b1010100001011101111111111001111100011111011101011010001100000101)  
) LUT6_314 (
   .O(gates[167]),
   .I0(InputBits[1149]),
   .I1(InputBits[1592]),
   .I2(InputBits[1621]),
   .I3(InputBits[1705]),
   .I4(InputBits[5]),
   .I5(InputBits[1645])
);
LUT6 #(
   .INIT(64'b1100110011111000000101010011100101101010101010111011110101101101)  
) LUT6_315 (
   .O(gates[48]),
   .I0(InputBits[1481]),
   .I1(InputBits[207]),
   .I2(InputBits[613]),
   .I3(InputBits[1525]),
   .I4(InputBits[506]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0010001010110110011111100011000100110001110010010101101111100100)  
) LUT6_316 (
   .O(gates[360]),
   .I0(InputBits[1155]),
   .I1(InputBits[949]),
   .I2(InputBits[1243]),
   .I3(InputBits[1397]),
   .I4(InputBits[795]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b0001100000010101100000100001011001110101101101010110000101101101)  
) LUT6_317 (
   .O(gates[692]),
   .I0(InputBits[924]),
   .I1(InputBits[1066]),
   .I2(InputBits[1663]),
   .I3(InputBits[492]),
   .I4(InputBits[25]),
   .I5(InputBits[1719])
);
LUT6 #(
   .INIT(64'b1011111001110001010110100001001001000010111101110000111001111110)  
) LUT6_318 (
   .O(gates[663]),
   .I0(InputBits[1382]),
   .I1(InputBits[864]),
   .I2(InputBits[591]),
   .I3(InputBits[1602]),
   .I4(InputBits[1290]),
   .I5(InputBits[969])
);
LUT6 #(
   .INIT(64'b1100010011000111011011101000011101000010101100010111010100100010)  
) LUT6_319 (
   .O(gates[854]),
   .I0(InputBits[927]),
   .I1(InputBits[380]),
   .I2(InputBits[1164]),
   .I3(InputBits[1135]),
   .I4(InputBits[259]),
   .I5(InputBits[1172])
);
LUT6 #(
   .INIT(64'b0101010110011000011000010000101010100011001010101011010101111110)  
) LUT6_320 (
   .O(gates[969]),
   .I0(InputBits[650]),
   .I1(InputBits[1411]),
   .I2(InputBits[658]),
   .I3(InputBits[1253]),
   .I4(InputBits[523]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b1111000000010100110001100101101000011101000000100000000010100001)  
) LUT6_321 (
   .O(gates[1174]),
   .I0(InputBits[1470]),
   .I1(InputBits[1449]),
   .I2(InputBits[1385]),
   .I3(InputBits[1517]),
   .I4(InputBits[418]),
   .I5(InputBits[1355])
);
LUT6 #(
   .INIT(64'b1101011111000010100011110101010001000011000001101100010001111000)  
) LUT6_322 (
   .O(gates[1076]),
   .I0(InputBits[436]),
   .I1(InputBits[1472]),
   .I2(InputBits[197]),
   .I3(InputBits[21]),
   .I4(InputBits[1658]),
   .I5(InputBits[1625])
);
LUT6 #(
   .INIT(64'b0110101100110111010110111000111000011001010101111111111101010111)  
) LUT6_323 (
   .O(gates[510]),
   .I0(InputBits[747]),
   .I1(InputBits[1319]),
   .I2(InputBits[1126]),
   .I3(InputBits[203]),
   .I4(InputBits[67]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0011101011011100011111001011101100111001011100110010110101110110)  
) LUT6_324 (
   .O(gates[766]),
   .I0(InputBits[1190]),
   .I1(InputBits[1508]),
   .I2(InputBits[153]),
   .I3(InputBits[665]),
   .I4(InputBits[356]),
   .I5(InputBits[1301])
);
LUT6 #(
   .INIT(64'b0101110011111110010100111111010100100101111010101110010101011011)  
) LUT6_325 (
   .O(gates[393]),
   .I0(InputBits[973]),
   .I1(InputBits[36]),
   .I2(InputBits[122]),
   .I3(InputBits[1181]),
   .I4(InputBits[479]),
   .I5(InputBits[644])
);
LUT6 #(
   .INIT(64'b1001001010111101010101010101001010011010101111101110101111111101)  
) LUT6_326 (
   .O(gates[449]),
   .I0(InputBits[845]),
   .I1(InputBits[703]),
   .I2(InputBits[619]),
   .I3(InputBits[474]),
   .I4(InputBits[794]),
   .I5(InputBits[1447])
);
LUT6 #(
   .INIT(64'b1111111111000101011100010000101100011110001111100100010100100100)  
) LUT6_327 (
   .O(gates[1501]),
   .I0(InputBits[1197]),
   .I1(InputBits[1168]),
   .I2(InputBits[1558]),
   .I3(InputBits[438]),
   .I4(InputBits[338]),
   .I5(InputBits[91])
);
LUT6 #(
   .INIT(64'b1101001111011000001100110011101010100110110111001010110100100111)  
) LUT6_328 (
   .O(gates[658]),
   .I0(InputBits[788]),
   .I1(InputBits[1455]),
   .I2(InputBits[963]),
   .I3(InputBits[1489]),
   .I4(InputBits[553]),
   .I5(InputBits[821])
);
LUT6 #(
   .INIT(64'b1000001001101110011101010010100100001111110110000000011001000000)  
) LUT6_329 (
   .O(gates[274]),
   .I0(InputBits[428]),
   .I1(InputBits[1545]),
   .I2(InputBits[468]),
   .I3(InputBits[422]),
   .I4(InputBits[199]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b1101100101110000100010010100111101111001011110111111010000011001)  
) LUT6_330 (
   .O(gates[549]),
   .I0(InputBits[270]),
   .I1(InputBits[114]),
   .I2(InputBits[397]),
   .I3(InputBits[538]),
   .I4(InputBits[1475]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0111110000100001101000111001000110100000110111000100101100101100)  
) LUT6_331 (
   .O(gates[659]),
   .I0(InputBits[1298]),
   .I1(InputBits[1040]),
   .I2(InputBits[59]),
   .I3(InputBits[663]),
   .I4(InputBits[761]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0001111001011001111110000001001001100101111111110011001111111110)  
) LUT6_332 (
   .O(gates[877]),
   .I0(InputBits[404]),
   .I1(InputBits[520]),
   .I2(InputBits[426]),
   .I3(InputBits[1696]),
   .I4(InputBits[990]),
   .I5(InputBits[1206])
);
LUT6 #(
   .INIT(64'b1011000001101110000110101001011011011100001101100001011101100110)  
) LUT6_333 (
   .O(gates[1508]),
   .I0(InputBits[1441]),
   .I1(InputBits[319]),
   .I2(InputBits[1650]),
   .I3(InputBits[526]),
   .I4(InputBits[248]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b0011110100100001011000011110101011111000010100101101010001011100)  
) LUT6_334 (
   .O(gates[1141]),
   .I0(InputBits[967]),
   .I1(InputBits[753]),
   .I2(InputBits[12]),
   .I3(InputBits[896]),
   .I4(InputBits[221]),
   .I5(InputBits[1010])
);
LUT6 #(
   .INIT(64'b1101110100001111001011110000010011100001110001101000010011110011)  
) LUT6_335 (
   .O(gates[1128]),
   .I0(InputBits[603]),
   .I1(InputBits[1492]),
   .I2(InputBits[1021]),
   .I3(InputBits[637]),
   .I4(InputBits[1112]),
   .I5(InputBits[807])
);
LUT6 #(
   .INIT(64'b1001011110101110111110010010000001100010111111011101101000001001)  
) LUT6_336 (
   .O(gates[682]),
   .I0(InputBits[860]),
   .I1(InputBits[1028]),
   .I2(InputBits[1241]),
   .I3(InputBits[1034]),
   .I4(InputBits[440]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b1011010000100111110101011101011001110000111000101101100000110101)  
) LUT6_337 (
   .O(gates[353]),
   .I0(InputBits[1259]),
   .I1(InputBits[801]),
   .I2(InputBits[101]),
   .I3(InputBits[279]),
   .I4(InputBits[587]),
   .I5(InputBits[655])
);
LUT6 #(
   .INIT(64'b0000111001101001110110010011110110100000000111001101010011001010)  
) LUT6_338 (
   .O(gates[375]),
   .I0(InputBits[109]),
   .I1(InputBits[1656]),
   .I2(InputBits[1103]),
   .I3(InputBits[1178]),
   .I4(InputBits[912]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b1000110100011101101011010000101001111100101011101100111111001111)  
) LUT6_339 (
   .O(gates[984]),
   .I0(InputBits[1225]),
   .I1(InputBits[771]),
   .I2(InputBits[626]),
   .I3(InputBits[389]),
   .I4(InputBits[1534]),
   .I5(InputBits[674])
);
LUT6 #(
   .INIT(64'b1110010101000000010010100101110000011111010011011100111100111101)  
) LUT6_340 (
   .O(gates[1155]),
   .I0(InputBits[27]),
   .I1(InputBits[881]),
   .I2(InputBits[1287]),
   .I3(InputBits[44]),
   .I4(InputBits[1458]),
   .I5(InputBits[751])
);
LUT6 #(
   .INIT(64'b0001111010110010001111110100000111011011000110011110011001101100)  
) LUT6_341 (
   .O(gates[946]),
   .I0(InputBits[1345]),
   .I1(InputBits[1035]),
   .I2(InputBits[828]),
   .I3(InputBits[1559]),
   .I4(InputBits[1097]),
   .I5(InputBits[782])
);
LUT6 #(
   .INIT(64'b1000000101011101001111011101110100111101101101000011011010111111)  
) LUT6_342 (
   .O(gates[1485]),
   .I0(InputBits[728]),
   .I1(InputBits[1048]),
   .I2(InputBits[688]),
   .I3(InputBits[1131]),
   .I4(InputBits[852]),
   .I5(InputBits[1327])
);
LUT6 #(
   .INIT(64'b1011100000111111100101010011001111111111001100100111111100111100)  
) LUT6_343 (
   .O(gates[788]),
   .I0(InputBits[1679]),
   .I1(InputBits[107]),
   .I2(InputBits[544]),
   .I3(InputBits[1140]),
   .I4(InputBits[921]),
   .I5(InputBits[1433])
);
LUT6 #(
   .INIT(64'b0101000101001100100000101001001100000001001010000101011000100101)  
) LUT6_344 (
   .O(gates[128]),
   .I0(InputBits[32]),
   .I1(InputBits[366]),
   .I2(InputBits[4]),
   .I3(InputBits[1311]),
   .I4(InputBits[1662]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1100101100001001100011101011110001111111111110000101101111111000)  
) LUT6_345 (
   .O(gates[1520]),
   .I0(InputBits[146]),
   .I1(InputBits[305]),
   .I2(InputBits[561]),
   .I3(InputBits[888]),
   .I4(InputBits[695]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b1100100101001110000011000101001011110000011000110000010101101001)  
) LUT6_346 (
   .O(gates[303]),
   .I0(InputBits[346]),
   .I1(InputBits[382]),
   .I2(InputBits[675]),
   .I3(InputBits[330]),
   .I4(InputBits[1210]),
   .I5(InputBits[1350])
);
LUT6 #(
   .INIT(64'b0000111100011101001110111010011111100100101100000101100101000111)  
) LUT6_347 (
   .O(gates[250]),
   .I0(InputBits[262]),
   .I1(InputBits[744]),
   .I2(InputBits[1265]),
   .I3(InputBits[1053]),
   .I4(InputBits[1059]),
   .I5(InputBits[1152])
);
LUT6 #(
   .INIT(64'b1010000000001010010101011100010001101011110110010101110001110101)  
) LUT6_348 (
   .O(gates[1361]),
   .I0(InputBits[1262]),
   .I1(InputBits[1499]),
   .I2(InputBits[1068]),
   .I3(InputBits[694]),
   .I4(InputBits[302]),
   .I5(InputBits[868])
);
LUT6 #(
   .INIT(64'b1010001111110011001101011110110010101111000001010010010010111010)  
) LUT6_349 (
   .O(gates[614]),
   .I0(InputBits[50]),
   .I1(InputBits[352]),
   .I2(InputBits[876]),
   .I3(InputBits[1615]),
   .I4(InputBits[390]),
   .I5(InputBits[1605])
);
LUT6 #(
   .INIT(64'b1101000001110101010010110111010000010110100010100001111101001001)  
) LUT6_350 (
   .O(gates[501]),
   .I0(InputBits[1565]),
   .I1(InputBits[1724]),
   .I2(InputBits[766]),
   .I3(InputBits[433]),
   .I4(InputBits[1580]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0110000011011101011111110010110110000010110111011000110000111100)  
) LUT6_351 (
   .O(gates[1313]),
   .I0(InputBits[1527]),
   .I1(InputBits[1465]),
   .I2(InputBits[721]),
   .I3(InputBits[1707]),
   .I4(InputBits[19]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1111001111010001011010001110010100100100010110011100100111010001)  
) LUT6_352 (
   .O(gates[278]),
   .I0(InputBits[1219]),
   .I1(InputBits[1479]),
   .I2(InputBits[1208]),
   .I3(InputBits[216]),
   .I4(InputBits[1416]),
   .I5(InputBits[1434])
);
LUT6 #(
   .INIT(64'b1111110101010000001100110010010001001100101001011100010111110001)  
) LUT6_353 (
   .O(gates[490]),
   .I0(InputBits[1336]),
   .I1(InputBits[854]),
   .I2(InputBits[1278]),
   .I3(InputBits[169]),
   .I4(InputBits[1089]),
   .I5(InputBits[593])
);
LUT6 #(
   .INIT(64'b1000011010100100001001010011100111100110010011100010101110011110)  
) LUT6_354 (
   .O(gates[155]),
   .I0(InputBits[210]),
   .I1(InputBits[1408]),
   .I2(InputBits[1600]),
   .I3(InputBits[1389]),
   .I4(InputBits[1404]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b0010010100111000111000000010110110000000100100111111010001001000)  
) LUT6_355 (
   .O(gates[130]),
   .I0(InputBits[1589]),
   .I1(InputBits[1095]),
   .I2(InputBits[288]),
   .I3(InputBits[1725]),
   .I4(InputBits[1370]),
   .I5(InputBits[1435])
);
LUT6 #(
   .INIT(64'b0000011110101011101100010000110001100111011011110100000001100101)  
) LUT6_356 (
   .O(gates[53]),
   .I0(InputBits[1071]),
   .I1(InputBits[358]),
   .I2(InputBits[684]),
   .I3(InputBits[1474]),
   .I4(InputBits[1157]),
   .I5(InputBits[837])
);
LUT6 #(
   .INIT(64'b0000010010100110101101010110110011011111010000000000001000011001)  
) LUT6_357 (
   .O(gates[387]),
   .I0(InputBits[7]),
   .I1(InputBits[324]),
   .I2(InputBits[269]),
   .I3(InputBits[645]),
   .I4(InputBits[726]),
   .I5(InputBits[1362])
);
LUT6 #(
   .INIT(64'b0011100100111101000100111000011000011101000001011100101100100000)  
) LUT6_358 (
   .O(gates[1373]),
   .I0(InputBits[2]),
   .I1(InputBits[314]),
   .I2(InputBits[1635]),
   .I3(InputBits[1502]),
   .I4(InputBits[787]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b1011110100100111010100011101011000111011111011100101101001001111)  
) LUT6_359 (
   .O(gates[1465]),
   .I0(InputBits[749]),
   .I1(InputBits[1321]),
   .I2(InputBits[786]),
   .I3(InputBits[580]),
   .I4(InputBits[1249]),
   .I5(InputBits[1292])
);
LUT6 #(
   .INIT(64'b0110111000111010111010100111000100000101101011001010001010110011)  
) LUT6_360 (
   .O(gates[1302]),
   .I0(InputBits[1678]),
   .I1(InputBits[1460]),
   .I2(InputBits[365]),
   .I3(InputBits[276]),
   .I4(InputBits[910]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1001011101001111100011011110001010010011111101010010001000010101)  
) LUT6_361 (
   .O(gates[1112]),
   .I0(InputBits[1310]),
   .I1(InputBits[143]),
   .I2(InputBits[1227]),
   .I3(InputBits[1437]),
   .I4(InputBits[482]),
   .I5(InputBits[1084])
);
LUT6 #(
   .INIT(64'b0110101101101000011100001000100101001010100010011001101010001001)  
) LUT6_362 (
   .O(gates[626]),
   .I0(InputBits[900]),
   .I1(InputBits[843]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[1087]),
   .I5(InputBits[799])
);
LUT6 #(
   .INIT(64'b0101110101010000001001100101101111011011111101111000101001001011)  
) LUT6_363 (
   .O(gates[1397]),
   .I0(InputBits[70]),
   .I1(InputBits[281]),
   .I2(InputBits[1431]),
   .I3(InputBits[847]),
   .I4(InputBits[1176]),
   .I5(InputBits[1374])
);
LUT6 #(
   .INIT(64'b0111100110111011010100001011001101101000001011110100111010001110)  
) LUT6_364 (
   .O(gates[1294]),
   .I0(InputBits[740]),
   .I1(InputBits[898]),
   .I2(InputBits[286]),
   .I3(InputBits[327]),
   .I4(InputBits[1272]),
   .I5(InputBits[1183])
);
LUT6 #(
   .INIT(64'b0001111000110110000011101110111011110100101011101001010111010000)  
) LUT6_365 (
   .O(gates[941]),
   .I0(InputBits[1466]),
   .I1(InputBits[1031]),
   .I2(InputBits[1203]),
   .I3(InputBits[1610]),
   .I4(InputBits[978]),
   .I5(InputBits[1215])
);
LUT6 #(
   .INIT(64'b1110000101100010001000001000111010110001000101001110001100111010)  
) LUT6_366 (
   .O(gates[461]),
   .I0(InputBits[1086]),
   .I1(InputBits[1115]),
   .I2(InputBits[1532]),
   .I3(InputBits[1452]),
   .I4(InputBits[29]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b1111100110110111100001100010011001100110010111101100000000001101)  
) LUT6_367 (
   .O(gates[583]),
   .I0(InputBits[22]),
   .I1(InputBits[601]),
   .I2(InputBits[17]),
   .I3(InputBits[1296]),
   .I4(InputBits[1417]),
   .I5(InputBits[1574])
);
LUT6 #(
   .INIT(64'b1111101100111001101111111000000100100110111110011101000001010111)  
) LUT6_368 (
   .O(gates[1426]),
   .I0(InputBits[595]),
   .I1(InputBits[451]),
   .I2(InputBits[690]),
   .I3(InputBits[1623]),
   .I4(InputBits[1280]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b1101100000011001001111000010111111010101011001010011100010110010)  
) LUT6_369 (
   .O(gates[257]),
   .I0(InputBits[1314]),
   .I1(InputBits[575]),
   .I2(InputBits[353]),
   .I3(InputBits[170]),
   .I4(InputBits[34]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b1001001110010100101010111101001100111000000101000010110111110001)  
) LUT6_370 (
   .O(gates[1358]),
   .I0(InputBits[995]),
   .I1(InputBits[1237]),
   .I2(InputBits[824]),
   .I3(InputBits[1128]),
   .I4(InputBits[1688]),
   .I5(InputBits[1448])
);
LUT6 #(
   .INIT(64'b1100001110000100111001111010100111110111110100010100010110010100)  
) LUT6_371 (
   .O(gates[782]),
   .I0(InputBits[1064]),
   .I1(InputBits[464]),
   .I2(InputBits[115]),
   .I3(InputBits[455]),
   .I4(InputBits[1110]),
   .I5(InputBits[1279])
);
LUT6 #(
   .INIT(64'b0010110111010101000011011111000100011100111100101101110111000110)  
) LUT6_372 (
   .O(gates[951]),
   .I0(InputBits[57]),
   .I1(InputBits[913]),
   .I2(InputBits[1727]),
   .I3(InputBits[193]),
   .I4(InputBits[572]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1101010011000001110110100100111101110101001001111000000110010110)  
) LUT6_373 (
   .O(gates[85]),
   .I0(InputBits[628]),
   .I1(InputBits[667]),
   .I2(InputBits[15]),
   .I3(InputBits[1118]),
   .I4(InputBits[345]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b1100000011000111101101000000111111010011100101100010001010011101)  
) LUT6_374 (
   .O(gates[809]),
   .I0(InputBits[1023]),
   .I1(InputBits[116]),
   .I2(InputBits[486]),
   .I3(InputBits[507]),
   .I4(InputBits[1338]),
   .I5(InputBits[1596])
);
LUT6 #(
   .INIT(64'b1011001100010001111101100110110001111101110001001001010110000110)  
) LUT6_375 (
   .O(gates[1156]),
   .I0(InputBits[1506]),
   .I1(InputBits[1246]),
   .I2(InputBits[8]),
   .I3(InputBits[1536]),
   .I4(InputBits[611]),
   .I5(InputBits[1331])
);
LUT6 #(
   .INIT(64'b0000000111011000100110001100100100100111011100000100110010101100)  
) LUT6_376 (
   .O(gates[425]),
   .I0(InputBits[988]),
   .I1(InputBits[245]),
   .I2(InputBits[1266]),
   .I3(InputBits[546]),
   .I4(InputBits[162]),
   .I5(InputBits[1507])
);
LUT6 #(
   .INIT(64'b1101111110110001000101010010100111110100010101100010101111000110)  
) LUT6_377 (
   .O(gates[1486]),
   .I0(InputBits[1002]),
   .I1(InputBits[1160]),
   .I2(InputBits[550]),
   .I3(InputBits[79]),
   .I4(InputBits[1139]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1110111111000010001010100001111000011001110110111100101011011000)  
) LUT6_378 (
   .O(gates[591]),
   .I0(InputBits[293]),
   .I1(InputBits[621]),
   .I2(InputBits[1236]),
   .I3(InputBits[1159]),
   .I4(InputBits[1102]),
   .I5(InputBits[755])
);
LUT6 #(
   .INIT(64'b0010100111100110111001000111100010000011111001011010011011101001)  
) LUT6_379 (
   .O(gates[832]),
   .I0(InputBits[312]),
   .I1(InputBits[940]),
   .I2(InputBits[931]),
   .I3(InputBits[1497]),
   .I4(InputBits[767]),
   .I5(InputBits[883])
);
LUT6 #(
   .INIT(64'b0111011101001111010111101100000010110010111110010011110111100000)  
) LUT6_380 (
   .O(gates[736]),
   .I0(InputBits[762]),
   .I1(InputBits[1722]),
   .I2(InputBits[68]),
   .I3(InputBits[1691]),
   .I4(InputBits[950]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b1110101100111000011000001001111110101101001111010101011111010111)  
) LUT6_381 (
   .O(gates[539]),
   .I0(InputBits[1381]),
   .I1(InputBits[654]),
   .I2(InputBits[371]),
   .I3(InputBits[469]),
   .I4(InputBits[819]),
   .I5(InputBits[970])
);
LUT6 #(
   .INIT(64'b0100001010111001110001110010011001000110100011110011100011000100)  
) LUT6_382 (
   .O(gates[781]),
   .I0(InputBits[495]),
   .I1(InputBits[139]),
   .I2(InputBits[343]),
   .I3(InputBits[764]),
   .I4(InputBits[1186]),
   .I5(InputBits[1073])
);
LUT6 #(
   .INIT(64'b1011110101001011001010010100110010110111010010001010001111110110)  
) LUT6_383 (
   .O(gates[828]),
   .I0(InputBits[915]),
   .I1(InputBits[232]),
   .I2(InputBits[1217]),
   .I3(InputBits[196]),
   .I4(InputBits[696]),
   .I5(InputBits[582])
);
LUT6 #(
   .INIT(64'b0010100000111100001001101011001100011100000101001111100000110010)  
) LUT6_384 (
   .O(gates[276]),
   .I0(InputBits[1628]),
   .I1(InputBits[1260]),
   .I2(InputBits[1524]),
   .I3(InputBits[1239]),
   .I4(InputBits[566]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b1010001110010011101111010000110001100100101001100111100101001111)  
) LUT6_385 (
   .O(gates[102]),
   .I0(InputBits[1515]),
   .I1(InputBits[1153]),
   .I2(InputBits[1007]),
   .I3(InputBits[95]),
   .I4(InputBits[1196]),
   .I5(InputBits[1539])
);
LUT6 #(
   .INIT(64'b0011100110001111000101001110111100010110000000001110011001010000)  
) LUT6_386 (
   .O(gates[520]),
   .I0(InputBits[1234]),
   .I1(InputBits[519]),
   .I2(InputBits[984]),
   .I3(InputBits[1295]),
   .I4(InputBits[992]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0111000100101111011000010000000000001110111010001110010010100110)  
) LUT6_387 (
   .O(gates[532]),
   .I0(InputBits[1224]),
   .I1(InputBits[1693]),
   .I2(InputBits[1364]),
   .I3(InputBits[1398]),
   .I4(InputBits[584]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0000011001110011101110010000001011011111100000000111101010111001)  
) LUT6_388 (
   .O(gates[1218]),
   .I0(InputBits[228]),
   .I1(InputBits[373]),
   .I2(InputBits[201]),
   .I3(InputBits[700]),
   .I4(InputBits[81]),
   .I5(InputBits[936])
);
LUT6 #(
   .INIT(64'b0000010001101111100100010101111001010011110101110011001010000110)  
) LUT6_389 (
   .O(gates[1193]),
   .I0(InputBits[504]),
   .I1(InputBits[272]),
   .I2(InputBits[959]),
   .I3(InputBits[811]),
   .I4(InputBits[946]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b1111101100101100000100111101011010111011011000111110100100011111)  
) LUT6_390 (
   .O(gates[55]),
   .I0(InputBits[1550]),
   .I1(InputBits[441]),
   .I2(InputBits[1356]),
   .I3(InputBits[715]),
   .I4(InputBits[220]),
   .I5(InputBits[863])
);
LUT6 #(
   .INIT(64'b0001111011110011001111101001101011100111000010011001011001011011)  
) LUT6_391 (
   .O(gates[1404]),
   .I0(InputBits[1577]),
   .I1(InputBits[779]),
   .I2(InputBits[975]),
   .I3(InputBits[510]),
   .I4(InputBits[1401]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b0010010010010111101110010011010101110110000100101000110001111110)  
) LUT6_392 (
   .O(gates[1543]),
   .I0(InputBits[1698]),
   .I1(InputBits[834]),
   .I2(InputBits[1009]),
   .I3(InputBits[1690]),
   .I4(InputBits[827]),
   .I5(InputBits[1391])
);
LUT6 #(
   .INIT(64'b1010111000011110110110000101010110000100010101110111101011010101)  
) LUT6_393 (
   .O(gates[57]),
   .I0(InputBits[1093]),
   .I1(InputBits[1080]),
   .I2(InputBits[175]),
   .I3(InputBits[722]),
   .I4(InputBits[798]),
   .I5(InputBits[296])
);
LUT6 #(
   .INIT(64'b1100010100100010100000000101011111011101001111010101011111011100)  
) LUT6_394 (
   .O(gates[259]),
   .I0(InputBits[1643]),
   .I1(InputBits[1660]),
   .I2(InputBits[1075]),
   .I3(InputBits[604]),
   .I4(InputBits[1504]),
   .I5(InputBits[818])
);
LUT6 #(
   .INIT(64'b1100001110100100000111001001001111110111110000100110010000010001)  
) LUT6_395 (
   .O(gates[424]),
   .I0(InputBits[708]),
   .I1(InputBits[100]),
   .I2(InputBits[388]),
   .I3(InputBits[1708]),
   .I4(InputBits[1318]),
   .I5(InputBits[236])
);
LUT6 #(
   .INIT(64'b1011101110100010010001101001011111001101001000110001101111100100)  
) LUT6_396 (
   .O(gates[872]),
   .I0(InputBits[87]),
   .I1(InputBits[94]),
   .I2(InputBits[671]),
   .I3(InputBits[1323]),
   .I4(InputBits[625]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0111000000110100000010010001100110001110010110111111011011001011)  
) LUT6_397 (
   .O(gates[163]),
   .I0(InputBits[1214]),
   .I1(InputBits[1193]),
   .I2(InputBits[243]),
   .I3(InputBits[980]),
   .I4(InputBits[77]),
   .I5(InputBits[857])
);
LUT6 #(
   .INIT(64'b1011101011011110011001101111010100001110111000101011000011110110)  
) LUT6_398 (
   .O(gates[1106]),
   .I0(InputBits[132]),
   .I1(InputBits[597]),
   .I2(InputBits[724]),
   .I3(InputBits[278]),
   .I4(InputBits[1587]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0100111010010001101100110000000000001111110110100111001110111000)  
) LUT6_399 (
   .O(gates[1402]),
   .I0(InputBits[1251]),
   .I1(InputBits[1564]),
   .I2(InputBits[1307]),
   .I3(InputBits[9]),
   .I4(InputBits[234]),
   .I5(InputBits[1477])
);
LUT6 #(
   .INIT(64'b1010100001011110001110000100110101001110010111101100110111111000)  
) LUT6_400 (
   .O(gates[395]),
   .I0(InputBits[685]),
   .I1(InputBits[462]),
   .I2(InputBits[1108]),
   .I3(InputBits[1637]),
   .I4(InputBits[521]),
   .I5(InputBits[1468])
);
LUT6 #(
   .INIT(64'b1100000111101001011111110000011100000010100001101111110001000001)  
) LUT6_401 (
   .O(gates[1146]),
   .I0(InputBits[1329]),
   .I1(InputBits[1106]),
   .I2(InputBits[283]),
   .I3(InputBits[218]),
   .I4(InputBits[1611]),
   .I5(InputBits[1018])
);
LUT6 #(
   .INIT(64'b0001011111100111001101101011110111110100011100101101011100110010)  
) LUT6_402 (
   .O(gates[89]),
   .I0(InputBits[1429]),
   .I1(InputBits[1522]),
   .I2(InputBits[1379]),
   .I3(InputBits[1305]),
   .I4(InputBits[102]),
   .I5(InputBits[1586])
);
LUT6 #(
   .INIT(64'b0001000101001111110010110011101000001011011101101010010110011001)  
) LUT6_403 (
   .O(gates[175]),
   .I0(InputBits[835]),
   .I1(InputBits[1454]),
   .I2(InputBits[630]),
   .I3(InputBits[1162]),
   .I4(InputBits[1025]),
   .I5(InputBits[1572])
);
LUT6 #(
   .INIT(64'b0110011000010110110111010000111101000000001111101000001101010110)  
) LUT6_404 (
   .O(gates[1531]),
   .I0(InputBits[796]),
   .I1(InputBits[564]),
   .I2(InputBits[198]),
   .I3(InputBits[1632]),
   .I4(InputBits[570]),
   .I5(InputBits[1133])
);
LUT6 #(
   .INIT(64'b1101110000000110111010011101011100101100110111010010001001011001)  
) LUT6_405 (
   .O(gates[584]),
   .I0(InputBits[292]),
   .I1(InputBits[998]),
   .I2(InputBits[242]),
   .I3(InputBits[1424]),
   .I4(InputBits[359]),
   .I5(InputBits[1715])
);
LUT6 #(
   .INIT(64'b0010001100101000101101111100110100110110001011000111011011101110)  
) LUT6_406 (
   .O(gates[988]),
   .I0(InputBits[891]),
   .I1(InputBits[1484]),
   .I2(InputBits[1014]),
   .I3(InputBits[1406]),
   .I4(InputBits[364]),
   .I5(InputBits[1201])
);
LUT6 #(
   .INIT(64'b0110011000101110000000001111011011110100000111101110000101101111)  
) LUT6_407 (
   .O(gates[35]),
   .I0(InputBits[150]),
   .I1(InputBits[383]),
   .I2(InputBits[1445]),
   .I3(InputBits[540]),
   .I4(InputBits[1672]),
   .I5(InputBits[1046])
);
LUT6 #(
   .INIT(64'b0110100110101011010111110100100000111100000010100101111111000001)  
) LUT6_408 (
   .O(gates[1550]),
   .I0(InputBits[1044]),
   .I1(InputBits[1405]),
   .I2(InputBits[1552]),
   .I3(InputBits[1423]),
   .I4(InputBits[31]),
   .I5(InputBits[1016])
);
LUT6 #(
   .INIT(64'b0010110010111001011000111110111010010111100101010010011111110001)  
) LUT6_409 (
   .O(gates[1421]),
   .I0(InputBits[431]),
   .I1(InputBits[1302]),
   .I2(InputBits[1051]),
   .I3(InputBits[367]),
   .I4(InputBits[1493]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0111100001110111101000011101100011011010011010010110111010110000)  
) LUT6_410 (
   .O(gates[1454]),
   .I0(InputBits[258]),
   .I1(InputBits[1393]),
   .I2(InputBits[842]),
   .I3(InputBits[505]),
   .I4(InputBits[1074]),
   .I5(InputBits[113])
);
LUT6 #(
   .INIT(64'b0101010010001110111000110001111001010010110010010100111001100100)  
) LUT6_411 (
   .O(gates[347]),
   .I0(InputBits[160]),
   .I1(InputBits[742]),
   .I2(InputBits[608]),
   .I3(InputBits[659]),
   .I4(InputBits[58]),
   .I5(InputBits[1349])
);
LUT6 #(
   .INIT(64'b1101010101010001100010111111110001100011111010000110010001101011)  
) LUT6_412 (
   .O(gates[1333]),
   .I0(InputBits[548]),
   .I1(InputBits[1394]),
   .I2(InputBits[791]),
   .I3(InputBits[155]),
   .I4(InputBits[640]),
   .I5(InputBits[669])
);
LUT6 #(
   .INIT(64'b1000100001001100010010000101100000101111111000011001110010001000)  
) LUT6_413 (
   .O(gates[665]),
   .I0(InputBits[557]),
   .I1(InputBits[866]),
   .I2(InputBits[350]),
   .I3(InputBits[666]),
   .I4(InputBits[1282]),
   .I5(InputBits[1000])
);
LUT6 #(
   .INIT(64'b1110100011101011000100100100011011001111010111100111111100111001)  
) LUT6_414 (
   .O(gates[434]),
   .I0(InputBits[1648]),
   .I1(InputBits[1427]),
   .I2(InputBits[20]),
   .I3(InputBits[257]),
   .I4(InputBits[1681]),
   .I5(InputBits[873])
);
LUT6 #(
   .INIT(64'b0000100010010010011001111110001010010111000100000010011111001011)  
) LUT6_415 (
   .O(gates[1184]),
   .I0(InputBits[386]),
   .I1(InputBits[214]),
   .I2(InputBits[1271]),
   .I3(InputBits[652]),
   .I4(InputBits[920]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b0001001100000100011101101011010001110011110100011011001010111000)  
) LUT6_416 (
   .O(gates[1476]),
   .I0(InputBits[917]),
   .I1(InputBits[118]),
   .I2(InputBits[577]),
   .I3(InputBits[977]),
   .I4(InputBits[1626]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0011101011010101100000010111001101100001001000011001100100011111)  
) LUT6_417 (
   .O(gates[865]),
   .I0(InputBits[1057]),
   .I1(InputBits[166]),
   .I2(InputBits[942]),
   .I3(InputBits[624]),
   .I4(InputBits[617]),
   .I5(InputBits[476])
);
LUT6 #(
   .INIT(64'b0010011101100001111100100000011110101001010001100110111010011000)  
) LUT6_418 (
   .O(gates[1207]),
   .I0(InputBits[1495]),
   .I1(InputBits[717]),
   .I2(InputBits[334]),
   .I3(InputBits[1137]),
   .I4(InputBits[698]),
   .I5(InputBits[1091])
);
LUT6 #(
   .INIT(64'b0110001100001011100100100000001101100100011111111101011010100011)  
) LUT6_419 (
   .O(gates[904]),
   .I0(InputBits[878]),
   .I1(InputBits[41]),
   .I2(InputBits[1232]),
   .I3(InputBits[250]),
   .I4(InputBits[1671]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0111011110101110101000001100011011011111111111010001100100000101)  
) LUT6_420 (
   .O(gates[442]),
   .I0(InputBits[172]),
   .I1(InputBits[1367]),
   .I2(InputBits[542]),
   .I3(InputBits[1142]),
   .I4(InputBits[1269]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0001000110100011011010110100010011011101011011110010100100100111)  
) LUT6_421 (
   .O(gates[930]),
   .I0(InputBits[1184]),
   .I1(InputBits[181]),
   .I2(InputBits[14]),
   .I3(InputBits[623]),
   .I4(InputBits[460]),
   .I5(InputBits[1354])
);
LUT6 #(
   .INIT(64'b1010100010101101101110000011100010111101011110011011100111100101)  
) LUT6_422 (
   .O(gates[649]),
   .I0(InputBits[1653]),
   .I1(InputBits[987]),
   .I2(InputBits[423]),
   .I3(InputBits[568]),
   .I4(InputBits[809]),
   .I5(InputBits[734])
);
LUT6 #(
   .INIT(64'b0111010001110010100110101000011111011010111101101101010110000111)  
) LUT6_423 (
   .O(gates[689]),
   .I0(InputBits[1005]),
   .I1(InputBits[85]),
   .I2(InputBits[1728]),
   .I3(InputBits[757]),
   .I4(InputBits[1154]),
   .I5(InputBits[1512])
);
LUT6 #(
   .INIT(64'b0000010101101010001001001111000010101011010010011111110010111000)  
) LUT6_424 (
   .O(gates[886]),
   .I0(InputBits[1541]),
   .I1(InputBits[1120]),
   .I2(InputBits[1147]),
   .I3(InputBits[1175]),
   .I4(InputBits[1700]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1111000100010100101011001011110111100000111100100100001010000110)  
) LUT6_425 (
   .O(gates[1318]),
   .I0(InputBits[1038]),
   .I1(InputBits[1641]),
   .I2(InputBits[1575]),
   .I3(InputBits[466]),
   .I4(InputBits[805]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b0110011001110001011010000001101110101010010001011101000111101111)  
) LUT6_426 (
   .O(gates[642]),
   .I0(InputBits[1365]),
   .I1(InputBits[141]),
   .I2(InputBits[1613]),
   .I3(InputBits[848]),
   .I4(InputBits[483]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b1011010000110000010111001110011100010110111111011111100011110101)  
) LUT6_427 (
   .O(gates[648]),
   .I0(InputBits[1568]),
   .I1(InputBits[706]),
   .I2(InputBits[493]),
   .I3(InputBits[1555]),
   .I4(InputBits[536]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b1000000110000000100111101011111110011000110100010111000000011001)  
) LUT6_428 (
   .O(gates[1116]),
   .I0(InputBits[777]),
   .I1(InputBits[416]),
   .I2(InputBits[1375]),
   .I3(InputBits[803]),
   .I4(InputBits[943]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b1001000010001100010010100100000010101000101100000000001100010101)  
) LUT6_429 (
   .O(gates[1329]),
   .I0(InputBits[189]),
   .I1(InputBits[692]),
   .I2(InputBits[1619]),
   .I3(InputBits[1562]),
   .I4(InputBits[1312]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0111111010101111011110001110000011011011000010111100101010010000)  
) LUT6_430 (
   .O(gates[1028]),
   .I0(InputBits[1316]),
   .I1(InputBits[308]),
   .I2(InputBits[1720]),
   .I3(InputBits[1358]),
   .I4(InputBits[908]),
   .I5(InputBits[745])
);
LUT6 #(
   .INIT(64'b1111001010111011101000100110000111011110011001111001111111100001)  
) LUT6_431 (
   .O(gates[198]),
   .I0(InputBits[925]),
   .I1(InputBits[938]),
   .I2(InputBits[92]),
   .I3(InputBits[341]),
   .I4(InputBits[1340]),
   .I5(InputBits[825])
);
LUT6 #(
   .INIT(64'b1011001010001111001001010001111011010101110100100011110100100000)  
) LUT6_432 (
   .O(gates[1098]),
   .I0(InputBits[813]),
   .I1(InputBits[131]),
   .I2(InputBits[400]),
   .I3(InputBits[1710]),
   .I4(InputBits[1222]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0000100000010101011001101010100001010010000010110010100001000000)  
) LUT6_433 (
   .O(gates[1059]),
   .I0(InputBits[1229]),
   .I1(InputBits[119]),
   .I2(InputBits[1639]),
   .I3(InputBits[679]),
   .I4(InputBits[104]),
   .I5(InputBits[1191])
);
LUT6 #(
   .INIT(64'b1011000100010011100100000111110100110100010011000101011010101011)  
) LUT6_434 (
   .O(gates[727]),
   .I0(InputBits[240]),
   .I1(InputBits[1482]),
   .I2(InputBits[673]),
   .I3(InputBits[515]),
   .I4(InputBits[1245]),
   .I5(InputBits[618])
);
LUT6 #(
   .INIT(64'b1001101011111100011001100001001110101111010010111000011011101000)  
) LUT6_435 (
   .O(gates[939]),
   .I0(InputBits[213]),
   .I1(InputBits[1194]),
   .I2(InputBits[968]),
   .I3(InputBits[1718]),
   .I4(InputBits[840]),
   .I5(InputBits[810])
);
LUT6 #(
   .INIT(64'b0111011100110001010010110010010100011111000101010110010100001001)  
) LUT6_436 (
   .O(gates[320]),
   .I0(InputBits[134]),
   .I1(InputBits[306]),
   .I2(InputBits[752]),
   .I3(InputBits[434]),
   .I4(InputBits[1270]),
   .I5(InputBits[1151])
);
LUT6 #(
   .INIT(64'b0110100011010001000100001111110101011111110010110110101110110011)  
) LUT6_437 (
   .O(gates[811]),
   .I0(InputBits[606]),
   .I1(InputBits[1342]),
   .I2(InputBits[605]),
   .I3(InputBits[578]),
   .I4(InputBits[99]),
   .I5(InputBits[895])
);
LUT6 #(
   .INIT(64'b1111000011110111000001101110000101100100000100010000111101101101)  
) LUT6_438 (
   .O(gates[913]),
   .I0(InputBits[1713]),
   .I1(InputBits[1461]),
   .I2(InputBits[315]),
   .I3(InputBits[994]),
   .I4(InputBits[681]),
   .I5(InputBits[1674])
);
LUT6 #(
   .INIT(64'b1001010010110001001110001000001010011010000110100001111011010010)  
) LUT6_439 (
   .O(gates[202]),
   .I0(InputBits[1291]),
   .I1(InputBits[911]),
   .I2(InputBits[1591]),
   .I3(InputBits[1300]),
   .I4(InputBits[1188]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0101000011110001000010111001110101110011110110001001111111010110)  
) LUT6_440 (
   .O(gates[249]),
   .I0(InputBits[1721]),
   .I1(InputBits[1453]),
   .I2(InputBits[465]),
   .I3(InputBits[590]),
   .I4(InputBits[1020]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0100100000001111100001010110100010000111000100011000011111000011)  
) LUT6_441 (
   .O(gates[465]),
   .I0(InputBits[649]),
   .I1(InputBits[1067]),
   .I2(InputBits[1469]),
   .I3(InputBits[1244]),
   .I4(InputBits[237]),
   .I5(InputBits[1335])
);
LUT6 #(
   .INIT(64'b0101011010110110110010110010011011101001000110111010100100100010)  
) LUT6_442 (
   .O(gates[361]),
   .I0(InputBits[217]),
   .I1(InputBits[769]),
   .I2(InputBits[662]),
   .I3(InputBits[778]),
   .I4(InputBits[1119]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1001001110100100010100000110000100001101000111110100000011101011)  
) LUT6_443 (
   .O(gates[184]),
   .I0(InputBits[1601]),
   .I1(InputBits[1173]),
   .I2(InputBits[497]),
   .I3(InputBits[321]),
   .I4(InputBits[1313]),
   .I5(InputBits[1412])
);
LUT6 #(
   .INIT(64'b0101011011110111110110001011111001100010001111111011100011001111)  
) LUT6_444 (
   .O(gates[819]),
   .I0(InputBits[204]),
   .I1(InputBits[562]),
   .I2(InputBits[419]),
   .I3(InputBits[477]),
   .I4(InputBits[379]),
   .I5(InputBits[981])
);
LUT6 #(
   .INIT(64'b1101111111100000110011001000100001110001110111100101111100000110)  
) LUT6_445 (
   .O(gates[1177]),
   .I0(InputBits[948]),
   .I1(InputBits[646]),
   .I2(InputBits[361]),
   .I3(InputBits[928]),
   .I4(InputBits[1471]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b1010010010000100110010010000010001000110101110010110010110110110)  
) LUT6_446 (
   .O(gates[1189]),
   .I0(InputBits[1252]),
   .I1(InputBits[748]),
   .I2(InputBits[1514]),
   .I3(InputBits[137]),
   .I4(InputBits[1125]),
   .I5(InputBits[704])
);
LUT6 #(
   .INIT(64'b1001100101000110010001000001011110110000101101101011110111000010)  
) LUT6_447 (
   .O(gates[776]),
   .I0(InputBits[1122]),
   .I1(InputBits[1402]),
   .I2(InputBits[290]),
   .I3(InputBits[123]),
   .I4(InputBits[1509]),
   .I5(InputBits[657])
);
LUT6 #(
   .INIT(64'b1000000001000111111001101100110100011010001101000100111110110010)  
) LUT6_448 (
   .O(gates[1127]),
   .I0(InputBits[331]),
   .I1(InputBits[1528]),
   .I2(InputBits[266]),
   .I3(InputBits[417]),
   .I4(InputBits[437]),
   .I5(InputBits[1518])
);
LUT6 #(
   .INIT(64'b1011000010011011010101100100000001010101000010000111001101100111)  
) LUT6_449 (
   .O(gates[1537]),
   .I0(InputBits[923]),
   .I1(InputBits[287]),
   .I2(InputBits[785]),
   .I3(InputBits[588]),
   .I4(InputBits[710]),
   .I5(InputBits[822])
);
LUT6 #(
   .INIT(64'b1110110011100001111111110001011101010010101010011001100011000001)  
) LUT6_450 (
   .O(gates[894]),
   .I0(InputBits[894]),
   .I1(InputBits[90]),
   .I2(InputBits[574]),
   .I3(InputBits[945]),
   .I4(InputBits[1607]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b1001101110001010101111001000110010110011001100100101011011001111)  
) LUT6_451 (
   .O(gates[858]),
   .I0(InputBits[1665]),
   .I1(InputBits[1283]),
   .I2(InputBits[200]),
   .I3(InputBits[1256]),
   .I4(InputBits[299]),
   .I5(InputBits[1371])
);
LUT6 #(
   .INIT(64'b0110110101110111111101010110101011000111011111001111111111001011)  
) LUT6_452 (
   .O(gates[1298]),
   .I0(InputBits[1124]),
   .I1(InputBits[1344]),
   .I2(InputBits[1386]),
   .I3(InputBits[1490]),
   .I4(InputBits[627]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b0010100110101000010111001111010111011010110100000110011110001010)  
) LUT6_453 (
   .O(gates[140]),
   .I0(InputBits[84]),
   .I1(InputBits[636]),
   .I2(InputBits[1062]),
   .I3(InputBits[1376]),
   .I4(InputBits[339]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b0011111111101111101111101110011011101101001101000001000001110001)  
) LUT6_454 (
   .O(gates[1459]),
   .I0(InputBits[1583]),
   .I1(InputBits[1581]),
   .I2(InputBits[1328]),
   .I3(InputBits[634]),
   .I4(InputBits[732]),
   .I5(InputBits[985])
);
LUT6 #(
   .INIT(64'b1100000101110100100110010000000111111011110010101111000101110011)  
) LUT6_455 (
   .O(gates[1269]),
   .I0(InputBits[705]),
   .I1(InputBits[1553]),
   .I2(InputBits[729]),
   .I3(InputBits[1440]),
   .I4(InputBits[157]),
   .I5(InputBits[789])
);
LUT6 #(
   .INIT(64'b0010011001001110001100001111011110101100011110100000101011111101)  
) LUT6_456 (
   .O(gates[181]),
   .I0(InputBits[1198]),
   .I1(InputBits[997]),
   .I2(InputBits[966]),
   .I3(InputBits[73]),
   .I4(InputBits[906]),
   .I5(InputBits[1631])
);
LUT6 #(
   .INIT(64'b0001000111100001100010010010101111100100110100110100010011101100)  
) LUT6_457 (
   .O(gates[412]),
   .I0(InputBits[1664]),
   .I1(InputBits[880]),
   .I2(InputBits[1029]),
   .I3(InputBits[408]),
   .I4(InputBits[1167]),
   .I5(InputBits[816])
);
LUT6 #(
   .INIT(64'b1001001000111000001000011011010111011011101101011010011000011010)  
) LUT6_458 (
   .O(gates[954]),
   .I0(InputBits[179]),
   .I1(InputBits[964]),
   .I2(InputBits[530]),
   .I3(InputBits[1368]),
   .I4(InputBits[1055]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0111001011001111000111000100010100111010000110011100101000100111)  
) LUT6_459 (
   .O(gates[385]),
   .I0(InputBits[1675]),
   .I1(InputBits[1395]),
   .I2(InputBits[558]),
   .I3(InputBits[1560]),
   .I4(InputBits[1657]),
   .I5(InputBits[598])
);
LUT6 #(
   .INIT(64'b0010001000111011101001001101010101100010101101101000100011010101)  
) LUT6_460 (
   .O(gates[1479]),
   .I0(InputBits[1651]),
   .I1(InputBits[1419]),
   .I2(InputBits[524]),
   .I3(InputBits[850]),
   .I4(InputBits[1013]),
   .I5(InputBits[871])
);
LUT6 #(
   .INIT(64'b1110111100011100011011011000000011000000011011111010010110101110)  
) LUT6_461 (
   .O(gates[1359]),
   .I0(InputBits[677]),
   .I1(InputBits[831]),
   .I2(InputBits[758]),
   .I3(InputBits[1286]),
   .I4(InputBits[1570]),
   .I5(InputBits[877])
);
LUT6 #(
   .INIT(64'b0101010110011010000000001001100000000100101111011110010111101111)  
) LUT6_462 (
   .O(gates[307]),
   .I0(InputBits[687]),
   .I1(InputBits[1274]),
   .I2(InputBits[887]),
   .I3(InputBits[699]),
   .I4(InputBits[432]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0101100110011101011100100001001010100110010100010111000100110011)  
) LUT6_463 (
   .O(gates[801]),
   .I0(InputBits[1432]),
   .I1(InputBits[13]),
   .I2(InputBits[1026]),
   .I3(InputBits[252]),
   .I4(InputBits[144]),
   .I5(InputBits[1347])
);
LUT6 #(
   .INIT(64'b1011100010110000111011100010001011100010000101000011011001000111)  
) LUT6_464 (
   .O(gates[985]),
   .I0(InputBits[459]),
   .I1(InputBits[1047]),
   .I2(InputBits[922]),
   .I3(InputBits[265]),
   .I4(InputBits[1538]),
   .I5(InputBits[953])
);
LUT6 #(
   .INIT(64'b1000000011101110111110100110001101111001000010101101001001010010)  
) LUT6_465 (
   .O(gates[1463]),
   .I0(InputBits[741]),
   .I1(InputBits[736]),
   .I2(InputBits[632]),
   .I3(InputBits[376]),
   .I4(InputBits[1036]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1110100001001100010111001001100010101101101000001001001011010101)  
) LUT6_466 (
   .O(gates[154]),
   .I0(InputBits[555]),
   .I1(InputBits[1289]),
   .I2(InputBits[902]),
   .I3(InputBits[247]),
   .I4(InputBits[413]),
   .I5(InputBits[1220])
);
LUT6 #(
   .INIT(64'b0010000010100011000000110010110000001111110111001011110101010010)  
) LUT6_467 (
   .O(gates[830]),
   .I0(InputBits[1476]),
   .I1(InputBits[1456]),
   .I2(InputBits[689]),
   .I3(InputBits[1308]),
   .I4(InputBits[1593]),
   .I5(InputBits[1113])
);
LUT6 #(
   .INIT(64'b0100011101010001110101111111010111110010001000010010111010001110)  
) LUT6_468 (
   .O(gates[971]),
   .I0(InputBits[1543]),
   .I1(InputBits[1604]),
   .I2(InputBits[1695]),
   .I3(InputBits[718]),
   .I4(InputBits[856]),
   .I5(InputBits[1557])
);
LUT6 #(
   .INIT(64'b1011100010100001110111001100011100011011011101010001000001111010)  
) LUT6_469 (
   .O(gates[1467]),
   .I0(InputBits[1614]),
   .I1(InputBits[145]),
   .I2(InputBits[1293]),
   .I3(InputBits[676]),
   .I4(InputBits[1054]),
   .I5(InputBits[406])
);
LUT6 #(
   .INIT(64'b0100011110101010000111100000001101100001000110001000001100111010)  
) LUT6_470 (
   .O(gates[754]),
   .I0(InputBits[1540]),
   .I1(InputBits[1676]),
   .I2(InputBits[488]),
   .I3(InputBits[1706]),
   .I4(InputBits[576]),
   .I5(InputBits[1132])
);
LUT6 #(
   .INIT(64'b1001101101111101011100101001101001001111001001000001010111000000)  
) LUT6_471 (
   .O(gates[479]),
   .I0(InputBits[783]),
   .I1(InputBits[457]),
   .I2(InputBits[66]),
   .I3(InputBits[1415]),
   .I4(InputBits[347]),
   .I5(InputBits[776])
);
LUT6 #(
   .INIT(64'b0111100000010011100000000011100001010110000000011000010111110010)  
) LUT6_472 (
   .O(gates[847]),
   .I0(InputBits[6]),
   .I1(InputBits[1646]),
   .I2(InputBits[1702]),
   .I3(InputBits[311]),
   .I4(InputBits[329]),
   .I5(InputBits[565])
);
LUT6 #(
   .INIT(64'b0000001000000000101010111000010010001001011100001011100010010111)  
) LUT6_473 (
   .O(gates[1101]),
   .I0(InputBits[446]),
   .I1(InputBits[1661]),
   .I2(InputBits[560]),
   .I3(InputBits[303]),
   .I4(InputBits[763]),
   .I5(InputBits[592])
);
LUT6 #(
   .INIT(64'b1011111010100000010001000111001101100110000000101101110011111010)  
) LUT6_474 (
   .O(gates[1166]),
   .I0(InputBits[26]),
   .I1(InputBits[1096]),
   .I2(InputBits[49]),
   .I3(InputBits[1171]),
   .I4(InputBits[1480]),
   .I5(InputBits[1209])
);
LUT6 #(
   .INIT(64'b1101111110000100110000110100010100001000110100011001010001010100)  
) LUT6_475 (
   .O(gates[704]),
   .I0(InputBits[1242]),
   .I1(InputBits[1]),
   .I2(InputBits[254]),
   .I3(InputBits[480]),
   .I4(InputBits[1189]),
   .I5(InputBits[653])
);
LUT6 #(
   .INIT(64'b1111101111101000001111001000000011101101000101001011100111100010)  
) LUT6_476 (
   .O(gates[326]),
   .I0(InputBits[176]),
   .I1(InputBits[1004]),
   .I2(InputBits[1644]),
   .I3(InputBits[211]),
   .I4(InputBits[191]),
   .I5(InputBits[1060])
);
LUT6 #(
   .INIT(64'b1110100011001101001110001101011110000100001011111000001001110010)  
) LUT6_477 (
   .O(gates[1378]),
   .I0(InputBits[612]),
   .I1(InputBits[425]),
   .I2(InputBits[581]),
   .I3(InputBits[720]),
   .I4(InputBits[1130]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1010000101101101111100000110011000110001010110101111011010010100)  
) LUT6_478 (
   .O(gates[1003]),
   .I0(InputBits[1598]),
   .I1(InputBits[1579]),
   .I2(InputBits[1530]),
   .I3(InputBits[1473]),
   .I4(InputBits[1616]),
   .I5(InputBits[1277])
);
LUT6 #(
   .INIT(64'b1101100000011010000001110101101010011001111010010011100110011001)  
) LUT6_479 (
   .O(gates[1462]),
   .I0(InputBits[517]),
   .I1(InputBits[1726]),
   .I2(InputBits[1694]),
   .I3(InputBits[1566]),
   .I4(InputBits[647]),
   .I5(InputBits[1716])
);
LUT6 #(
   .INIT(64'b0010010111101001111000000100001001101100101100111101110010111000)  
) LUT6_480 (
   .O(gates[1165]),
   .I0(InputBits[683]),
   .I1(InputBits[313]),
   .I2(InputBits[1599]),
   .I3(InputBits[1069]),
   .I4(InputBits[208]),
   .I5(InputBits[1410])
);
LUT6 #(
   .INIT(64'b1001010010111010010000000101101100000001110010010111111011100100)  
) LUT6_481 (
   .O(gates[1054]),
   .I0(InputBits[355]),
   .I1(InputBits[235]),
   .I2(InputBits[323]),
   .I3(InputBits[1207]),
   .I4(InputBits[1521]),
   .I5(InputBits[833])
);
LUT6 #(
   .INIT(64'b0011111000001000000001001111111010011110010001001111010010110010)  
) LUT6_482 (
   .O(gates[681]),
   .I0(InputBits[1383]),
   .I1(InputBits[709]),
   .I2(InputBits[135]),
   .I3(InputBits[1409]),
   .I4(InputBits[1709]),
   .I5(InputBits[1156])
);
LUT6 #(
   .INIT(64'b1100010110010100100100101100000010001011100011110111110000010110)  
) LUT6_483 (
   .O(gates[619]),
   .I0(InputBits[545]),
   .I1(InputBits[427]),
   .I2(InputBits[947]),
   .I3(InputBits[1363]),
   .I4(InputBits[838]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1100100111001101110101001011111000011110011001010111000001101101)  
) LUT6_484 (
   .O(gates[335]),
   .I0(InputBits[1248]),
   .I1(InputBits[1320]),
   .I2(InputBits[1667]),
   .I3(InputBits[1450]),
   .I4(InputBits[285]),
   .I5(InputBits[853])
);
LUT6 #(
   .INIT(64'b1101101101100111000100010010110111000001100011110000001010101011)  
) LUT6_485 (
   .O(gates[1029]),
   .I0(InputBits[514]),
   .I1(InputBits[1590]),
   .I2(InputBits[268]),
   .I3(InputBits[500]),
   .I4(InputBits[712]),
   .I5(InputBits[982])
);
LUT6 #(
   .INIT(64'b0011111100111100000011010100101100010101001011100000000001001001)  
) LUT6_486 (
   .O(gates[5]),
   .I0(InputBits[1396]),
   .I1(InputBits[1255]),
   .I2(InputBits[1649]),
   .I3(InputBits[473]),
   .I4(InputBits[106]),
   .I5(InputBits[1520])
);
LUT6 #(
   .INIT(64'b1111011001000111001010010111000101011011101011111110111010011100)  
) LUT6_487 (
   .O(gates[698]),
   .I0(InputBits[750]),
   .I1(InputBits[1486]),
   .I2(InputBits[51]),
   .I3(InputBits[509]),
   .I4(InputBits[37]),
   .I5(InputBits[378])
);
LUT6 #(
   .INIT(64'b0000101101000001010101000101100110101001000001111000011011001101)  
) LUT6_488 (
   .O(gates[621]),
   .I0(InputBits[202]),
   .I1(InputBits[467]),
   .I2(InputBits[127]),
   .I3(InputBits[525]),
   .I4(InputBits[1226]),
   .I5(InputBits[1442])
);
LUT6 #(
   .INIT(64'b0100010101101010101101001101000110010101111100011000010101011110)  
) LUT6_489 (
   .O(gates[524]),
   .I0(InputBits[861]),
   .I1(InputBits[552]),
   .I2(InputBits[142]),
   .I3(InputBits[43]),
   .I4(InputBits[656]),
   .I5(InputBits[727])
);
LUT6 #(
   .INIT(64'b1111100110000001110101110101111000110001110000110111011010101011)  
) LUT6_490 (
   .O(gates[554]),
   .I0(InputBits[215]),
   .I1(InputBits[1205]),
   .I2(InputBits[301]),
   .I3(InputBits[974]),
   .I4(InputBits[1180]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b1011001001111001000101010010001011101110110001000000110011000001)  
) LUT6_491 (
   .O(gates[552]),
   .I0(InputBits[760]),
   .I1(InputBits[802]),
   .I2(InputBits[929]),
   .I3(InputBits[702]),
   .I4(InputBits[889]),
   .I5(InputBits[1104])
);
LUT6 #(
   .INIT(64'b0011011011111010111000010001110110011010010001000011010010001100)  
) LUT6_492 (
   .O(gates[598]),
   .I0(InputBits[1430]),
   .I1(InputBits[793]),
   .I2(InputBits[691]),
   .I3(InputBits[1090]),
   .I4(InputBits[439]),
   .I5(InputBits[1697])
);
LUT6 #(
   .INIT(64'b0110001011011100111111100111000000110010000100000000010011111011)  
) LUT6_493 (
   .O(gates[780]),
   .I0(InputBits[1078]),
   .I1(InputBits[1655]),
   .I2(InputBits[71]),
   .I3(InputBits[1618]),
   .I4(InputBits[664]),
   .I5(InputBits[586])
);
LUT6 #(
   .INIT(64'b0100100001000000110011100110110110001101010111000101111111101100)  
) LUT6_494 (
   .O(gates[1433]),
   .I0(InputBits[904]),
   .I1(InputBits[909]),
   .I2(InputBits[642]),
   .I3(InputBits[161]),
   .I4(InputBits[1299]),
   .I5(InputBits[226])
);
LUT6 #(
   .INIT(64'b1001110100110110110110100100000110000111001111101000001010011001)  
) LUT6_495 (
   .O(gates[74]),
   .I0(InputBits[108]),
   .I1(InputBits[1333]),
   .I2(InputBits[128]),
   .I3(InputBits[602]),
   .I4(InputBits[56]),
   .I5(InputBits[858])
);
LUT6 #(
   .INIT(64'b0011010000010010111011001101010110100100101100111000101010011100)  
) LUT6_496 (
   .O(gates[240]),
   .I0(InputBits[1011]),
   .I1(InputBits[1491]),
   .I2(InputBits[280]),
   .I3(InputBits[11]),
   .I4(InputBits[829]),
   .I5(InputBits[1326])
);
LUT6 #(
   .INIT(64'b1101011100010101001001010110111001000101101010011101101111110100)  
) LUT6_497 (
   .O(gates[890]),
   .I0(InputBits[260]),
   .I1(InputBits[1082]),
   .I2(InputBits[534]),
   .I3(InputBits[532]),
   .I4(InputBits[1546]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0001000011111000111000101011100000010000011011011000110101001011)  
) LUT6_498 (
   .O(gates[440]),
   .I0(InputBits[629]),
   .I1(InputBits[743]),
   .I2(InputBits[1606]),
   .I3(InputBits[1463]),
   .I4(InputBits[808]),
   .I5(InputBits[781])
);
LUT6 #(
   .INIT(64'b1101110110001011101101000010011001100100010100110010110111100000)  
) LUT6_499 (
   .O(gates[230]),
   .I0(InputBits[1353]),
   .I1(InputBits[738]),
   .I2(InputBits[152]),
   .I3(InputBits[956]),
   .I4(InputBits[1548]),
   .I5(InputBits[1049])
);
LUT6 #(
   .INIT(64'b0100101011110101101001011110010101111001001010111001000101111010)  
) LUT6_500 (
   .O(gates[115]),
   .I0(InputBits[1533]),
   .I1(InputBits[337]),
   .I2(InputBits[635]),
   .I3(InputBits[222]),
   .I4(InputBits[489]),
   .I5(InputBits[991])
);
LUT6 #(
   .INIT(64'b0101011111111001011111100100001000110000010110110101011000001110)  
) LUT6_501 (
   .O(gates[1289]),
   .I0(InputBits[1258]),
   .I1(InputBits[939]),
   .I2(InputBits[1169]),
   .I3(InputBits[962]),
   .I4(InputBits[1022]),
   .I5(InputBits[1111])
);
LUT6 #(
   .INIT(64'b1100101010001001001101100110010000110010101011110111011001110111)  
) LUT6_502 (
   .O(gates[299]),
   .I0(InputBits[1457]),
   .I1(InputBits[774]),
   .I2(InputBits[1179]),
   .I3(InputBits[410]),
   .I4(InputBits[45]),
   .I5(InputBits[1685])
);
LUT6 #(
   .INIT(64'b0010100110100000011111100011100000110010001101101111100111011111)  
) LUT6_503 (
   .O(gates[377]),
   .I0(InputBits[185]),
   .I1(InputBits[1425]),
   .I2(InputBits[1098]),
   .I3(InputBits[1195]),
   .I4(InputBits[1101]),
   .I5(InputBits[972])
);
LUT6 #(
   .INIT(64'b0101110000100010101000110100001101011111011010010001110010110001)  
) LUT6_504 (
   .O(gates[1282]),
   .I0(InputBits[993]),
   .I1(InputBits[527]),
   .I2(InputBits[295]),
   .I3(InputBits[1501]),
   .I4(InputBits[1058]),
   .I5(InputBits[1138])
);
LUT6 #(
   .INIT(64'b1101001101010000010110111110110111001101011100100101010010000010)  
) LUT6_505 (
   .O(gates[922]),
   .I0(InputBits[409]),
   .I1(InputBits[1547]),
   .I2(InputBits[1692]),
   .I3(InputBits[1070]),
   .I4(InputBits[1158]),
   .I5(InputBits[1263])
);
LUT6 #(
   .INIT(64'b1001101111000011111101001110100110001011010000010011011011101101)  
) LUT6_506 (
   .O(gates[602]),
   .I0(InputBits[869]),
   .I1(InputBits[916]),
   .I2(InputBits[64]),
   .I3(InputBits[1711]),
   .I4(InputBits[551]),
   .I5(InputBits[1141])
);
LUT6 #(
   .INIT(64'b0001010010001110111011111000101000001011001001111100111010001110)  
) LUT6_507 (
   .O(gates[841]),
   .I0(InputBits[1325]),
   .I1(InputBits[756]),
   .I2(InputBits[1523]),
   .I3(InputBits[643]),
   .I4(InputBits[138]),
   .I5(InputBits[1001])
);
LUT6 #(
   .INIT(64'b0110011111101100101110001100001010111101111000010010000111000100)  
) LUT6_508 (
   .O(gates[1311]),
   .I0(InputBits[1392]),
   .I1(InputBits[251]),
   .I2(InputBits[733]),
   .I3(InputBits[183]),
   .I4(InputBits[231]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b1100111101011111011110011000011101000000001100000001010011110010)  
) LUT6_509 (
   .O(gates[1044]),
   .I0(InputBits[294]),
   .I1(InputBits[1399]),
   .I2(InputBits[765]),
   .I3(InputBits[1094]),
   .I4(InputBits[1185]),
   .I5(InputBits[885])
);
LUT6 #(
   .INIT(64'b1011010100000100000101100111001101100000001000101111100011010000)  
) LUT6_510 (
   .O(gates[1072]),
   .I0(InputBits[585]),
   .I1(InputBits[1233]),
   .I2(InputBits[716]),
   .I3(InputBits[1670]),
   .I4(InputBits[812]),
   .I5(InputBits[1218])
);
LUT6 #(
   .INIT(64'b1000100011011001111000011100111001001011101010111011111000110000)  
) LUT6_511 (
   .O(gates[1394]),
   .I0(InputBits[1500]),
   .I1(InputBits[1704]),
   .I2(InputBits[445]),
   .I3(InputBits[882]),
   .I4(InputBits[976]),
   .I5(InputBits[890])
);
LUT6 #(
   .INIT(64'b0001101000110011000010011010100011110111100111000101010000110110)  
) LUT6_512 (
   .O(gates[612]),
   .I0(InputBits[1576]),
   .I1(InputBits[1134]),
   .I2(InputBits[1485]),
   .I3(InputBits[874]),
   .I4(InputBits[1516]),
   .I5(InputBits[1235])
);
LUT6 #(
   .INIT(64'b0100001001011010011011110101101001011000110010100100010000000111)  
) LUT6_513 (
   .O(gates[1350]),
   .I0(InputBits[1717]),
   .I1(InputBits[384]),
   .I2(InputBits[855]),
   .I3(InputBits[424]),
   .I4(InputBits[1542]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b1111011010111010000110010010011101100101110010001101111101001101)  
) LUT6_514 (
   .O(gates[936]),
   .I0(InputBits[1511]),
   .I1(InputBits[374]),
   .I2(InputBits[930]),
   .I3(InputBits[182]),
   .I4(InputBits[393]),
   .I5(InputBits[1588])
);
LUT6 #(
   .INIT(64'b1110101001110110011111000110110010100001010010001110111001101101)  
) LUT6_515 (
   .O(gates[1391]),
   .I0(InputBits[403]),
   .I1(InputBits[407]),
   .I2(InputBits[1578]),
   .I3(InputBits[1006]),
   .I4(InputBits[54]),
   .I5(InputBits[415])
);
LUT6 #(
   .INIT(64'b0010111100111000000011011110110101001001011010101000101111100101)  
) LUT6_516 (
   .O(gates[1277]),
   .I0(InputBits[836]),
   .I1(InputBits[225]),
   .I2(InputBits[1668]),
   .I3(InputBits[1689]),
   .I4(InputBits[567]),
   .I5(InputBits[1264])
);
LUT6 #(
   .INIT(64'b0001101110101001110010101001101000101010101100110011000000010111)  
) LUT6_517 (
   .O(gates[91]),
   .I0(InputBits[309]),
   .I1(InputBits[725]),
   .I2(InputBits[1659]),
   .I3(InputBits[48]),
   .I4(InputBits[875]),
   .I5(InputBits[678])
);
LUT6 #(
   .INIT(64'b1101010011111111100011100001110000011010111010111101010111011100)  
) LUT6_518 (
   .O(gates[1086]),
   .I0(InputBits[1388]),
   .I1(InputBits[326]),
   .I2(InputBits[1041]),
   .I3(InputBits[826]),
   .I4(InputBits[707]),
   .I5(InputBits[1216])
);
LUT6 #(
   .INIT(64'b1111111010100100111000100101010010111000100100011000010011100101)  
) LUT6_519 (
   .O(gates[1240]),
   .I0(InputBits[820]),
   .I1(InputBits[381]),
   .I2(InputBits[701]),
   .I3(InputBits[1204]),
   .I4(InputBits[494]),
   .I5(InputBits[103])
);
LUT6 #(
   .INIT(64'b1111010011001111010011101011100000110010100011000110110011100000)  
) LUT6_520 (
   .O(gates[467]),
   .I0(InputBits[1357]),
   .I1(InputBits[1642]),
   .I2(InputBits[88]),
   .I3(InputBits[957]),
   .I4(InputBits[10]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0100110111001110010010000010000110001011110100000001111000110001)  
) LUT6_521 (
   .O(gates[701]),
   .I0(InputBits[502]),
   .I1(InputBits[241]),
   .I2(InputBits[80]),
   .I3(InputBits[806]),
   .I4(InputBits[1443]),
   .I5(InputBits[620])
);
LUT6 #(
   .INIT(64'b0010010000111100100011101110011100000001100000100101111101001001)  
) LUT6_522 (
   .O(gates[474]),
   .I0(InputBits[1083]),
   .I1(InputBits[317]),
   .I2(InputBits[935]),
   .I3(InputBits[1008]),
   .I4(InputBits[503]),
   .I5(InputBits[1531])
);
LUT6 #(
   .INIT(64'b1010001000111101010111100110001111111101000010110011101100011100)  
) LUT6_523 (
   .O(gates[481]),
   .I0(InputBits[78]),
   .I1(InputBits[1088]),
   .I2(InputBits[1322]),
   .I3(InputBits[1380]),
   .I4(InputBits[387]),
   .I5(InputBits[958])
);
LUT6 #(
   .INIT(64'b0100100000000101100111101001010000111111001010001101111000101111)  
) LUT6_524 (
   .O(gates[867]),
   .I0(InputBits[487]),
   .I1(InputBits[450]),
   .I2(InputBits[151]),
   .I3(InputBits[284]),
   .I4(InputBits[1273]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1000000010001100000101000110001010001101011011011010001000100100)  
) LUT6_525 (
   .O(gates[214]),
   .I0(InputBits[631]),
   .I1(InputBits[1285]),
   .I2(InputBits[47]),
   .I3(InputBits[452]),
   .I4(InputBits[405]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b0011101011010110011111111101001010011100011011011000110110000111)  
) LUT6_526 (
   .O(gates[564]),
   .I0(InputBits[800]),
   .I1(InputBits[1228]),
   .I2(InputBits[357]),
   .I3(InputBits[609]),
   .I4(InputBits[737]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b1000010111011111101010100111100110001010111000110011010001011100)  
) LUT6_527 (
   .O(gates[817]),
   .I0(InputBits[1467]),
   .I1(InputBits[125]),
   .I2(InputBits[398]),
   .I3(InputBits[1324]),
   .I4(InputBits[1202]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0100000000000001110011101111101111001000111101010111010101111000)  
) LUT6_528 (
   .O(gates[563]),
   .I0(InputBits[899]),
   .I1(InputBits[522]),
   .I2(InputBits[481]),
   .I3(InputBits[484]),
   .I4(InputBits[192]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1010101101001110101100011110111001011000101010101011110011011110)  
) LUT6_529 (
   .O(gates[731]),
   .I0(InputBits[1573]),
   .I1(InputBits[1030]),
   .I2(InputBits[69]),
   .I3(InputBits[244]),
   .I4(InputBits[1337]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0011000111100100011101000111000110110011101001011001001101001111)  
) LUT6_530 (
   .O(gates[657]),
   .I0(InputBits[140]),
   .I1(InputBits[979]),
   .I2(InputBits[823]),
   .I3(InputBits[1428]),
   .I4(InputBits[149]),
   .I5(InputBits[1459])
);
LUT6 #(
   .INIT(64'b1100001010110101000110010101000010111110101011101100011011001000)  
) LUT6_531 (
   .O(gates[229]),
   .I0(InputBits[1529]),
   .I1(InputBits[1332]),
   .I2(InputBits[194]),
   .I3(InputBits[897]),
   .I4(InputBits[573]),
   .I5(InputBits[668])
);
LUT6 #(
   .INIT(64'b1010001001110011000000111011011010101000010100000101111000011010)  
) LUT6_532 (
   .O(gates[768]),
   .I0(InputBits[1146]),
   .I1(InputBits[1129]),
   .I2(InputBits[1597]),
   .I3(InputBits[1015]),
   .I4(InputBits[385]),
   .I5(InputBits[754])
);
LUT6 #(
   .INIT(64'b1111110110101010011011101001011110000000000001111001001001001001)  
) LUT6_533 (
   .O(gates[1092]),
   .I0(InputBits[86]),
   .I1(InputBits[360]),
   .I2(InputBits[1407]),
   .I3(InputBits[1109]),
   .I4(InputBits[1182]),
   .I5(InputBits[1629])
);
LUT6 #(
   .INIT(64'b1000001110010111000011100100010100001111010000010001011110100111)  
) LUT6_534 (
   .O(gates[673]),
   .I0(InputBits[513]),
   .I1(InputBits[171]),
   .I2(InputBits[1003]),
   .I3(InputBits[1348]),
   .I4(InputBits[1117]),
   .I5(InputBits[610])
);
LUT6 #(
   .INIT(64'b0101111011001010010001110011001100011010001110111010011011010011)  
) LUT6_535 (
   .O(gates[503]),
   .I0(InputBits[263]),
   .I1(InputBits[792]),
   .I2(InputBits[539]),
   .I3(InputBits[282]),
   .I4(InputBits[159]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b1011010011110000010110110110110100100001110101011110000011011001)  
) LUT6_536 (
   .O(gates[68]),
   .I0(InputBits[351]),
   .I1(InputBits[1231]),
   .I2(InputBits[1535]),
   .I3(InputBits[117]),
   .I4(InputBits[1422]),
   .I5(InputBits[1680])
);
LUT6 #(
   .INIT(64'b1110000101101101001000011010000111001111011100001110101111100101)  
) LUT6_537 (
   .O(gates[1483]),
   .I0(InputBits[768]),
   .I1(InputBits[770]),
   .I2(InputBits[130]),
   .I3(InputBits[456]),
   .I4(InputBits[336]),
   .I5(InputBits[1494])
);
LUT6 #(
   .INIT(64'b1110001111000110001101101000111001001011001101000011101101000110)  
) LUT6_538 (
   .O(gates[315]),
   .I0(InputBits[1267]),
   .I1(InputBits[1213]),
   .I2(InputBits[713]),
   .I3(InputBits[1478]),
   .I4(InputBits[772]),
   .I5(InputBits[714])
);
LUT6 #(
   .INIT(64'b0010010100010101011011011010100101101100111110101101100100110010)  
) LUT6_539 (
   .O(gates[338]),
   .I0(InputBits[1624]),
   .I1(InputBits[1634]),
   .I2(InputBits[1359]),
   .I3(InputBits[989]),
   .I4(InputBits[1351]),
   .I5(InputBits[986])
);
LUT6 #(
   .INIT(64'b1010001010010100000001100011100100101010110001001110010100001001)  
) LUT6_540 (
   .O(gates[1347]),
   .I0(InputBits[1666]),
   .I1(InputBits[1177]),
   .I2(InputBits[1297]),
   .I3(InputBits[600]),
   .I4(InputBits[38]),
   .I5(InputBits[844])
);
LUT6 #(
   .INIT(64'b1100011110010010010000001010100101110000010111010011010001100100)  
) LUT6_541 (
   .O(gates[576]),
   .I0(InputBits[156]),
   .I1(InputBits[1436]),
   .I2(InputBits[1052]),
   .I3(InputBits[1281]),
   .I4(InputBits[547]),
   .I5(InputBits[1024])
);
LUT6 #(
   .INIT(64'b1111110111000001011001101001000010100010010001110101001011101000)  
) LUT6_542 (
   .O(gates[761]),
   .I0(InputBits[1687]),
   .I1(InputBits[461]),
   .I2(InputBits[1627]),
   .I3(InputBits[1513]),
   .I4(InputBits[165]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b1001010011001111000100010000000111001010010101100011110111101001)  
) LUT6_543 (
   .O(gates[222]),
   .I0(InputBits[1498]),
   .I1(InputBits[651]),
   .I2(InputBits[622]),
   .I3(InputBits[333]),
   .I4(InputBits[941]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0110011111110100100100000010010011011000101111011001001000001110)  
) LUT6_544 (
   .O(gates[1504]),
   .I0(InputBits[1712]),
   .I1(InputBits[731]),
   .I2(InputBits[814]),
   .I3(InputBits[375]),
   .I4(InputBits[1092]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b1000111010011101001000100110000001010010001010000000000110000110)  
) LUT6_545 (
   .O(gates[25]),
   .I0(InputBits[1261]),
   .I1(InputBits[195]),
   .I2(InputBits[253]),
   .I3(InputBits[184]),
   .I4(InputBits[1247]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b0101101110110001100011010000100010110001001000111110011100101010)  
) LUT6_546 (
   .O(gates[738]),
   .I0(InputBits[496]),
   .I1(InputBits[1127]),
   .I2(InputBits[1268]),
   .I3(InputBits[1446]),
   .I4(InputBits[934]),
   .I5(InputBits[849])
);
LUT6 #(
   .INIT(64'b0101010001110111011111111001101010100100001100010001110110110110)  
) LUT6_547 (
   .O(gates[1415]),
   .I0(InputBits[1100]),
   .I1(InputBits[1622]),
   .I2(InputBits[954]),
   .I3(InputBits[1148]),
   .I4(InputBits[1400]),
   .I5(InputBits[616])
);
LUT6 #(
   .INIT(64'b1110001100000100001100011111100011101110101110010100110001111010)  
) LUT6_548 (
   .O(gates[484]),
   .I0(InputBits[1056]),
   .I1(InputBits[411]),
   .I2(InputBits[454]),
   .I3(InputBits[110]),
   .I4(InputBits[354]),
   .I5(InputBits[1072])
);
LUT6 #(
   .INIT(64'b1011010101111100110101110100001110101011110011000101010011010101)  
) LUT6_549 (
   .O(gates[1036]),
   .I0(InputBits[227]),
   .I1(InputBits[884]),
   .I2(InputBits[1143]),
   .I3(InputBits[697]),
   .I4(InputBits[1187]),
   .I5(InputBits[951])
);
LUT6 #(
   .INIT(64'b0101010011110010101100000011011111110101001101100100000011101110)  
) LUT6_550 (
   .O(gates[1078]),
   .I0(InputBits[529]),
   .I1(InputBits[918]),
   .I2(InputBits[1043]),
   .I3(InputBits[1654]),
   .I4(InputBits[1567]),
   .I5(InputBits[615])
);
LUT6 #(
   .INIT(64'b0100010111011000101000001100110111111100110100010010101100011010)  
) LUT6_551 (
   .O(gates[1243]),
   .I0(InputBits[1341]),
   .I1(InputBits[780]),
   .I2(InputBits[867]),
   .I3(InputBits[1366]),
   .I4(InputBits[435]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1011000111000011111101111011010001001011001101011011110100110001)  
) LUT6_552 (
   .O(gates[305]),
   .I0(InputBits[1699]),
   .I1(InputBits[97]),
   .I2(InputBits[846]),
   .I3(InputBits[1640]),
   .I4(InputBits[937]),
   .I5(InputBits[907])
);
LUT6 #(
   .INIT(64'b0110100101110111000110110110001000100001101000011000001100010010)  
) LUT6_553 (
   .O(gates[1253]),
   .I0(InputBits[498]),
   .I1(InputBits[1378]),
   .I2(InputBits[554]),
   .I3(InputBits[154]),
   .I4(InputBits[746]),
   .I5(InputBits[472])
);
LUT6 #(
   .INIT(64'b0011001111110010100010111010100010000111000100000000110110000011)  
) LUT6_554 (
   .O(gates[928]),
   .I0(InputBits[926]),
   .I1(InputBits[914]),
   .I2(InputBits[1317]),
   .I3(InputBits[190]),
   .I4(InputBits[1039]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b0011000000000000101011101111100001110111011110100001001100011111)  
) LUT6_555 (
   .O(gates[1265]),
   .I0(InputBits[535]),
   .I1(InputBits[307]),
   .I2(InputBits[797]),
   .I3(InputBits[569]),
   .I4(InputBits[342]),
   .I5(InputBits[1105])
);
LUT6 #(
   .INIT(64'b1000001011101101110011010111101110001110100111010011111001011011)  
) LUT6_556 (
   .O(gates[544]),
   .I0(InputBits[297]),
   .I1(InputBits[1136]),
   .I2(InputBits[817]),
   .I3(InputBits[1503]),
   .I4(InputBits[401]),
   .I5(InputBits[1390])
);
LUT6 #(
   .INIT(64'b1000000011110001111100101001010001111011101100101111111001010110)  
) LUT6_557 (
   .O(gates[623]),
   .I0(InputBits[693]),
   .I1(InputBits[1223]),
   .I2(InputBits[680]),
   .I3(InputBits[1620]),
   .I4(InputBits[1526]),
   .I5(InputBits[1254])
);
LUT6 #(
   .INIT(64'b0111101100000010000101001001001101101001001001010111001110100110)  
) LUT6_558 (
   .O(gates[1512]),
   .I0(InputBits[1544]),
   .I1(InputBits[1723]),
   .I2(InputBits[1076]),
   .I3(InputBits[723]),
   .I4(InputBits[872]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0100000001111101110110001111010111010011101000110101101101110011)  
) LUT6_559 (
   .O(gates[1526]),
   .I0(InputBits[82]),
   .I1(InputBits[1211]),
   .I2(InputBits[1373]),
   .I3(InputBits[239]),
   .I4(InputBits[638]),
   .I5(InputBits[1081])
);
LUT6 #(
   .INIT(64'b0011100111011111101011000111110110111111110101010000001111000100)  
) LUT6_560 (
   .O(gates[1196]),
   .I0(InputBits[537]),
   .I1(InputBits[1413]),
   .I2(InputBits[944]),
   .I3(InputBits[901]),
   .I4(InputBits[1636]),
   .I5(InputBits[1250])
);
LUT6 #(
   .INIT(64'b0101001100010011000100011111101110000101001110011100110101111100)  
) LUT6_561 (
   .O(gates[1114]),
   .I0(InputBits[541]),
   .I1(InputBits[229]),
   .I2(InputBits[1284]),
   .I3(InputBits[124]),
   .I4(InputBits[594]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0001111001110001001101110101101101110010111000111001001001011010)  
) LUT6_562 (
   .O(gates[217]),
   .I0(InputBits[1462]),
   .I1(InputBits[1085]),
   .I2(InputBits[65]),
   .I3(InputBits[1145]),
   .I4(InputBits[686]),
   .I5(InputBits[1549])
);
LUT6 #(
   .INIT(64'b0111001010101011110000010111101111111001111010100001010001011110)  
) LUT6_563 (
   .O(gates[328]),
   .I0(InputBits[1420]),
   .I1(InputBits[1505]),
   .I2(InputBits[1612]),
   .I3(InputBits[1192]),
   .I4(InputBits[328]),
   .I5(InputBits[607])
);
LUT6 #(
   .INIT(64'b1111010111111101000101000101110100110011001100100110110111101000)  
) LUT6_564 (
   .O(gates[239]),
   .I0(InputBits[815]),
   .I1(InputBits[291]),
   .I2(InputBits[660]),
   .I3(InputBits[1116]),
   .I4(InputBits[370]),
   .I5(InputBits[999])
);
LUT6 #(
   .INIT(64'b1000101110011001101100000001010011110111011110011100101011101110)  
) LUT6_565 (
   .O(gates[122]),
   .I0(InputBits[1019]),
   .I1(InputBits[1361]),
   .I2(InputBits[1571]),
   .I3(InputBits[1045]),
   .I4(InputBits[960]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b0111001100001101111111111001100011110101110111101111101111000011)  
) LUT6_566 (
   .O(gates[1223]),
   .I0(InputBits[28]),
   .I1(InputBits[862]),
   .I2(InputBits[76]),
   .I3(InputBits[273]),
   .I4(InputBits[1050]),
   .I5(InputBits[1065])
);
LUT6 #(
   .INIT(64'b0100110100111001000101110001001000100001100001110011010000001100)  
) LUT6_567 (
   .O(gates[878]),
   .I0(InputBits[739]),
   .I1(InputBits[1451]),
   .I2(InputBits[583]),
   .I3(InputBits[965]),
   .I4(InputBits[892]),
   .I5(InputBits[670])
);
LUT6 #(
   .INIT(64'b0001101011000111010011000100000100001111000011101100001110000100)  
) LUT6_568 (
   .O(gates[281]),
   .I0(InputBits[23]),
   .I1(InputBits[1673]),
   .I2(InputBits[1585]),
   .I3(InputBits[1488]),
   .I4(InputBits[1063]),
   .I5(InputBits[1426])
);
LUT6 #(
   .INIT(64'b0000110110001100001010100101001010111110010000010001010001000011)  
) LUT6_569 (
   .O(gates[269]),
   .I0(InputBits[1483]),
   .I1(InputBits[596]),
   .I2(InputBits[1238]),
   .I3(InputBits[274]),
   .I4(InputBits[362]),
   .I5(InputBits[1033])
);
LUT6 #(
   .INIT(64'b0111111010010110101110001001001010011100111001010111101111110001)  
) LUT6_570 (
   .O(gates[628]),
   .I0(InputBits[1438]),
   .I1(InputBits[349]),
   .I2(InputBits[206]),
   .I3(InputBits[74]),
   .I4(InputBits[363]),
   .I5(InputBits[1200])
);
LUT6 #(
   .INIT(64'b0100101011110110010001011101010110100011100100011001111011100000)  
) LUT6_571 (
   .O(gates[158]),
   .I0(InputBits[641]),
   .I1(InputBits[147]),
   .I2(InputBits[1682]),
   .I3(InputBits[1563]),
   .I4(InputBits[158]),
   .I5(InputBits[1595])
);
LUT6 #(
   .INIT(64'b0010100001010110111100100111100000100011111110011110010000000001)  
) LUT6_572 (
   .O(gates[363]),
   .I0(InputBits[1107]),
   .I1(InputBits[865]),
   .I2(InputBits[1174]),
   .I3(InputBits[549]),
   .I4(InputBits[1609]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1011010001011001001111011111111111011011111001101011000001001101)  
) LUT6_573 (
   .O(gates[46]),
   .I0(InputBits[1339]),
   .I1(InputBits[1303]),
   .I2(InputBits[174]),
   .I3(InputBits[971]),
   .I4(InputBits[1330]),
   .I5(InputBits[1306])
);
LUT6 #(
   .INIT(64'b1000111001001110010110000000011000100110001111001000000100100110)  
) LUT6_574 (
   .O(gates[1316]),
   .I0(InputBits[933]),
   .I1(InputBits[1551]),
   .I2(InputBits[1017]),
   .I3(InputBits[219]),
   .I4(InputBits[932]),
   .I5(InputBits[1633])
);
LUT6 #(
   .INIT(64'b1010001000100110111000101010100101000000100010100100001000100111)  
) LUT6_575 (
   .O(gates[733]),
   .I0(InputBits[1647]),
   .I1(InputBits[841]),
   .I2(InputBits[164]),
   .I3(InputBits[1165]),
   .I4(InputBits[1161]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b0101010000011000001001010001111010011101100110000000010101110001)  
) LUT6_576 (
   .O(gates[36]),
   .I0(InputBits[508]),
   .I1(InputBits[1114]),
   .I2(InputBits[136]),
   .I3(InputBits[448]),
   .I4(InputBits[1714]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0101011001110011100110011110011001000110001110000000111101111100)  
) LUT6_577 (
   .O(gates[1418]),
   .I0(InputBits[1077]),
   .I1(InputBits[1123]),
   .I2(InputBits[246]),
   .I3(InputBits[93]),
   .I4(InputBits[1343]),
   .I5(InputBits[1519])
);
LUT6 #(
   .INIT(64'b0101111110110100100001001001101100001000000001011011000010000110)  
) LUT6_578 (
   .O(gates[997]),
   .I0(InputBits[1372]),
   .I1(InputBits[1257]),
   .I2(InputBits[711]),
   .I3(InputBits[1608]),
   .I4(InputBits[1275]),
   .I5(InputBits[1360])
);
LUT6 #(
   .INIT(64'b1011011110110111110001011010100010110110010011001011110001011010)  
) LUT6_579 (
   .O(gates[630]),
   .I0(InputBits[1170]),
   .I1(InputBits[377]),
   .I2(InputBits[1387]),
   .I3(InputBits[961]),
   .I4(InputBits[1061]),
   .I5(InputBits[1079])
);
LUT6 #(
   .INIT(64'b0001100001011101100001111001001110110101101100001100101111000001)  
) LUT6_580 (
   .O(gates[1368]),
   .I0(InputBits[230]),
   .I1(InputBits[1584]),
   .I2(InputBits[983]),
   .I3(InputBits[893]),
   .I4(InputBits[1414]),
   .I5(InputBits[952])
);
LUT6 #(
   .INIT(64'b0010110011110010010000101111001110001111010000011010100011011101)  
) LUT6_581 (
   .O(gates[472]),
   .I0(InputBits[1166]),
   .I1(InputBits[1496]),
   .I2(InputBits[512]),
   .I3(InputBits[75]),
   .I4(InputBits[996]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0110011011100001001010110110001000100010111100001101101011111111)  
) LUT6_582 (
   .O(gates[748]),
   .I0(InputBits[1554]),
   .I1(InputBits[1630]),
   .I2(InputBits[599]),
   .I3(InputBits[83]),
   .I4(InputBits[589]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0100010100011101001010101100000010001010000011101000110010001001)  
) LUT6_583 (
   .O(gates[1449]),
   .I0(InputBits[255]),
   .I1(InputBits[648]),
   .I2(InputBits[60]),
   .I3(InputBits[1582]),
   .I4(InputBits[1276]),
   .I5(InputBits[1510])
);
LUT6 #(
   .INIT(64'b1100100001111010000011011000010010001001101010100000110000100011)  
) LUT6_584 (
   .O(gates[317]),
   .I0(InputBits[1377]),
   .I1(InputBits[177]),
   .I2(InputBits[518]),
   .I3(InputBits[832]),
   .I4(InputBits[1199]),
   .I5(InputBits[851])
);
LUT6 #(
   .INIT(64'b0000111001110001111110110011000111000100000000100110100011011111)  
) LUT6_585 (
   .O(gates[608]),
   .I0(InputBits[1617]),
   .I1(InputBits[1439]),
   .I2(InputBits[369]),
   .I3(InputBits[1701]),
   .I4(InputBits[1163]),
   .I5(InputBits[1487])
);
LUT6 #(
   .INIT(64'b1011111010000100010011001011011111001011111001100110100111100011)  
) LUT6_586 (
   .O(gates[711]),
   .I0(InputBits[1037]),
   .I1(InputBits[105]),
   .I2(InputBits[870]),
   .I3(InputBits[148]),
   .I4(InputBits[1652]),
   .I5(InputBits[735])
);
LUT6 #(
   .INIT(64'b0101111000010010001001001010011011100000001101011101010000100100)  
) LUT6_587 (
   .O(gates[132]),
   .I0(InputBits[759]),
   .I1(InputBits[531]),
   .I2(InputBits[661]),
   .I3(InputBits[261]),
   .I4(InputBits[905]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b1110000011111001111110111001000010010110111110110011101001111110)  
) LUT6_588 (
   .O(gates[1254]),
   .I0(InputBits[1288]),
   .I1(InputBits[955]),
   .I2(InputBits[1144]),
   .I3(InputBits[790]),
   .I4(InputBits[903]),
   .I5(InputBits[1032])
);
LUT6 #(
   .INIT(64'b0101100110010111010011000001010011111100100011111011110000001011)  
) LUT6_589 (
   .O(gates[1234]),
   .I0(InputBits[1569]),
   .I1(InputBits[53]),
   .I2(InputBits[773]),
   .I3(InputBits[1418]),
   .I4(InputBits[1012]),
   .I5(InputBits[1444])
);
LUT6 #(
   .INIT(64'b1011101111100110011100010000001001110101100101101011100000111111)  
) LUT6_590 (
   .O(gates[892]),
   .I0(InputBits[886]),
   .I1(InputBits[1421]),
   .I2(InputBits[919]),
   .I3(InputBits[1677]),
   .I4(InputBits[1334]),
   .I5(InputBits[859])
);
LUT6 #(
   .INIT(64'b0101001001010010101111000001111100001010000111001101000001110101)  
) LUT6_591 (
   .O(gates[1314]),
   .I0(InputBits[1369]),
   .I1(InputBits[1683]),
   .I2(InputBits[348]),
   .I3(InputBits[719]),
   .I4(InputBits[639]),
   .I5(InputBits[730])
);
LUT6 #(
   .INIT(64'b0001000111101111100101101101010100111110001101001000000110000110)  
) LUT6_592 (
   .O(gates[546]),
   .I0(InputBits[1603]),
   .I1(InputBits[1537]),
   .I2(InputBits[447]),
   .I3(InputBits[1309]),
   .I4(InputBits[1212]),
   .I5(InputBits[633])
);
LUT6 #(
   .INIT(64'b0101101010111011010011001100010011100111100110011110111011000111)  
) LUT6_593 (
   .O(gates[1428]),
   .I0(InputBits[533]),
   .I1(InputBits[223]),
   .I2(InputBits[112]),
   .I3(InputBits[304]),
   .I4(InputBits[784]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b0010000110011111010011000110001010001100110010001011000110111001)  
) LUT6_594 (
   .O(gates[537]),
   .I0(InputBits[579]),
   .I1(InputBits[1561]),
   .I2(InputBits[1221]),
   .I3(InputBits[804]),
   .I4(InputBits[1684]),
   .I5(InputBits[1346])
);
LUT6 #(
   .INIT(64'b1011000100010101101101100000101111110110101100001000111001000101)  
) LUT6_595 (
   .O(gates[1474]),
   .I0(InputBits[1556]),
   .I1(InputBits[879]),
   .I2(InputBits[490]),
   .I3(InputBits[1594]),
   .I4(InputBits[1027]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b0110011001111100011111010010110001111100111010111100101100111100)  
) LUT6_596 (
   .O(gates[125]),
   .I0(InputBits[478]),
   .I1(InputBits[499]),
   .I2(InputBits[173]),
   .I3(InputBits[1230]),
   .I4(InputBits[1669]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b1111000001000001101110111100111010010100110001110001010000100010)  
) LUT6_597 (
   .O(gates[522]),
   .I0(InputBits[1121]),
   .I1(InputBits[1352]),
   .I2(InputBits[1315]),
   .I3(InputBits[30]),
   .I4(InputBits[322]),
   .I5(InputBits[1384])
);
LUT6 #(
   .INIT(64'b1011001010101011010000010010011011111011001110111000011001110011)  
) LUT6_598 (
   .O(gates[1423]),
   .I0(InputBits[1304]),
   .I1(InputBits[1150]),
   .I2(InputBits[1638]),
   .I3(InputBits[672]),
   .I4(InputBits[1686]),
   .I5(InputBits[1464])
);
LUT6 #(
   .INIT(64'b0100001110010110111110000001110101000011000011001111001000101010)  
) LUT6_599 (
   .O(gates[44]),
   .I0(InputBits[614]),
   .I1(InputBits[1703]),
   .I2(InputBits[186]),
   .I3(InputBits[212]),
   .I4(InputBits[563]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b0110101111100100111000000100100001101101001100100111111010111100)  
) LUT6_600 (
   .O(gates[1018]),
   .I0(InputBits[682]),
   .I1(InputBits[133]),
   .I2(InputBits[839]),
   .I3(InputBits[1042]),
   .I4(InputBits[775]),
   .I5(InputBits[1294])
);
LUT6 #(
   .INIT(64'b1000001100110110001000110000111100011101110001101100100010100001)  
) LUT6_601 (
   .O(gates[1125]),
   .I0(InputBits[316]),
   .I1(InputBits[1099]),
   .I2(InputBits[830]),
   .I3(InputBits[1403]),
   .I4(InputBits[277]),
   .I5(InputBits[1240])
);
LUT6 #(
   .INIT(64'b0001101100010111000111000000011110100010001100011110100111010000)  
) LUT6_602 (
   .O(gates[667]),
   .I0(InputBits[1149]),
   .I1(InputBits[1592]),
   .I2(InputBits[1621]),
   .I3(InputBits[1705]),
   .I4(InputBits[5]),
   .I5(InputBits[1645])
);
LUT6 #(
   .INIT(64'b0010011111111010000010010101011001010011111011001100010111111010)  
) LUT6_603 (
   .O(gates[1007]),
   .I0(InputBits[1481]),
   .I1(InputBits[207]),
   .I2(InputBits[613]),
   .I3(InputBits[1525]),
   .I4(InputBits[506]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b1110000100000000100111110000001001001101110111100100011011001100)  
) LUT6_604 (
   .O(gates[1443]),
   .I0(InputBits[1155]),
   .I1(InputBits[949]),
   .I2(InputBits[1243]),
   .I3(InputBits[1397]),
   .I4(InputBits[795]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b1010001110100111010011001100000010111111011110011100011101110100)  
) LUT6_605 (
   .O(gates[741]),
   .I0(InputBits[924]),
   .I1(InputBits[1066]),
   .I2(InputBits[1663]),
   .I3(InputBits[492]),
   .I4(InputBits[25]),
   .I5(InputBits[1719])
);
LUT6 #(
   .INIT(64'b1001111000000101011111101001010100111100001110101111010101001111)  
) LUT6_606 (
   .O(gates[1188]),
   .I0(InputBits[1382]),
   .I1(InputBits[864]),
   .I2(InputBits[591]),
   .I3(InputBits[1602]),
   .I4(InputBits[1290]),
   .I5(InputBits[969])
);
LUT6 #(
   .INIT(64'b0010101000010011000011010100000111001100011000000101110101000101)  
) LUT6_607 (
   .O(gates[1186]),
   .I0(InputBits[927]),
   .I1(InputBits[380]),
   .I2(InputBits[1164]),
   .I3(InputBits[1135]),
   .I4(InputBits[259]),
   .I5(InputBits[1172])
);
LUT6 #(
   .INIT(64'b0001010001111111110001101001110011111000011110010011010001101010)  
) LUT6_608 (
   .O(gates[998]),
   .I0(InputBits[650]),
   .I1(InputBits[1411]),
   .I2(InputBits[658]),
   .I3(InputBits[1253]),
   .I4(InputBits[523]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b1100111001010001100111110101111001110100101111000001100010000011)  
) LUT6_609 (
   .O(gates[714]),
   .I0(InputBits[1470]),
   .I1(InputBits[1449]),
   .I2(InputBits[1385]),
   .I3(InputBits[1517]),
   .I4(InputBits[418]),
   .I5(InputBits[1355])
);
LUT6 #(
   .INIT(64'b0100100110110100011110001111110111100001001011101000001101000100)  
) LUT6_610 (
   .O(gates[1280]),
   .I0(InputBits[436]),
   .I1(InputBits[1472]),
   .I2(InputBits[197]),
   .I3(InputBits[21]),
   .I4(InputBits[1658]),
   .I5(InputBits[1625])
);
LUT6 #(
   .INIT(64'b0001110010000111100011100111110101101111001011101011011100000110)  
) LUT6_611 (
   .O(gates[313]),
   .I0(InputBits[747]),
   .I1(InputBits[1319]),
   .I2(InputBits[1126]),
   .I3(InputBits[203]),
   .I4(InputBits[67]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0001001111100110001000110110100001011101010011001100001111110001)  
) LUT6_612 (
   .O(gates[529]),
   .I0(InputBits[1190]),
   .I1(InputBits[1508]),
   .I2(InputBits[153]),
   .I3(InputBits[665]),
   .I4(InputBits[356]),
   .I5(InputBits[1301])
);
LUT6 #(
   .INIT(64'b0001001111111100100000100010100000110010101110110001001100110000)  
) LUT6_613 (
   .O(gates[1545]),
   .I0(InputBits[973]),
   .I1(InputBits[36]),
   .I2(InputBits[122]),
   .I3(InputBits[1181]),
   .I4(InputBits[479]),
   .I5(InputBits[644])
);
LUT6 #(
   .INIT(64'b1000011111101110010010111100101000111111101011010101111100100101)  
) LUT6_614 (
   .O(gates[1058]),
   .I0(InputBits[845]),
   .I1(InputBits[703]),
   .I2(InputBits[619]),
   .I3(InputBits[474]),
   .I4(InputBits[794]),
   .I5(InputBits[1447])
);
LUT6 #(
   .INIT(64'b1000001110101011011101000001000100101011111101000110011111011111)  
) LUT6_615 (
   .O(gates[987]),
   .I0(InputBits[1197]),
   .I1(InputBits[1168]),
   .I2(InputBits[1558]),
   .I3(InputBits[438]),
   .I4(InputBits[338]),
   .I5(InputBits[91])
);
LUT6 #(
   .INIT(64'b1111000111110110101010101011101110100110101101110000000100110000)  
) LUT6_616 (
   .O(gates[1324]),
   .I0(InputBits[788]),
   .I1(InputBits[1455]),
   .I2(InputBits[963]),
   .I3(InputBits[1489]),
   .I4(InputBits[553]),
   .I5(InputBits[821])
);
LUT6 #(
   .INIT(64'b1010100001001111111001010111011011010101111001010010101111101110)  
) LUT6_617 (
   .O(gates[397]),
   .I0(InputBits[428]),
   .I1(InputBits[1545]),
   .I2(InputBits[468]),
   .I3(InputBits[422]),
   .I4(InputBits[199]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b0111000011111000011101001001100110010100011100111100110110110110)  
) LUT6_618 (
   .O(gates[1150]),
   .I0(InputBits[270]),
   .I1(InputBits[114]),
   .I2(InputBits[397]),
   .I3(InputBits[538]),
   .I4(InputBits[1475]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b1001100000011001100101111001100011001000001011101011001001001111)  
) LUT6_619 (
   .O(gates[1096]),
   .I0(InputBits[1298]),
   .I1(InputBits[1040]),
   .I2(InputBits[59]),
   .I3(InputBits[663]),
   .I4(InputBits[761]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0111001111010101000101000111010111100000110000001111001111000000)  
) LUT6_620 (
   .O(gates[1535]),
   .I0(InputBits[404]),
   .I1(InputBits[520]),
   .I2(InputBits[426]),
   .I3(InputBits[1696]),
   .I4(InputBits[990]),
   .I5(InputBits[1206])
);
LUT6 #(
   .INIT(64'b0111010110100111110101000001000100001111011001111101000111001011)  
) LUT6_621 (
   .O(gates[1335]),
   .I0(InputBits[1441]),
   .I1(InputBits[319]),
   .I2(InputBits[1650]),
   .I3(InputBits[526]),
   .I4(InputBits[248]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b0000101110010111101101000011000001011000100111000010000011011011)  
) LUT6_622 (
   .O(gates[908]),
   .I0(InputBits[967]),
   .I1(InputBits[753]),
   .I2(InputBits[12]),
   .I3(InputBits[896]),
   .I4(InputBits[221]),
   .I5(InputBits[1010])
);
LUT6 #(
   .INIT(64'b0001010100111000110100011111101111000010100101111100101101111011)  
) LUT6_623 (
   .O(gates[1191]),
   .I0(InputBits[603]),
   .I1(InputBits[1492]),
   .I2(InputBits[1021]),
   .I3(InputBits[637]),
   .I4(InputBits[1112]),
   .I5(InputBits[807])
);
LUT6 #(
   .INIT(64'b0011101100100010101100001111100100001001001100101111100110111100)  
) LUT6_624 (
   .O(gates[459]),
   .I0(InputBits[860]),
   .I1(InputBits[1028]),
   .I2(InputBits[1241]),
   .I3(InputBits[1034]),
   .I4(InputBits[440]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b0100000001101101101000000001101001001100010111000001000010000101)  
) LUT6_625 (
   .O(gates[284]),
   .I0(InputBits[1259]),
   .I1(InputBits[801]),
   .I2(InputBits[101]),
   .I3(InputBits[279]),
   .I4(InputBits[587]),
   .I5(InputBits[655])
);
LUT6 #(
   .INIT(64'b0111101011000101010110111011001000010000111000001010001001001100)  
) LUT6_626 (
   .O(gates[823]),
   .I0(InputBits[109]),
   .I1(InputBits[1656]),
   .I2(InputBits[1103]),
   .I3(InputBits[1178]),
   .I4(InputBits[912]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b0011000111101010001100100100001011011011110110101101000101110000)  
) LUT6_627 (
   .O(gates[903]),
   .I0(InputBits[1225]),
   .I1(InputBits[771]),
   .I2(InputBits[626]),
   .I3(InputBits[389]),
   .I4(InputBits[1534]),
   .I5(InputBits[674])
);
LUT6 #(
   .INIT(64'b1110110000011011000101100101001011010011100010101001011000100100)  
) LUT6_628 (
   .O(gates[247]),
   .I0(InputBits[27]),
   .I1(InputBits[881]),
   .I2(InputBits[1287]),
   .I3(InputBits[44]),
   .I4(InputBits[1458]),
   .I5(InputBits[751])
);
LUT6 #(
   .INIT(64'b1110101011000001100100001010011011011110000111011011000110011111)  
) LUT6_629 (
   .O(gates[1340]),
   .I0(InputBits[1345]),
   .I1(InputBits[1035]),
   .I2(InputBits[828]),
   .I3(InputBits[1559]),
   .I4(InputBits[1097]),
   .I5(InputBits[782])
);
LUT6 #(
   .INIT(64'b0000001001110011000011001011101001000100000000100111110010011101)  
) LUT6_630 (
   .O(gates[165]),
   .I0(InputBits[728]),
   .I1(InputBits[1048]),
   .I2(InputBits[688]),
   .I3(InputBits[1131]),
   .I4(InputBits[852]),
   .I5(InputBits[1327])
);
LUT6 #(
   .INIT(64'b0010011011111110011111000011111010001000111111110000010111110011)  
) LUT6_631 (
   .O(gates[289]),
   .I0(InputBits[1679]),
   .I1(InputBits[107]),
   .I2(InputBits[544]),
   .I3(InputBits[1140]),
   .I4(InputBits[921]),
   .I5(InputBits[1433])
);
LUT6 #(
   .INIT(64'b1101110011110000101011000111011001000101110111010000101111101011)  
) LUT6_632 (
   .O(gates[1495]),
   .I0(InputBits[32]),
   .I1(InputBits[366]),
   .I2(InputBits[4]),
   .I3(InputBits[1311]),
   .I4(InputBits[1662]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b0001011111000101011100001111110101110101010001011111011111000110)  
) LUT6_633 (
   .O(gates[729]),
   .I0(InputBits[146]),
   .I1(InputBits[305]),
   .I2(InputBits[561]),
   .I3(InputBits[888]),
   .I4(InputBits[695]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b1100101110111101000001011011100100100000111101111111010001000110)  
) LUT6_634 (
   .O(gates[2]),
   .I0(InputBits[346]),
   .I1(InputBits[382]),
   .I2(InputBits[675]),
   .I3(InputBits[330]),
   .I4(InputBits[1210]),
   .I5(InputBits[1350])
);
LUT6 #(
   .INIT(64'b0100101100011111001100100110000011010010111011110111111010101010)  
) LUT6_635 (
   .O(gates[771]),
   .I0(InputBits[262]),
   .I1(InputBits[744]),
   .I2(InputBits[1265]),
   .I3(InputBits[1053]),
   .I4(InputBits[1059]),
   .I5(InputBits[1152])
);
LUT6 #(
   .INIT(64'b0101101000100010111010101100010111111100111001100010101100101101)  
) LUT6_636 (
   .O(gates[808]),
   .I0(InputBits[1262]),
   .I1(InputBits[1499]),
   .I2(InputBits[1068]),
   .I3(InputBits[694]),
   .I4(InputBits[302]),
   .I5(InputBits[868])
);
LUT6 #(
   .INIT(64'b1100010100001110110111111101010111001110110000101011111101011111)  
) LUT6_637 (
   .O(gates[401]),
   .I0(InputBits[50]),
   .I1(InputBits[352]),
   .I2(InputBits[876]),
   .I3(InputBits[1615]),
   .I4(InputBits[390]),
   .I5(InputBits[1605])
);
LUT6 #(
   .INIT(64'b0000101110101100101100100010111110001000110000010001111000001110)  
) LUT6_638 (
   .O(gates[845]),
   .I0(InputBits[1565]),
   .I1(InputBits[1724]),
   .I2(InputBits[766]),
   .I3(InputBits[433]),
   .I4(InputBits[1580]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0111000111000001110111011001011010011000100100110111111010100000)  
) LUT6_639 (
   .O(gates[186]),
   .I0(InputBits[1527]),
   .I1(InputBits[1465]),
   .I2(InputBits[721]),
   .I3(InputBits[1707]),
   .I4(InputBits[19]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0110111100110000100111100010011110000110010110100111101000110110)  
) LUT6_640 (
   .O(gates[1231]),
   .I0(InputBits[1219]),
   .I1(InputBits[1479]),
   .I2(InputBits[1208]),
   .I3(InputBits[216]),
   .I4(InputBits[1416]),
   .I5(InputBits[1434])
);
LUT6 #(
   .INIT(64'b1110001001000100001101001100000110111100000111001100100001111111)  
) LUT6_641 (
   .O(gates[1119]),
   .I0(InputBits[1336]),
   .I1(InputBits[854]),
   .I2(InputBits[1278]),
   .I3(InputBits[169]),
   .I4(InputBits[1089]),
   .I5(InputBits[593])
);
LUT6 #(
   .INIT(64'b0000000101111001101001011111101100111001001001110001110101101100)  
) LUT6_642 (
   .O(gates[147]),
   .I0(InputBits[210]),
   .I1(InputBits[1408]),
   .I2(InputBits[1600]),
   .I3(InputBits[1389]),
   .I4(InputBits[1404]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1001001000100100010000011010111011000001010101110110101111111110)  
) LUT6_643 (
   .O(gates[1249]),
   .I0(InputBits[1589]),
   .I1(InputBits[1095]),
   .I2(InputBits[288]),
   .I3(InputBits[1725]),
   .I4(InputBits[1370]),
   .I5(InputBits[1435])
);
LUT6 #(
   .INIT(64'b1011110000010000010100110010000011111110000011001011110110011000)  
) LUT6_644 (
   .O(gates[973]),
   .I0(InputBits[1071]),
   .I1(InputBits[358]),
   .I2(InputBits[684]),
   .I3(InputBits[1474]),
   .I4(InputBits[1157]),
   .I5(InputBits[837])
);
LUT6 #(
   .INIT(64'b1111101011111111010110001101001000001101010001101000011101101110)  
) LUT6_645 (
   .O(gates[1046]),
   .I0(InputBits[7]),
   .I1(InputBits[324]),
   .I2(InputBits[269]),
   .I3(InputBits[645]),
   .I4(InputBits[726]),
   .I5(InputBits[1362])
);
LUT6 #(
   .INIT(64'b1000000110111001010011011101110010111101111011110110001110011100)  
) LUT6_646 (
   .O(gates[1142]),
   .I0(InputBits[2]),
   .I1(InputBits[314]),
   .I2(InputBits[1635]),
   .I3(InputBits[1502]),
   .I4(InputBits[787]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b1001111110010101000101101001000010010001111111111011000101101011)  
) LUT6_647 (
   .O(gates[1291]),
   .I0(InputBits[749]),
   .I1(InputBits[1321]),
   .I2(InputBits[786]),
   .I3(InputBits[580]),
   .I4(InputBits[1249]),
   .I5(InputBits[1292])
);
LUT6 #(
   .INIT(64'b1100110110111100000111111010111110111001100110110101111100111010)  
) LUT6_648 (
   .O(gates[319]),
   .I0(InputBits[1678]),
   .I1(InputBits[1460]),
   .I2(InputBits[365]),
   .I3(InputBits[276]),
   .I4(InputBits[910]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1001011011100010011110010110011011100001010001011001110101101101)  
) LUT6_649 (
   .O(gates[915]),
   .I0(InputBits[1310]),
   .I1(InputBits[143]),
   .I2(InputBits[1227]),
   .I3(InputBits[1437]),
   .I4(InputBits[482]),
   .I5(InputBits[1084])
);
LUT6 #(
   .INIT(64'b0011100011110100111011100001000101100110100101011101000101000001)  
) LUT6_650 (
   .O(gates[1179]),
   .I0(InputBits[900]),
   .I1(InputBits[843]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[1087]),
   .I5(InputBits[799])
);
LUT6 #(
   .INIT(64'b0111000010101110011001110010111000100010010101010011001111110011)  
) LUT6_651 (
   .O(gates[1456]),
   .I0(InputBits[70]),
   .I1(InputBits[281]),
   .I2(InputBits[1431]),
   .I3(InputBits[847]),
   .I4(InputBits[1176]),
   .I5(InputBits[1374])
);
LUT6 #(
   .INIT(64'b0010110001101011100001101001001110100001001011011010100011001100)  
) LUT6_652 (
   .O(gates[1052]),
   .I0(InputBits[740]),
   .I1(InputBits[898]),
   .I2(InputBits[286]),
   .I3(InputBits[327]),
   .I4(InputBits[1272]),
   .I5(InputBits[1183])
);
LUT6 #(
   .INIT(64'b1101000001100010111010111101011000111100111110011000110010000100)  
) LUT6_653 (
   .O(gates[404]),
   .I0(InputBits[1466]),
   .I1(InputBits[1031]),
   .I2(InputBits[1203]),
   .I3(InputBits[1610]),
   .I4(InputBits[978]),
   .I5(InputBits[1215])
);
LUT6 #(
   .INIT(64'b1001010011100001010101000010110000101100000010100011011111111011)  
) LUT6_654 (
   .O(gates[735]),
   .I0(InputBits[1086]),
   .I1(InputBits[1115]),
   .I2(InputBits[1532]),
   .I3(InputBits[1452]),
   .I4(InputBits[29]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b0100111001010101010010101010001001000000100011000111100111101100)  
) LUT6_655 (
   .O(gates[516]),
   .I0(InputBits[22]),
   .I1(InputBits[601]),
   .I2(InputBits[17]),
   .I3(InputBits[1296]),
   .I4(InputBits[1417]),
   .I5(InputBits[1574])
);
LUT6 #(
   .INIT(64'b1000010010110011010001010111001001011000101100011010001011001100)  
) LUT6_656 (
   .O(gates[1493]),
   .I0(InputBits[595]),
   .I1(InputBits[451]),
   .I2(InputBits[690]),
   .I3(InputBits[1623]),
   .I4(InputBits[1280]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b0111001111110110100001011011011001010111110110111110001000010001)  
) LUT6_657 (
   .O(gates[974]),
   .I0(InputBits[1314]),
   .I1(InputBits[575]),
   .I2(InputBits[353]),
   .I3(InputBits[170]),
   .I4(InputBits[34]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b0001000110010100000000000000100010110110111011010000110011000101)  
) LUT6_658 (
   .O(gates[1551]),
   .I0(InputBits[995]),
   .I1(InputBits[1237]),
   .I2(InputBits[824]),
   .I3(InputBits[1128]),
   .I4(InputBits[1688]),
   .I5(InputBits[1448])
);
LUT6 #(
   .INIT(64'b1110011111100111011110111001001110100010000000001001011010011101)  
) LUT6_659 (
   .O(gates[702]),
   .I0(InputBits[1064]),
   .I1(InputBits[464]),
   .I2(InputBits[115]),
   .I3(InputBits[455]),
   .I4(InputBits[1110]),
   .I5(InputBits[1279])
);
LUT6 #(
   .INIT(64'b0110100110010001100001101010000011011001001101001110110011101001)  
) LUT6_660 (
   .O(gates[1271]),
   .I0(InputBits[57]),
   .I1(InputBits[913]),
   .I2(InputBits[1727]),
   .I3(InputBits[193]),
   .I4(InputBits[572]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1000000100110001110001111101110011111011011100010111000010010101)  
) LUT6_661 (
   .O(gates[344]),
   .I0(InputBits[628]),
   .I1(InputBits[667]),
   .I2(InputBits[15]),
   .I3(InputBits[1118]),
   .I4(InputBits[345]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b1001011001111000111100010000011011010011000001010011100010001000)  
) LUT6_662 (
   .O(gates[636]),
   .I0(InputBits[1023]),
   .I1(InputBits[116]),
   .I2(InputBits[486]),
   .I3(InputBits[507]),
   .I4(InputBits[1338]),
   .I5(InputBits[1596])
);
LUT6 #(
   .INIT(64'b1001001101000110110101010111001001110111110101111000011101010110)  
) LUT6_663 (
   .O(gates[1104]),
   .I0(InputBits[1506]),
   .I1(InputBits[1246]),
   .I2(InputBits[8]),
   .I3(InputBits[1536]),
   .I4(InputBits[611]),
   .I5(InputBits[1331])
);
LUT6 #(
   .INIT(64'b0001010101000101010111000111111101011110010000100110101111010000)  
) LUT6_664 (
   .O(gates[1406]),
   .I0(InputBits[988]),
   .I1(InputBits[245]),
   .I2(InputBits[1266]),
   .I3(InputBits[546]),
   .I4(InputBits[162]),
   .I5(InputBits[1507])
);
LUT6 #(
   .INIT(64'b1110011010100100011000010110010011010001111000101111000100001101)  
) LUT6_665 (
   .O(gates[561]),
   .I0(InputBits[1002]),
   .I1(InputBits[1160]),
   .I2(InputBits[550]),
   .I3(InputBits[79]),
   .I4(InputBits[1139]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0010000010001111001000100000111111000101100000000100100001001000)  
) LUT6_666 (
   .O(gates[1133]),
   .I0(InputBits[293]),
   .I1(InputBits[621]),
   .I2(InputBits[1236]),
   .I3(InputBits[1159]),
   .I4(InputBits[1102]),
   .I5(InputBits[755])
);
LUT6 #(
   .INIT(64'b0001101000100001000010100000011001001010001101111101110001111001)  
) LUT6_667 (
   .O(gates[209]),
   .I0(InputBits[312]),
   .I1(InputBits[940]),
   .I2(InputBits[931]),
   .I3(InputBits[1497]),
   .I4(InputBits[767]),
   .I5(InputBits[883])
);
LUT6 #(
   .INIT(64'b1000011011110010110011111011000110101000110000010001000001000110)  
) LUT6_668 (
   .O(gates[1118]),
   .I0(InputBits[762]),
   .I1(InputBits[1722]),
   .I2(InputBits[68]),
   .I3(InputBits[1691]),
   .I4(InputBits[950]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b1100000000110101001100111101110010010110011101100001001001000100)  
) LUT6_669 (
   .O(gates[357]),
   .I0(InputBits[1381]),
   .I1(InputBits[654]),
   .I2(InputBits[371]),
   .I3(InputBits[469]),
   .I4(InputBits[819]),
   .I5(InputBits[970])
);
LUT6 #(
   .INIT(64'b0001011101010000100111011000111111001011010000010011110111111001)  
) LUT6_670 (
   .O(gates[117]),
   .I0(InputBits[495]),
   .I1(InputBits[139]),
   .I2(InputBits[343]),
   .I3(InputBits[764]),
   .I4(InputBits[1186]),
   .I5(InputBits[1073])
);
LUT6 #(
   .INIT(64'b1010000110110110111001111110010001011000100110100000110001010010)  
) LUT6_671 (
   .O(gates[1307]),
   .I0(InputBits[915]),
   .I1(InputBits[232]),
   .I2(InputBits[1217]),
   .I3(InputBits[196]),
   .I4(InputBits[696]),
   .I5(InputBits[582])
);
LUT6 #(
   .INIT(64'b0101100101000000101000100000010000001100100110000101100000100011)  
) LUT6_672 (
   .O(gates[455]),
   .I0(InputBits[1628]),
   .I1(InputBits[1260]),
   .I2(InputBits[1524]),
   .I3(InputBits[1239]),
   .I4(InputBits[566]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0010001101100111100111000001111111110011000110110001011011010011)  
) LUT6_673 (
   .O(gates[80]),
   .I0(InputBits[1515]),
   .I1(InputBits[1153]),
   .I2(InputBits[1007]),
   .I3(InputBits[95]),
   .I4(InputBits[1196]),
   .I5(InputBits[1539])
);
LUT6 #(
   .INIT(64'b0000001111111011100001010101011111001000111001010101001011101011)  
) LUT6_674 (
   .O(gates[600]),
   .I0(InputBits[1234]),
   .I1(InputBits[519]),
   .I2(InputBits[984]),
   .I3(InputBits[1295]),
   .I4(InputBits[992]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0110000100000110110001100111100101100001101111010001100001100000)  
) LUT6_675 (
   .O(gates[336]),
   .I0(InputBits[1224]),
   .I1(InputBits[1693]),
   .I2(InputBits[1364]),
   .I3(InputBits[1398]),
   .I4(InputBits[584]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b1101100111001010100110001000101010010011111111101011000100101010)  
) LUT6_676 (
   .O(gates[457]),
   .I0(InputBits[228]),
   .I1(InputBits[373]),
   .I2(InputBits[201]),
   .I3(InputBits[700]),
   .I4(InputBits[81]),
   .I5(InputBits[936])
);
LUT6 #(
   .INIT(64'b1010000101110011101000001000101111101100100111101111001001111001)  
) LUT6_677 (
   .O(gates[1301]),
   .I0(InputBits[504]),
   .I1(InputBits[272]),
   .I2(InputBits[959]),
   .I3(InputBits[811]),
   .I4(InputBits[946]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b0000110001110110011110111111011011111001100100010010100111100000)  
) LUT6_678 (
   .O(gates[821]),
   .I0(InputBits[1550]),
   .I1(InputBits[441]),
   .I2(InputBits[1356]),
   .I3(InputBits[715]),
   .I4(InputBits[220]),
   .I5(InputBits[863])
);
LUT6 #(
   .INIT(64'b1000101110010000000110011010011011101000111001100001011000001101)  
) LUT6_679 (
   .O(gates[383]),
   .I0(InputBits[1577]),
   .I1(InputBits[779]),
   .I2(InputBits[975]),
   .I3(InputBits[510]),
   .I4(InputBits[1401]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b0011000010000111110001010000000000110100101001100111001010000000)  
) LUT6_680 (
   .O(gates[696]),
   .I0(InputBits[1698]),
   .I1(InputBits[834]),
   .I2(InputBits[1009]),
   .I3(InputBits[1690]),
   .I4(InputBits[827]),
   .I5(InputBits[1391])
);
LUT6 #(
   .INIT(64'b1010011000101000101101100000100000100111111000111110011111011011)  
) LUT6_681 (
   .O(gates[297]),
   .I0(InputBits[1093]),
   .I1(InputBits[1080]),
   .I2(InputBits[175]),
   .I3(InputBits[722]),
   .I4(InputBits[798]),
   .I5(InputBits[296])
);
LUT6 #(
   .INIT(64'b1011100001001000010000000011101101010100101000000010100001111010)  
) LUT6_682 (
   .O(gates[963]),
   .I0(InputBits[1643]),
   .I1(InputBits[1660]),
   .I2(InputBits[1075]),
   .I3(InputBits[604]),
   .I4(InputBits[1504]),
   .I5(InputBits[818])
);
LUT6 #(
   .INIT(64'b0101001101010110110001010011010000101111100111001110100101111001)  
) LUT6_683 (
   .O(gates[1431]),
   .I0(InputBits[708]),
   .I1(InputBits[100]),
   .I2(InputBits[388]),
   .I3(InputBits[1708]),
   .I4(InputBits[1318]),
   .I5(InputBits[236])
);
LUT6 #(
   .INIT(64'b0001101101100100001110000001010110011000000110011110010110010101)  
) LUT6_684 (
   .O(gates[92]),
   .I0(InputBits[87]),
   .I1(InputBits[94]),
   .I2(InputBits[671]),
   .I3(InputBits[1323]),
   .I4(InputBits[625]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0111110111110110101111001100001101000101100000011111010111100100)  
) LUT6_685 (
   .O(gates[1489]),
   .I0(InputBits[1214]),
   .I1(InputBits[1193]),
   .I2(InputBits[243]),
   .I3(InputBits[980]),
   .I4(InputBits[77]),
   .I5(InputBits[857])
);
LUT6 #(
   .INIT(64'b0011101011110011000000001000110000001110101000110010111011111100)  
) LUT6_686 (
   .O(gates[1212]),
   .I0(InputBits[132]),
   .I1(InputBits[597]),
   .I2(InputBits[724]),
   .I3(InputBits[278]),
   .I4(InputBits[1587]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0011000000111100111111111010001011111100111001010001001111111000)  
) LUT6_687 (
   .O(gates[10]),
   .I0(InputBits[1251]),
   .I1(InputBits[1564]),
   .I2(InputBits[1307]),
   .I3(InputBits[9]),
   .I4(InputBits[234]),
   .I5(InputBits[1477])
);
LUT6 #(
   .INIT(64'b0111001010101000100100101001101100100110100100001011010001111011)  
) LUT6_688 (
   .O(gates[980]),
   .I0(InputBits[685]),
   .I1(InputBits[462]),
   .I2(InputBits[1108]),
   .I3(InputBits[1637]),
   .I4(InputBits[521]),
   .I5(InputBits[1468])
);
LUT6 #(
   .INIT(64'b0000010000001010111100100010011101101001001110011101000001100010)  
) LUT6_689 (
   .O(gates[550]),
   .I0(InputBits[1329]),
   .I1(InputBits[1106]),
   .I2(InputBits[283]),
   .I3(InputBits[218]),
   .I4(InputBits[1611]),
   .I5(InputBits[1018])
);
LUT6 #(
   .INIT(64'b0101001010101100111010101011111000011110000010001111101100111111)  
) LUT6_690 (
   .O(gates[1477]),
   .I0(InputBits[1429]),
   .I1(InputBits[1522]),
   .I2(InputBits[1379]),
   .I3(InputBits[1305]),
   .I4(InputBits[102]),
   .I5(InputBits[1586])
);
LUT6 #(
   .INIT(64'b1011111100011101000001110110111101100011101010010000000010101011)  
) LUT6_691 (
   .O(gates[1164]),
   .I0(InputBits[835]),
   .I1(InputBits[1454]),
   .I2(InputBits[630]),
   .I3(InputBits[1162]),
   .I4(InputBits[1025]),
   .I5(InputBits[1572])
);
LUT6 #(
   .INIT(64'b1001111001000100111100001110100011101010011101111110100110011010)  
) LUT6_692 (
   .O(gates[1081]),
   .I0(InputBits[796]),
   .I1(InputBits[564]),
   .I2(InputBits[198]),
   .I3(InputBits[1632]),
   .I4(InputBits[570]),
   .I5(InputBits[1133])
);
LUT6 #(
   .INIT(64'b0101000101101111101110000000111001011111100010000001010110100101)  
) LUT6_693 (
   .O(gates[505]),
   .I0(InputBits[292]),
   .I1(InputBits[998]),
   .I2(InputBits[242]),
   .I3(InputBits[1424]),
   .I4(InputBits[359]),
   .I5(InputBits[1715])
);
LUT6 #(
   .INIT(64'b1111110100001011101000111011110000001101001011100111011011000101)  
) LUT6_694 (
   .O(gates[670]),
   .I0(InputBits[891]),
   .I1(InputBits[1484]),
   .I2(InputBits[1014]),
   .I3(InputBits[1406]),
   .I4(InputBits[364]),
   .I5(InputBits[1201])
);
LUT6 #(
   .INIT(64'b1101111010000000000110110101001011000111110011110010110000011101)  
) LUT6_695 (
   .O(gates[1094]),
   .I0(InputBits[150]),
   .I1(InputBits[383]),
   .I2(InputBits[1445]),
   .I3(InputBits[540]),
   .I4(InputBits[1672]),
   .I5(InputBits[1046])
);
LUT6 #(
   .INIT(64'b1111001011100001011011110000101000101111001111100100001110000101)  
) LUT6_696 (
   .O(gates[958]),
   .I0(InputBits[1044]),
   .I1(InputBits[1405]),
   .I2(InputBits[1552]),
   .I3(InputBits[1423]),
   .I4(InputBits[31]),
   .I5(InputBits[1016])
);
LUT6 #(
   .INIT(64'b1111111111010000111010010001000011101000101000001010111101001000)  
) LUT6_697 (
   .O(gates[419]),
   .I0(InputBits[431]),
   .I1(InputBits[1302]),
   .I2(InputBits[1051]),
   .I3(InputBits[367]),
   .I4(InputBits[1493]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b1100100000101011001010111011001000010011001101001100000100100000)  
) LUT6_698 (
   .O(gates[995]),
   .I0(InputBits[258]),
   .I1(InputBits[1393]),
   .I2(InputBits[842]),
   .I3(InputBits[505]),
   .I4(InputBits[1074]),
   .I5(InputBits[113])
);
LUT6 #(
   .INIT(64'b0010001111100110111001110001111100010110100111110001001000001010)  
) LUT6_699 (
   .O(gates[1225]),
   .I0(InputBits[160]),
   .I1(InputBits[742]),
   .I2(InputBits[608]),
   .I3(InputBits[659]),
   .I4(InputBits[58]),
   .I5(InputBits[1349])
);
LUT6 #(
   .INIT(64'b0100001110011100110010101111011111000001011110000011000110101100)  
) LUT6_700 (
   .O(gates[837]),
   .I0(InputBits[548]),
   .I1(InputBits[1394]),
   .I2(InputBits[791]),
   .I3(InputBits[155]),
   .I4(InputBits[640]),
   .I5(InputBits[669])
);
LUT6 #(
   .INIT(64'b1001101000111100111110010110101010111000001111110000111100000000)  
) LUT6_701 (
   .O(gates[290]),
   .I0(InputBits[557]),
   .I1(InputBits[866]),
   .I2(InputBits[350]),
   .I3(InputBits[666]),
   .I4(InputBits[1282]),
   .I5(InputBits[1000])
);
LUT6 #(
   .INIT(64'b1001001100111001000000100011011010101001000111010000000110101101)  
) LUT6_702 (
   .O(gates[592]),
   .I0(InputBits[1648]),
   .I1(InputBits[1427]),
   .I2(InputBits[20]),
   .I3(InputBits[257]),
   .I4(InputBits[1681]),
   .I5(InputBits[873])
);
LUT6 #(
   .INIT(64'b0111111101000100101110100101000100100000110000111011000000011001)  
) LUT6_703 (
   .O(gates[149]),
   .I0(InputBits[386]),
   .I1(InputBits[214]),
   .I2(InputBits[1271]),
   .I3(InputBits[652]),
   .I4(InputBits[920]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b1010111111100101011100101111100110101110100110010110101101000101)  
) LUT6_704 (
   .O(gates[625]),
   .I0(InputBits[917]),
   .I1(InputBits[118]),
   .I2(InputBits[577]),
   .I3(InputBits[977]),
   .I4(InputBits[1626]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0101111101100110000001101001101000110011101011101010110011001000)  
) LUT6_705 (
   .O(gates[712]),
   .I0(InputBits[1057]),
   .I1(InputBits[166]),
   .I2(InputBits[942]),
   .I3(InputBits[624]),
   .I4(InputBits[617]),
   .I5(InputBits[476])
);
LUT6 #(
   .INIT(64'b1110000001011111011000100100100100010101001011001000010001000000)  
) LUT6_706 (
   .O(gates[210]),
   .I0(InputBits[1495]),
   .I1(InputBits[717]),
   .I2(InputBits[334]),
   .I3(InputBits[1137]),
   .I4(InputBits[698]),
   .I5(InputBits[1091])
);
LUT6 #(
   .INIT(64'b1000001010101011000100100001100111010000001001010111111000000011)  
) LUT6_707 (
   .O(gates[406]),
   .I0(InputBits[878]),
   .I1(InputBits[41]),
   .I2(InputBits[1232]),
   .I3(InputBits[250]),
   .I4(InputBits[1671]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b1010110100010110101110110100010000111101100100001001001100111110)  
) LUT6_708 (
   .O(gates[173]),
   .I0(InputBits[172]),
   .I1(InputBits[1367]),
   .I2(InputBits[542]),
   .I3(InputBits[1142]),
   .I4(InputBits[1269]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0000111110110011000001011110101101110111111001100111101110001001)  
) LUT6_709 (
   .O(gates[530]),
   .I0(InputBits[1184]),
   .I1(InputBits[181]),
   .I2(InputBits[14]),
   .I3(InputBits[623]),
   .I4(InputBits[460]),
   .I5(InputBits[1354])
);
LUT6 #(
   .INIT(64'b1101101010110000101001100110011001000011100100100100100001011000)  
) LUT6_710 (
   .O(gates[66]),
   .I0(InputBits[1653]),
   .I1(InputBits[987]),
   .I2(InputBits[423]),
   .I3(InputBits[568]),
   .I4(InputBits[809]),
   .I5(InputBits[734])
);
LUT6 #(
   .INIT(64'b0111101110000100101011110100101000111011100011100100110000100011)  
) LUT6_711 (
   .O(gates[19]),
   .I0(InputBits[1005]),
   .I1(InputBits[85]),
   .I2(InputBits[1728]),
   .I3(InputBits[757]),
   .I4(InputBits[1154]),
   .I5(InputBits[1512])
);
LUT6 #(
   .INIT(64'b0101010111000111001110101110010001100101011110010111000001101001)  
) LUT6_712 (
   .O(gates[1030]),
   .I0(InputBits[1541]),
   .I1(InputBits[1120]),
   .I2(InputBits[1147]),
   .I3(InputBits[1175]),
   .I4(InputBits[1700]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0010010010101111100100010011001001001111110101101000010111110101)  
) LUT6_713 (
   .O(gates[365]),
   .I0(InputBits[1038]),
   .I1(InputBits[1641]),
   .I2(InputBits[1575]),
   .I3(InputBits[466]),
   .I4(InputBits[805]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1110010001010010111000100010100011011111101101011110100110111001)  
) LUT6_714 (
   .O(gates[763]),
   .I0(InputBits[1365]),
   .I1(InputBits[141]),
   .I2(InputBits[1613]),
   .I3(InputBits[848]),
   .I4(InputBits[483]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b1110101100001101110010111001111100101101001001000011111111100011)  
) LUT6_715 (
   .O(gates[470]),
   .I0(InputBits[1568]),
   .I1(InputBits[706]),
   .I2(InputBits[493]),
   .I3(InputBits[1555]),
   .I4(InputBits[536]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b1100111010011111101101110101100100100100110100001011011101010010)  
) LUT6_716 (
   .O(gates[1524]),
   .I0(InputBits[777]),
   .I1(InputBits[416]),
   .I2(InputBits[1375]),
   .I3(InputBits[803]),
   .I4(InputBits[943]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b0000010100110111111111011111011110100000111110110110000001001001)  
) LUT6_717 (
   .O(gates[793]),
   .I0(InputBits[189]),
   .I1(InputBits[692]),
   .I2(InputBits[1619]),
   .I3(InputBits[1562]),
   .I4(InputBits[1312]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0111000100100110010101001001110111100111111111000110110010000000)  
) LUT6_718 (
   .O(gates[1205]),
   .I0(InputBits[1316]),
   .I1(InputBits[308]),
   .I2(InputBits[1720]),
   .I3(InputBits[1358]),
   .I4(InputBits[908]),
   .I5(InputBits[745])
);
LUT6 #(
   .INIT(64'b1011110110101010011110011111101010000010101111001001100110001000)  
) LUT6_719 (
   .O(gates[1287]),
   .I0(InputBits[925]),
   .I1(InputBits[938]),
   .I2(InputBits[92]),
   .I3(InputBits[341]),
   .I4(InputBits[1340]),
   .I5(InputBits[825])
);
LUT6 #(
   .INIT(64'b1010011100010111001110010011001101010101000100011011001101111000)  
) LUT6_720 (
   .O(gates[654]),
   .I0(InputBits[813]),
   .I1(InputBits[131]),
   .I2(InputBits[400]),
   .I3(InputBits[1710]),
   .I4(InputBits[1222]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b1100110000010111001011111111100010101100001001101100011001010100)  
) LUT6_721 (
   .O(gates[570]),
   .I0(InputBits[1229]),
   .I1(InputBits[119]),
   .I2(InputBits[1639]),
   .I3(InputBits[679]),
   .I4(InputBits[104]),
   .I5(InputBits[1191])
);
LUT6 #(
   .INIT(64'b1100110110010111010011110000001111100101100100100100110111010101)  
) LUT6_722 (
   .O(gates[252]),
   .I0(InputBits[240]),
   .I1(InputBits[1482]),
   .I2(InputBits[673]),
   .I3(InputBits[515]),
   .I4(InputBits[1245]),
   .I5(InputBits[618])
);
LUT6 #(
   .INIT(64'b1101011100100110000010000001110010001000010100001011000001010101)  
) LUT6_723 (
   .O(gates[1159]),
   .I0(InputBits[213]),
   .I1(InputBits[1194]),
   .I2(InputBits[968]),
   .I3(InputBits[1718]),
   .I4(InputBits[840]),
   .I5(InputBits[810])
);
LUT6 #(
   .INIT(64'b0110111101100100001111001110100011101000010000001110111110101111)  
) LUT6_724 (
   .O(gates[883]),
   .I0(InputBits[134]),
   .I1(InputBits[306]),
   .I2(InputBits[752]),
   .I3(InputBits[434]),
   .I4(InputBits[1270]),
   .I5(InputBits[1151])
);
LUT6 #(
   .INIT(64'b0100111100110010000101100101001110100001110110001011100000101100)  
) LUT6_725 (
   .O(gates[283]),
   .I0(InputBits[606]),
   .I1(InputBits[1342]),
   .I2(InputBits[605]),
   .I3(InputBits[578]),
   .I4(InputBits[99]),
   .I5(InputBits[895])
);
LUT6 #(
   .INIT(64'b0001100100011000001100000010001111000110110110010110111111000010)  
) LUT6_726 (
   .O(gates[156]),
   .I0(InputBits[1713]),
   .I1(InputBits[1461]),
   .I2(InputBits[315]),
   .I3(InputBits[994]),
   .I4(InputBits[681]),
   .I5(InputBits[1674])
);
LUT6 #(
   .INIT(64'b1100010100111010001000110001110001100100110001110110110001111001)  
) LUT6_727 (
   .O(gates[655]),
   .I0(InputBits[1291]),
   .I1(InputBits[911]),
   .I2(InputBits[1591]),
   .I3(InputBits[1300]),
   .I4(InputBits[1188]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b0000101001110111101010111000101100100000011000010000111101101001)  
) LUT6_728 (
   .O(gates[421]),
   .I0(InputBits[1721]),
   .I1(InputBits[1453]),
   .I2(InputBits[465]),
   .I3(InputBits[590]),
   .I4(InputBits[1020]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0101111010001011001101011000110011010100101101101111100100001001)  
) LUT6_729 (
   .O(gates[59]),
   .I0(InputBits[649]),
   .I1(InputBits[1067]),
   .I2(InputBits[1469]),
   .I3(InputBits[1244]),
   .I4(InputBits[237]),
   .I5(InputBits[1335])
);
LUT6 #(
   .INIT(64'b0100111101101010000100100011100011001010110000010011010010101001)  
) LUT6_730 (
   .O(gates[1367]),
   .I0(InputBits[217]),
   .I1(InputBits[769]),
   .I2(InputBits[662]),
   .I3(InputBits[778]),
   .I4(InputBits[1119]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1010111110100011011110111101010111000010010001101100011011100000)  
) LUT6_731 (
   .O(gates[271]),
   .I0(InputBits[1601]),
   .I1(InputBits[1173]),
   .I2(InputBits[497]),
   .I3(InputBits[321]),
   .I4(InputBits[1313]),
   .I5(InputBits[1412])
);
LUT6 #(
   .INIT(64'b1000001011101101110011111100100010001010101100101000011111000110)  
) LUT6_732 (
   .O(gates[1226]),
   .I0(InputBits[204]),
   .I1(InputBits[562]),
   .I2(InputBits[419]),
   .I3(InputBits[477]),
   .I4(InputBits[379]),
   .I5(InputBits[981])
);
LUT6 #(
   .INIT(64'b1110010010100101011000011100000100011011000001001010111000000000)  
) LUT6_733 (
   .O(gates[1256]),
   .I0(InputBits[948]),
   .I1(InputBits[646]),
   .I2(InputBits[361]),
   .I3(InputBits[928]),
   .I4(InputBits[1471]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0011001011110110110001011010101000101111101010100101110001010001)  
) LUT6_734 (
   .O(gates[1070]),
   .I0(InputBits[1252]),
   .I1(InputBits[748]),
   .I2(InputBits[1514]),
   .I3(InputBits[137]),
   .I4(InputBits[1125]),
   .I5(InputBits[704])
);
LUT6 #(
   .INIT(64'b1101001100010100101100100101001100011000111010100010101010101000)  
) LUT6_735 (
   .O(gates[1024]),
   .I0(InputBits[1122]),
   .I1(InputBits[1402]),
   .I2(InputBits[290]),
   .I3(InputBits[123]),
   .I4(InputBits[1509]),
   .I5(InputBits[657])
);
LUT6 #(
   .INIT(64'b1100111000001110100100001101100001100010111100010001101000100001)  
) LUT6_736 (
   .O(gates[491]),
   .I0(InputBits[331]),
   .I1(InputBits[1528]),
   .I2(InputBits[266]),
   .I3(InputBits[417]),
   .I4(InputBits[437]),
   .I5(InputBits[1518])
);
LUT6 #(
   .INIT(64'b0010010010101111001001010100011000100001100000000100111010010001)  
) LUT6_737 (
   .O(gates[864]),
   .I0(InputBits[923]),
   .I1(InputBits[287]),
   .I2(InputBits[785]),
   .I3(InputBits[588]),
   .I4(InputBits[710]),
   .I5(InputBits[822])
);
LUT6 #(
   .INIT(64'b1111011000001000000111110010011010111010100001011000001001000111)  
) LUT6_738 (
   .O(gates[219]),
   .I0(InputBits[894]),
   .I1(InputBits[90]),
   .I2(InputBits[574]),
   .I3(InputBits[945]),
   .I4(InputBits[1607]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b1110111100001110111111000111100111101100111011100111000010011100)  
) LUT6_739 (
   .O(gates[1016]),
   .I0(InputBits[1665]),
   .I1(InputBits[1283]),
   .I2(InputBits[200]),
   .I3(InputBits[1256]),
   .I4(InputBits[299]),
   .I5(InputBits[1371])
);
LUT6 #(
   .INIT(64'b0100101001100000111101101111110010100010010001010111001011101011)  
) LUT6_740 (
   .O(gates[13]),
   .I0(InputBits[1124]),
   .I1(InputBits[1344]),
   .I2(InputBits[1386]),
   .I3(InputBits[1490]),
   .I4(InputBits[627]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b1000100100110110001000001010110000011010100011010110001101001010)  
) LUT6_741 (
   .O(gates[799]),
   .I0(InputBits[84]),
   .I1(InputBits[636]),
   .I2(InputBits[1062]),
   .I3(InputBits[1376]),
   .I4(InputBits[339]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b1001000001101101111001100100100101011111011010100010001000001110)  
) LUT6_742 (
   .O(gates[1170]),
   .I0(InputBits[1583]),
   .I1(InputBits[1581]),
   .I2(InputBits[1328]),
   .I3(InputBits[634]),
   .I4(InputBits[732]),
   .I5(InputBits[985])
);
LUT6 #(
   .INIT(64'b0111101111101000110110011001011001010101100101111001011010001010)  
) LUT6_743 (
   .O(gates[105]),
   .I0(InputBits[705]),
   .I1(InputBits[1553]),
   .I2(InputBits[729]),
   .I3(InputBits[1440]),
   .I4(InputBits[157]),
   .I5(InputBits[789])
);
LUT6 #(
   .INIT(64'b1110110000001110001111001100010110111111010001001001100011110111)  
) LUT6_744 (
   .O(gates[1514]),
   .I0(InputBits[1198]),
   .I1(InputBits[997]),
   .I2(InputBits[966]),
   .I3(InputBits[73]),
   .I4(InputBits[906]),
   .I5(InputBits[1631])
);
LUT6 #(
   .INIT(64'b1011100001110110100011100111011011111000111100001010101000100000)  
) LUT6_745 (
   .O(gates[925]),
   .I0(InputBits[1664]),
   .I1(InputBits[880]),
   .I2(InputBits[1029]),
   .I3(InputBits[408]),
   .I4(InputBits[1167]),
   .I5(InputBits[816])
);
LUT6 #(
   .INIT(64'b1010100110010100000100101000000110100001101000000001100000010101)  
) LUT6_746 (
   .O(gates[840]),
   .I0(InputBits[179]),
   .I1(InputBits[964]),
   .I2(InputBits[530]),
   .I3(InputBits[1368]),
   .I4(InputBits[1055]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b1100000011101001101000010001011110011101000011111011010101101010)  
) LUT6_747 (
   .O(gates[597]),
   .I0(InputBits[1675]),
   .I1(InputBits[1395]),
   .I2(InputBits[558]),
   .I3(InputBits[1560]),
   .I4(InputBits[1657]),
   .I5(InputBits[598])
);
LUT6 #(
   .INIT(64'b1110110000110010101111010010110001111010110000110110110001101001)  
) LUT6_748 (
   .O(gates[390]),
   .I0(InputBits[1651]),
   .I1(InputBits[1419]),
   .I2(InputBits[524]),
   .I3(InputBits[850]),
   .I4(InputBits[1013]),
   .I5(InputBits[871])
);
LUT6 #(
   .INIT(64'b1111111000100010101100000000011101110101101110001100010100101100)  
) LUT6_749 (
   .O(gates[111]),
   .I0(InputBits[677]),
   .I1(InputBits[831]),
   .I2(InputBits[758]),
   .I3(InputBits[1286]),
   .I4(InputBits[1570]),
   .I5(InputBits[877])
);
LUT6 #(
   .INIT(64'b1001101110110110010101001000110000101001111110110001100100100101)  
) LUT6_750 (
   .O(gates[1042]),
   .I0(InputBits[687]),
   .I1(InputBits[1274]),
   .I2(InputBits[887]),
   .I3(InputBits[699]),
   .I4(InputBits[432]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b0011000101100100101100101100101101010111100101111100010100100100)  
) LUT6_751 (
   .O(gates[1515]),
   .I0(InputBits[1432]),
   .I1(InputBits[13]),
   .I2(InputBits[1026]),
   .I3(InputBits[252]),
   .I4(InputBits[144]),
   .I5(InputBits[1347])
);
LUT6 #(
   .INIT(64'b0111010100100011111101000010001011111110010101010110001001100001)  
) LUT6_752 (
   .O(gates[38]),
   .I0(InputBits[459]),
   .I1(InputBits[1047]),
   .I2(InputBits[922]),
   .I3(InputBits[265]),
   .I4(InputBits[1538]),
   .I5(InputBits[953])
);
LUT6 #(
   .INIT(64'b1111001110110011000001111000001011000010001000100000100010110100)  
) LUT6_753 (
   .O(gates[408]),
   .I0(InputBits[741]),
   .I1(InputBits[736]),
   .I2(InputBits[632]),
   .I3(InputBits[376]),
   .I4(InputBits[1036]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0001100100111110001110010100010000011110000110111101101000000101)  
) LUT6_754 (
   .O(gates[1411]),
   .I0(InputBits[555]),
   .I1(InputBits[1289]),
   .I2(InputBits[902]),
   .I3(InputBits[247]),
   .I4(InputBits[413]),
   .I5(InputBits[1220])
);
LUT6 #(
   .INIT(64'b1101001111110000110110011111000000000101100110111101101011001011)  
) LUT6_755 (
   .O(gates[1480]),
   .I0(InputBits[1476]),
   .I1(InputBits[1456]),
   .I2(InputBits[689]),
   .I3(InputBits[1308]),
   .I4(InputBits[1593]),
   .I5(InputBits[1113])
);
LUT6 #(
   .INIT(64'b1100100010001111101100000000011111100000001111000010011000011001)  
) LUT6_756 (
   .O(gates[196]),
   .I0(InputBits[1543]),
   .I1(InputBits[1604]),
   .I2(InputBits[1695]),
   .I3(InputBits[718]),
   .I4(InputBits[856]),
   .I5(InputBits[1557])
);
LUT6 #(
   .INIT(64'b1111001001000101111111001001011001001010101000111100100000001110)  
) LUT6_757 (
   .O(gates[945]),
   .I0(InputBits[1614]),
   .I1(InputBits[145]),
   .I2(InputBits[1293]),
   .I3(InputBits[676]),
   .I4(InputBits[1054]),
   .I5(InputBits[406])
);
LUT6 #(
   .INIT(64'b1100100001010101011110001001011010011111000110000111000111100011)  
) LUT6_758 (
   .O(gates[242]),
   .I0(InputBits[1540]),
   .I1(InputBits[1676]),
   .I2(InputBits[488]),
   .I3(InputBits[1706]),
   .I4(InputBits[576]),
   .I5(InputBits[1132])
);
LUT6 #(
   .INIT(64'b1101010101111011100110110110000000001110101111010100101110101101)  
) LUT6_759 (
   .O(gates[1169]),
   .I0(InputBits[783]),
   .I1(InputBits[457]),
   .I2(InputBits[66]),
   .I3(InputBits[1415]),
   .I4(InputBits[347]),
   .I5(InputBits[776])
);
LUT6 #(
   .INIT(64'b0111000100001010111000100110111100110001101111011100111111101111)  
) LUT6_760 (
   .O(gates[559]),
   .I0(InputBits[6]),
   .I1(InputBits[1646]),
   .I2(InputBits[1702]),
   .I3(InputBits[311]),
   .I4(InputBits[329]),
   .I5(InputBits[565])
);
LUT6 #(
   .INIT(64'b1000101101001101100001010011101100010100110100101001101010101000)  
) LUT6_761 (
   .O(gates[32]),
   .I0(InputBits[446]),
   .I1(InputBits[1661]),
   .I2(InputBits[560]),
   .I3(InputBits[303]),
   .I4(InputBits[763]),
   .I5(InputBits[592])
);
LUT6 #(
   .INIT(64'b0000101001110111010000101001011111001001110111111101101101010011)  
) LUT6_762 (
   .O(gates[118]),
   .I0(InputBits[26]),
   .I1(InputBits[1096]),
   .I2(InputBits[49]),
   .I3(InputBits[1171]),
   .I4(InputBits[1480]),
   .I5(InputBits[1209])
);
LUT6 #(
   .INIT(64'b0101011001010111110110100100110010110111010011000011000000000101)  
) LUT6_763 (
   .O(gates[443]),
   .I0(InputBits[1242]),
   .I1(InputBits[1]),
   .I2(InputBits[254]),
   .I3(InputBits[480]),
   .I4(InputBits[1189]),
   .I5(InputBits[653])
);
LUT6 #(
   .INIT(64'b0001100010011001010000010001011010111000100101011101101110001000)  
) LUT6_764 (
   .O(gates[206]),
   .I0(InputBits[176]),
   .I1(InputBits[1004]),
   .I2(InputBits[1644]),
   .I3(InputBits[211]),
   .I4(InputBits[191]),
   .I5(InputBits[1060])
);
LUT6 #(
   .INIT(64'b1011001001101000111001110111000100100001011111100110011001000110)  
) LUT6_765 (
   .O(gates[959]),
   .I0(InputBits[612]),
   .I1(InputBits[425]),
   .I2(InputBits[581]),
   .I3(InputBits[720]),
   .I4(InputBits[1130]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1110100010111001010010000011001100110110101001000101001010110001)  
) LUT6_766 (
   .O(gates[358]),
   .I0(InputBits[1598]),
   .I1(InputBits[1579]),
   .I2(InputBits[1530]),
   .I3(InputBits[1473]),
   .I4(InputBits[1616]),
   .I5(InputBits[1277])
);
LUT6 #(
   .INIT(64'b0000111101100101101000011010010010101100101100000100010001000000)  
) LUT6_767 (
   .O(gates[331]),
   .I0(InputBits[517]),
   .I1(InputBits[1726]),
   .I2(InputBits[1694]),
   .I3(InputBits[1566]),
   .I4(InputBits[647]),
   .I5(InputBits[1716])
);
LUT6 #(
   .INIT(64'b0100011010001101100101001000010010011101101101111111000001001000)  
) LUT6_768 (
   .O(gates[1065]),
   .I0(InputBits[683]),
   .I1(InputBits[313]),
   .I2(InputBits[1599]),
   .I3(InputBits[1069]),
   .I4(InputBits[208]),
   .I5(InputBits[1410])
);
LUT6 #(
   .INIT(64'b1000110100101101111001011011100101001110011001111011001100001100)  
) LUT6_769 (
   .O(gates[737]),
   .I0(InputBits[355]),
   .I1(InputBits[235]),
   .I2(InputBits[323]),
   .I3(InputBits[1207]),
   .I4(InputBits[1521]),
   .I5(InputBits[833])
);
LUT6 #(
   .INIT(64'b1000101011101100001001101011101101111011111010110110010011100110)  
) LUT6_770 (
   .O(gates[580]),
   .I0(InputBits[1383]),
   .I1(InputBits[709]),
   .I2(InputBits[135]),
   .I3(InputBits[1409]),
   .I4(InputBits[1709]),
   .I5(InputBits[1156])
);
LUT6 #(
   .INIT(64'b0100010000101100111100000001111100101101110101011110100110110111)  
) LUT6_771 (
   .O(gates[767]),
   .I0(InputBits[545]),
   .I1(InputBits[427]),
   .I2(InputBits[947]),
   .I3(InputBits[1363]),
   .I4(InputBits[838]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1100100100101101101010010011000100010000001000000000111100000100)  
) LUT6_772 (
   .O(gates[84]),
   .I0(InputBits[1248]),
   .I1(InputBits[1320]),
   .I2(InputBits[1667]),
   .I3(InputBits[1450]),
   .I4(InputBits[285]),
   .I5(InputBits[853])
);
LUT6 #(
   .INIT(64'b1011101111111100000011100110110110110111010101110011001010001000)  
) LUT6_773 (
   .O(gates[805]),
   .I0(InputBits[514]),
   .I1(InputBits[1590]),
   .I2(InputBits[268]),
   .I3(InputBits[500]),
   .I4(InputBits[712]),
   .I5(InputBits[982])
);
LUT6 #(
   .INIT(64'b0001001101101110001001010001111000011110100010100000010101111011)  
) LUT6_774 (
   .O(gates[1020]),
   .I0(InputBits[1396]),
   .I1(InputBits[1255]),
   .I2(InputBits[1649]),
   .I3(InputBits[473]),
   .I4(InputBits[106]),
   .I5(InputBits[1520])
);
LUT6 #(
   .INIT(64'b1110001101111011011011101001110101001110011111011001001100000111)  
) LUT6_775 (
   .O(gates[437]),
   .I0(InputBits[750]),
   .I1(InputBits[1486]),
   .I2(InputBits[51]),
   .I3(InputBits[509]),
   .I4(InputBits[37]),
   .I5(InputBits[378])
);
LUT6 #(
   .INIT(64'b0000110101110000001011100001000101010001001111101011010110011000)  
) LUT6_776 (
   .O(gates[194]),
   .I0(InputBits[202]),
   .I1(InputBits[467]),
   .I2(InputBits[127]),
   .I3(InputBits[525]),
   .I4(InputBits[1226]),
   .I5(InputBits[1442])
);
LUT6 #(
   .INIT(64'b0101011000111010111101010110000101101100010111110011110010100000)  
) LUT6_777 (
   .O(gates[220]),
   .I0(InputBits[861]),
   .I1(InputBits[552]),
   .I2(InputBits[142]),
   .I3(InputBits[43]),
   .I4(InputBits[656]),
   .I5(InputBits[727])
);
LUT6 #(
   .INIT(64'b1001010011101101011111011001101011110110000100000001000101110011)  
) LUT6_778 (
   .O(gates[1312]),
   .I0(InputBits[215]),
   .I1(InputBits[1205]),
   .I2(InputBits[301]),
   .I3(InputBits[974]),
   .I4(InputBits[1180]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b0001111111110011101001100011000110101000100100000010100110110000)  
) LUT6_779 (
   .O(gates[1257]),
   .I0(InputBits[760]),
   .I1(InputBits[802]),
   .I2(InputBits[929]),
   .I3(InputBits[702]),
   .I4(InputBits[889]),
   .I5(InputBits[1104])
);
LUT6 #(
   .INIT(64'b0111011001111000011111101001001111010110010010001000000011001100)  
) LUT6_780 (
   .O(gates[846]),
   .I0(InputBits[1430]),
   .I1(InputBits[793]),
   .I2(InputBits[691]),
   .I3(InputBits[1090]),
   .I4(InputBits[439]),
   .I5(InputBits[1697])
);
LUT6 #(
   .INIT(64'b1011100000110101011011111010101101001110110000110101110100111000)  
) LUT6_781 (
   .O(gates[1021]),
   .I0(InputBits[1078]),
   .I1(InputBits[1655]),
   .I2(InputBits[71]),
   .I3(InputBits[1618]),
   .I4(InputBits[664]),
   .I5(InputBits[586])
);
LUT6 #(
   .INIT(64'b1010101101000100000011000001111111001100100001000010010110110010)  
) LUT6_782 (
   .O(gates[31]),
   .I0(InputBits[904]),
   .I1(InputBits[909]),
   .I2(InputBits[642]),
   .I3(InputBits[161]),
   .I4(InputBits[1299]),
   .I5(InputBits[226])
);
LUT6 #(
   .INIT(64'b1010010111001010011010000111011100100100001010000011011101001101)  
) LUT6_783 (
   .O(gates[1263]),
   .I0(InputBits[108]),
   .I1(InputBits[1333]),
   .I2(InputBits[128]),
   .I3(InputBits[602]),
   .I4(InputBits[56]),
   .I5(InputBits[858])
);
LUT6 #(
   .INIT(64'b0111010110011111001000100111010001011101010101110111110011100001)  
) LUT6_784 (
   .O(gates[934]),
   .I0(InputBits[1011]),
   .I1(InputBits[1491]),
   .I2(InputBits[280]),
   .I3(InputBits[11]),
   .I4(InputBits[829]),
   .I5(InputBits[1326])
);
LUT6 #(
   .INIT(64'b0110100100001101100011011010111100111011100001001001001101001000)  
) LUT6_785 (
   .O(gates[1296]),
   .I0(InputBits[260]),
   .I1(InputBits[1082]),
   .I2(InputBits[534]),
   .I3(InputBits[532]),
   .I4(InputBits[1546]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0001011010000111011110100100111110011001001101101010010011101001)  
) LUT6_786 (
   .O(gates[1553]),
   .I0(InputBits[629]),
   .I1(InputBits[743]),
   .I2(InputBits[1606]),
   .I3(InputBits[1463]),
   .I4(InputBits[808]),
   .I5(InputBits[781])
);
LUT6 #(
   .INIT(64'b1110110111001001101001101000000010010011100000001101000110000111)  
) LUT6_787 (
   .O(gates[948]),
   .I0(InputBits[1353]),
   .I1(InputBits[738]),
   .I2(InputBits[152]),
   .I3(InputBits[956]),
   .I4(InputBits[1548]),
   .I5(InputBits[1049])
);
LUT6 #(
   .INIT(64'b1110000000101110011011100011001010111111111110111010111100010111)  
) LUT6_788 (
   .O(gates[1303]),
   .I0(InputBits[1533]),
   .I1(InputBits[337]),
   .I2(InputBits[635]),
   .I3(InputBits[222]),
   .I4(InputBits[489]),
   .I5(InputBits[991])
);
LUT6 #(
   .INIT(64'b0001000010011001000011100100110110011000000010101011000110100011)  
) LUT6_789 (
   .O(gates[572]),
   .I0(InputBits[1258]),
   .I1(InputBits[939]),
   .I2(InputBits[1169]),
   .I3(InputBits[962]),
   .I4(InputBits[1022]),
   .I5(InputBits[1111])
);
LUT6 #(
   .INIT(64'b0101110110100100011001101110001110101010101010101111011011010011)  
) LUT6_790 (
   .O(gates[968]),
   .I0(InputBits[1457]),
   .I1(InputBits[774]),
   .I2(InputBits[1179]),
   .I3(InputBits[410]),
   .I4(InputBits[45]),
   .I5(InputBits[1685])
);
LUT6 #(
   .INIT(64'b1001101110100110111110110111100111110100011101100101011111001011)  
) LUT6_791 (
   .O(gates[675]),
   .I0(InputBits[185]),
   .I1(InputBits[1425]),
   .I2(InputBits[1098]),
   .I3(InputBits[1195]),
   .I4(InputBits[1101]),
   .I5(InputBits[972])
);
LUT6 #(
   .INIT(64'b1101101000101000011110101110000111110011110011010111010100000001)  
) LUT6_792 (
   .O(gates[1398]),
   .I0(InputBits[993]),
   .I1(InputBits[527]),
   .I2(InputBits[295]),
   .I3(InputBits[1501]),
   .I4(InputBits[1058]),
   .I5(InputBits[1138])
);
LUT6 #(
   .INIT(64'b0111111100011011001100110010001001001101010110000001110111000000)  
) LUT6_793 (
   .O(gates[226]),
   .I0(InputBits[409]),
   .I1(InputBits[1547]),
   .I2(InputBits[1692]),
   .I3(InputBits[1070]),
   .I4(InputBits[1158]),
   .I5(InputBits[1263])
);
LUT6 #(
   .INIT(64'b1101000010010000111100100011011011001001000011111011101111011110)  
) LUT6_794 (
   .O(gates[15]),
   .I0(InputBits[869]),
   .I1(InputBits[916]),
   .I2(InputBits[64]),
   .I3(InputBits[1711]),
   .I4(InputBits[551]),
   .I5(InputBits[1141])
);
LUT6 #(
   .INIT(64'b0011100010011011000101101100001010111100110100110001000100000111)  
) LUT6_795 (
   .O(gates[527]),
   .I0(InputBits[1325]),
   .I1(InputBits[756]),
   .I2(InputBits[1523]),
   .I3(InputBits[643]),
   .I4(InputBits[138]),
   .I5(InputBits[1001])
);
LUT6 #(
   .INIT(64'b0010001101111011100110011010111100000001110011110100010101100100)  
) LUT6_796 (
   .O(gates[431]),
   .I0(InputBits[1392]),
   .I1(InputBits[251]),
   .I2(InputBits[733]),
   .I3(InputBits[183]),
   .I4(InputBits[231]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b1101001011000011101001101011001001001110111001111000111010111111)  
) LUT6_797 (
   .O(gates[1430]),
   .I0(InputBits[294]),
   .I1(InputBits[1399]),
   .I2(InputBits[765]),
   .I3(InputBits[1094]),
   .I4(InputBits[1185]),
   .I5(InputBits[885])
);
LUT6 #(
   .INIT(64'b0100000101110100011110101111010010111110001110111110001010111011)  
) LUT6_798 (
   .O(gates[1145]),
   .I0(InputBits[585]),
   .I1(InputBits[1233]),
   .I2(InputBits[716]),
   .I3(InputBits[1670]),
   .I4(InputBits[812]),
   .I5(InputBits[1218])
);
LUT6 #(
   .INIT(64'b0010111010010111101101000001010000010011001111100001000101000111)  
) LUT6_799 (
   .O(gates[382]),
   .I0(InputBits[1500]),
   .I1(InputBits[1704]),
   .I2(InputBits[445]),
   .I3(InputBits[882]),
   .I4(InputBits[976]),
   .I5(InputBits[890])
);
LUT6 #(
   .INIT(64'b1111010101001111000010110000000001010000110001000111101100111100)  
) LUT6_800 (
   .O(gates[1448]),
   .I0(InputBits[1576]),
   .I1(InputBits[1134]),
   .I2(InputBits[1485]),
   .I3(InputBits[874]),
   .I4(InputBits[1516]),
   .I5(InputBits[1235])
);
LUT6 #(
   .INIT(64'b1011011101110101110011101000011111001000010000111001000100100101)  
) LUT6_801 (
   .O(gates[1506]),
   .I0(InputBits[1717]),
   .I1(InputBits[384]),
   .I2(InputBits[855]),
   .I3(InputBits[424]),
   .I4(InputBits[1542]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b1100101101000110000001011011101011100001101000101011100101100101)  
) LUT6_802 (
   .O(gates[62]),
   .I0(InputBits[1511]),
   .I1(InputBits[374]),
   .I2(InputBits[930]),
   .I3(InputBits[182]),
   .I4(InputBits[393]),
   .I5(InputBits[1588])
);
LUT6 #(
   .INIT(64'b0101010011011011010001001110011100001000100110101111101111111101)  
) LUT6_803 (
   .O(gates[833]),
   .I0(InputBits[403]),
   .I1(InputBits[407]),
   .I2(InputBits[1578]),
   .I3(InputBits[1006]),
   .I4(InputBits[54]),
   .I5(InputBits[415])
);
LUT6 #(
   .INIT(64'b1110011001011000101110111000101011111001100111111010010001010010)  
) LUT6_804 (
   .O(gates[139]),
   .I0(InputBits[836]),
   .I1(InputBits[225]),
   .I2(InputBits[1668]),
   .I3(InputBits[1689]),
   .I4(InputBits[567]),
   .I5(InputBits[1264])
);
LUT6 #(
   .INIT(64'b0110010111111011001101101101110011000010011001100100010000001010)  
) LUT6_805 (
   .O(gates[129]),
   .I0(InputBits[309]),
   .I1(InputBits[725]),
   .I2(InputBits[1659]),
   .I3(InputBits[48]),
   .I4(InputBits[875]),
   .I5(InputBits[678])
);
LUT6 #(
   .INIT(64'b0011010100110000100101001011100111010011010010101000001000011110)  
) LUT6_806 (
   .O(gates[1472]),
   .I0(InputBits[1388]),
   .I1(InputBits[326]),
   .I2(InputBits[1041]),
   .I3(InputBits[826]),
   .I4(InputBits[707]),
   .I5(InputBits[1216])
);
LUT6 #(
   .INIT(64'b1111011010000001111100110100111011010010110100011101100100000100)  
) LUT6_807 (
   .O(gates[548]),
   .I0(InputBits[820]),
   .I1(InputBits[381]),
   .I2(InputBits[701]),
   .I3(InputBits[1204]),
   .I4(InputBits[494]),
   .I5(InputBits[103])
);
LUT6 #(
   .INIT(64'b0110111110111010001100010101101111010111110010100000110100000100)  
) LUT6_808 (
   .O(gates[926]),
   .I0(InputBits[1357]),
   .I1(InputBits[1642]),
   .I2(InputBits[88]),
   .I3(InputBits[957]),
   .I4(InputBits[10]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1001000001110001001010100110001011110111011110101000001111110111)  
) LUT6_809 (
   .O(gates[859]),
   .I0(InputBits[502]),
   .I1(InputBits[241]),
   .I2(InputBits[80]),
   .I3(InputBits[806]),
   .I4(InputBits[1443]),
   .I5(InputBits[620])
);
LUT6 #(
   .INIT(64'b1110100110011101001001100111000100101110100001001001101101101111)  
) LUT6_810 (
   .O(gates[1246]),
   .I0(InputBits[1083]),
   .I1(InputBits[317]),
   .I2(InputBits[935]),
   .I3(InputBits[1008]),
   .I4(InputBits[503]),
   .I5(InputBits[1531])
);
LUT6 #(
   .INIT(64'b1010010101111010101110010111111001100101110110100001111000011011)  
) LUT6_811 (
   .O(gates[1083]),
   .I0(InputBits[78]),
   .I1(InputBits[1088]),
   .I2(InputBits[1322]),
   .I3(InputBits[1380]),
   .I4(InputBits[387]),
   .I5(InputBits[958])
);
LUT6 #(
   .INIT(64'b0111011001000101001101111010000001010110001000011110111001010001)  
) LUT6_812 (
   .O(gates[739]),
   .I0(InputBits[487]),
   .I1(InputBits[450]),
   .I2(InputBits[151]),
   .I3(InputBits[284]),
   .I4(InputBits[1273]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b0010001000011101001111110010100111010010001110111110011110101101)  
) LUT6_813 (
   .O(gates[1110]),
   .I0(InputBits[631]),
   .I1(InputBits[1285]),
   .I2(InputBits[47]),
   .I3(InputBits[452]),
   .I4(InputBits[405]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b1010010011010100101111010101110001110011100110001000110101010010)  
) LUT6_814 (
   .O(gates[1293]),
   .I0(InputBits[800]),
   .I1(InputBits[1228]),
   .I2(InputBits[357]),
   .I3(InputBits[609]),
   .I4(InputBits[737]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b0111011011001110010101101101010000101011101000100101010001000110)  
) LUT6_815 (
   .O(gates[876]),
   .I0(InputBits[1467]),
   .I1(InputBits[125]),
   .I2(InputBits[398]),
   .I3(InputBits[1324]),
   .I4(InputBits[1202]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1110111010010001000101100010110010010110101110011100101111010011)  
) LUT6_816 (
   .O(gates[662]),
   .I0(InputBits[899]),
   .I1(InputBits[522]),
   .I2(InputBits[481]),
   .I3(InputBits[484]),
   .I4(InputBits[192]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b1101011000111110010110010101100110001000000101101001010000011010)  
) LUT6_817 (
   .O(gates[418]),
   .I0(InputBits[1573]),
   .I1(InputBits[1030]),
   .I2(InputBits[69]),
   .I3(InputBits[244]),
   .I4(InputBits[1337]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1111011001111110100101101010110001110100000111110010100111010010)  
) LUT6_818 (
   .O(gates[783]),
   .I0(InputBits[140]),
   .I1(InputBits[979]),
   .I2(InputBits[823]),
   .I3(InputBits[1428]),
   .I4(InputBits[149]),
   .I5(InputBits[1459])
);
LUT6 #(
   .INIT(64'b0111011101110000000000011000001111000010101011000111010011100100)  
) LUT6_819 (
   .O(gates[933]),
   .I0(InputBits[1529]),
   .I1(InputBits[1332]),
   .I2(InputBits[194]),
   .I3(InputBits[897]),
   .I4(InputBits[573]),
   .I5(InputBits[668])
);
LUT6 #(
   .INIT(64'b1101110000000000001110111000101110100111001011111011011001011001)  
) LUT6_820 (
   .O(gates[168]),
   .I0(InputBits[1146]),
   .I1(InputBits[1129]),
   .I2(InputBits[1597]),
   .I3(InputBits[1015]),
   .I4(InputBits[385]),
   .I5(InputBits[754])
);
LUT6 #(
   .INIT(64'b1110000011101110101011000110110110101001100100100011111100110011)  
) LUT6_821 (
   .O(gates[1357]),
   .I0(InputBits[86]),
   .I1(InputBits[360]),
   .I2(InputBits[1407]),
   .I3(InputBits[1109]),
   .I4(InputBits[1182]),
   .I5(InputBits[1629])
);
LUT6 #(
   .INIT(64'b1101010001100001010100001110000010110111110000101101010111011111)  
) LUT6_822 (
   .O(gates[135]),
   .I0(InputBits[513]),
   .I1(InputBits[171]),
   .I2(InputBits[1003]),
   .I3(InputBits[1348]),
   .I4(InputBits[1117]),
   .I5(InputBits[610])
);
LUT6 #(
   .INIT(64'b0011110100000001111110000000100010000001111010000010000000110101)  
) LUT6_823 (
   .O(gates[348]),
   .I0(InputBits[263]),
   .I1(InputBits[792]),
   .I2(InputBits[539]),
   .I3(InputBits[282]),
   .I4(InputBits[159]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b0001100001111111011111011011001100110000011100001100000010100011)  
) LUT6_824 (
   .O(gates[1518]),
   .I0(InputBits[351]),
   .I1(InputBits[1231]),
   .I2(InputBits[1535]),
   .I3(InputBits[117]),
   .I4(InputBits[1422]),
   .I5(InputBits[1680])
);
LUT6 #(
   .INIT(64'b1101000010101110001101001101000111010011110011110011010001000010)  
) LUT6_825 (
   .O(gates[1152]),
   .I0(InputBits[768]),
   .I1(InputBits[770]),
   .I2(InputBits[130]),
   .I3(InputBits[456]),
   .I4(InputBits[336]),
   .I5(InputBits[1494])
);
LUT6 #(
   .INIT(64'b0000010100011001010000100111011010110100101110100001111000110010)  
) LUT6_826 (
   .O(gates[145]),
   .I0(InputBits[1267]),
   .I1(InputBits[1213]),
   .I2(InputBits[713]),
   .I3(InputBits[1478]),
   .I4(InputBits[772]),
   .I5(InputBits[714])
);
LUT6 #(
   .INIT(64'b1011101010101001110101101011100110101100111110110001101011000101)  
) LUT6_827 (
   .O(gates[789]),
   .I0(InputBits[1624]),
   .I1(InputBits[1634]),
   .I2(InputBits[1359]),
   .I3(InputBits[989]),
   .I4(InputBits[1351]),
   .I5(InputBits[986])
);
LUT6 #(
   .INIT(64'b1010100110000110000000010000010000101101110000111011011111101111)  
) LUT6_828 (
   .O(gates[49]),
   .I0(InputBits[1666]),
   .I1(InputBits[1177]),
   .I2(InputBits[1297]),
   .I3(InputBits[600]),
   .I4(InputBits[38]),
   .I5(InputBits[844])
);
LUT6 #(
   .INIT(64'b1000010000011100010011010000000010010001000000110100000000011110)  
) LUT6_829 (
   .O(gates[178]),
   .I0(InputBits[156]),
   .I1(InputBits[1436]),
   .I2(InputBits[1052]),
   .I3(InputBits[1281]),
   .I4(InputBits[547]),
   .I5(InputBits[1024])
);
LUT6 #(
   .INIT(64'b0101010000110001011010000111110011110101000101101011101011111011)  
) LUT6_830 (
   .O(gates[1131]),
   .I0(InputBits[1687]),
   .I1(InputBits[461]),
   .I2(InputBits[1627]),
   .I3(InputBits[1513]),
   .I4(InputBits[165]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0110010100000101010010010010110001111001100001101000111110101101)  
) LUT6_831 (
   .O(gates[124]),
   .I0(InputBits[1498]),
   .I1(InputBits[651]),
   .I2(InputBits[622]),
   .I3(InputBits[333]),
   .I4(InputBits[941]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0010001000001111001010001101111011010011101000101010100101100101)  
) LUT6_832 (
   .O(gates[772]),
   .I0(InputBits[1712]),
   .I1(InputBits[731]),
   .I2(InputBits[814]),
   .I3(InputBits[375]),
   .I4(InputBits[1092]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0111011011110010110101111110111110101111101111001111001110010011)  
) LUT6_833 (
   .O(gates[993]),
   .I0(InputBits[1261]),
   .I1(InputBits[195]),
   .I2(InputBits[253]),
   .I3(InputBits[184]),
   .I4(InputBits[1247]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b1001101100000000110000110101100000000001110001001000111010101111)  
) LUT6_834 (
   .O(gates[1090]),
   .I0(InputBits[496]),
   .I1(InputBits[1127]),
   .I2(InputBits[1268]),
   .I3(InputBits[1446]),
   .I4(InputBits[934]),
   .I5(InputBits[849])
);
LUT6 #(
   .INIT(64'b0011001101110101001100111110011101011000101000110111111001011110)  
) LUT6_835 (
   .O(gates[627]),
   .I0(InputBits[1100]),
   .I1(InputBits[1622]),
   .I2(InputBits[954]),
   .I3(InputBits[1148]),
   .I4(InputBits[1400]),
   .I5(InputBits[616])
);
LUT6 #(
   .INIT(64'b1001011111101010001011001000100110010100010010100100000110010110)  
) LUT6_836 (
   .O(gates[1308]),
   .I0(InputBits[1056]),
   .I1(InputBits[411]),
   .I2(InputBits[454]),
   .I3(InputBits[110]),
   .I4(InputBits[354]),
   .I5(InputBits[1072])
);
LUT6 #(
   .INIT(64'b1010011011111010001111110010111010111000100010110100100011101001)  
) LUT6_837 (
   .O(gates[1429]),
   .I0(InputBits[227]),
   .I1(InputBits[884]),
   .I2(InputBits[1143]),
   .I3(InputBits[697]),
   .I4(InputBits[1187]),
   .I5(InputBits[951])
);
LUT6 #(
   .INIT(64'b1000000100111001000110001110101110001100011110000111010011010001)  
) LUT6_838 (
   .O(gates[715]),
   .I0(InputBits[529]),
   .I1(InputBits[918]),
   .I2(InputBits[1043]),
   .I3(InputBits[1654]),
   .I4(InputBits[1567]),
   .I5(InputBits[615])
);
LUT6 #(
   .INIT(64'b1111000010100000000100010000011111001011000010100000100010000000)  
) LUT6_839 (
   .O(gates[1374]),
   .I0(InputBits[1341]),
   .I1(InputBits[780]),
   .I2(InputBits[867]),
   .I3(InputBits[1366]),
   .I4(InputBits[435]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b1110001111111101011111110111011100010011100100011110111011100101)  
) LUT6_840 (
   .O(gates[23]),
   .I0(InputBits[1699]),
   .I1(InputBits[97]),
   .I2(InputBits[846]),
   .I3(InputBits[1640]),
   .I4(InputBits[937]),
   .I5(InputBits[907])
);
LUT6 #(
   .INIT(64'b0011001101101010000110000111100100011000101010011100100001010000)  
) LUT6_841 (
   .O(gates[388]),
   .I0(InputBits[498]),
   .I1(InputBits[1378]),
   .I2(InputBits[554]),
   .I3(InputBits[154]),
   .I4(InputBits[746]),
   .I5(InputBits[472])
);
LUT6 #(
   .INIT(64'b0011101011000111000101011100011100100110000111101011101101001001)  
) LUT6_842 (
   .O(gates[364]),
   .I0(InputBits[926]),
   .I1(InputBits[914]),
   .I2(InputBits[1317]),
   .I3(InputBits[190]),
   .I4(InputBits[1039]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b0110000001000110001011000101111001000001011101110100001110100001)  
) LUT6_843 (
   .O(gates[1528]),
   .I0(InputBits[535]),
   .I1(InputBits[307]),
   .I2(InputBits[797]),
   .I3(InputBits[569]),
   .I4(InputBits[342]),
   .I5(InputBits[1105])
);
LUT6 #(
   .INIT(64'b0011001000001101011010010001110100100111011110011101110000110111)  
) LUT6_844 (
   .O(gates[653]),
   .I0(InputBits[297]),
   .I1(InputBits[1136]),
   .I2(InputBits[817]),
   .I3(InputBits[1503]),
   .I4(InputBits[401]),
   .I5(InputBits[1390])
);
LUT6 #(
   .INIT(64'b1001101110011101110111111110011010010111111011100100001110110101)  
) LUT6_845 (
   .O(gates[1425]),
   .I0(InputBits[693]),
   .I1(InputBits[1223]),
   .I2(InputBits[680]),
   .I3(InputBits[1620]),
   .I4(InputBits[1526]),
   .I5(InputBits[1254])
);
LUT6 #(
   .INIT(64'b1000100010001000001001101010111001001011010101010110101000100111)  
) LUT6_846 (
   .O(gates[950]),
   .I0(InputBits[1544]),
   .I1(InputBits[1723]),
   .I2(InputBits[1076]),
   .I3(InputBits[723]),
   .I4(InputBits[872]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0001111011000111110101000110100100110000011111111011100100011111)  
) LUT6_847 (
   .O(gates[1445]),
   .I0(InputBits[82]),
   .I1(InputBits[1211]),
   .I2(InputBits[1373]),
   .I3(InputBits[239]),
   .I4(InputBits[638]),
   .I5(InputBits[1081])
);
LUT6 #(
   .INIT(64'b1010001001001111000110101111001001111000100111010010101101100111)  
) LUT6_848 (
   .O(gates[1025]),
   .I0(InputBits[537]),
   .I1(InputBits[1413]),
   .I2(InputBits[944]),
   .I3(InputBits[901]),
   .I4(InputBits[1636]),
   .I5(InputBits[1250])
);
LUT6 #(
   .INIT(64'b1011010111000011110100110000011000100100100110011101010111000001)  
) LUT6_849 (
   .O(gates[509]),
   .I0(InputBits[541]),
   .I1(InputBits[229]),
   .I2(InputBits[1284]),
   .I3(InputBits[124]),
   .I4(InputBits[594]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0111010001100011010111111011101000011100000110100011111010111111)  
) LUT6_850 (
   .O(gates[1015]),
   .I0(InputBits[1462]),
   .I1(InputBits[1085]),
   .I2(InputBits[65]),
   .I3(InputBits[1145]),
   .I4(InputBits[686]),
   .I5(InputBits[1549])
);
LUT6 #(
   .INIT(64'b0011001011100010101000010100001100001011101100001011000100100001)  
) LUT6_851 (
   .O(gates[976]),
   .I0(InputBits[1420]),
   .I1(InputBits[1505]),
   .I2(InputBits[1612]),
   .I3(InputBits[1192]),
   .I4(InputBits[328]),
   .I5(InputBits[607])
);
LUT6 #(
   .INIT(64'b0010100010101000101101100101010000011000111010111110001111010001)  
) LUT6_852 (
   .O(gates[367]),
   .I0(InputBits[815]),
   .I1(InputBits[291]),
   .I2(InputBits[660]),
   .I3(InputBits[1116]),
   .I4(InputBits[370]),
   .I5(InputBits[999])
);
LUT6 #(
   .INIT(64'b0001101001010000011100001001010000110110001001100001011000111010)  
) LUT6_853 (
   .O(gates[716]),
   .I0(InputBits[1019]),
   .I1(InputBits[1361]),
   .I2(InputBits[1571]),
   .I3(InputBits[1045]),
   .I4(InputBits[960]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b1100010100111110011001110000100011011001010001100100111111101001)  
) LUT6_854 (
   .O(gates[940]),
   .I0(InputBits[28]),
   .I1(InputBits[862]),
   .I2(InputBits[76]),
   .I3(InputBits[273]),
   .I4(InputBits[1050]),
   .I5(InputBits[1065])
);
LUT6 #(
   .INIT(64'b0010101100000100010010011101100110100111111001101100010111110100)  
) LUT6_855 (
   .O(gates[1466]),
   .I0(InputBits[739]),
   .I1(InputBits[1451]),
   .I2(InputBits[583]),
   .I3(InputBits[965]),
   .I4(InputBits[892]),
   .I5(InputBits[670])
);
LUT6 #(
   .INIT(64'b1110110111000110100100011101100000010011001010100000010100100110)  
) LUT6_856 (
   .O(gates[485]),
   .I0(InputBits[23]),
   .I1(InputBits[1673]),
   .I2(InputBits[1585]),
   .I3(InputBits[1488]),
   .I4(InputBits[1063]),
   .I5(InputBits[1426])
);
LUT6 #(
   .INIT(64'b1001001111111000101111011000100000001100010010001000111110101110)  
) LUT6_857 (
   .O(gates[743]),
   .I0(InputBits[1483]),
   .I1(InputBits[596]),
   .I2(InputBits[1238]),
   .I3(InputBits[274]),
   .I4(InputBits[362]),
   .I5(InputBits[1033])
);
LUT6 #(
   .INIT(64'b0100010011011101100010100001010111101000011010110010000011111101)  
) LUT6_858 (
   .O(gates[778]),
   .I0(InputBits[1438]),
   .I1(InputBits[349]),
   .I2(InputBits[206]),
   .I3(InputBits[74]),
   .I4(InputBits[363]),
   .I5(InputBits[1200])
);
LUT6 #(
   .INIT(64'b0011100010001011110111100001001111101110010001110000111111001100)  
) LUT6_859 (
   .O(gates[685]),
   .I0(InputBits[641]),
   .I1(InputBits[147]),
   .I2(InputBits[1682]),
   .I3(InputBits[1563]),
   .I4(InputBits[158]),
   .I5(InputBits[1595])
);
LUT6 #(
   .INIT(64'b1100011000000000100000100101101011001001101110000101010110000100)  
) LUT6_860 (
   .O(gates[21]),
   .I0(InputBits[1107]),
   .I1(InputBits[865]),
   .I2(InputBits[1174]),
   .I3(InputBits[549]),
   .I4(InputBits[1609]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b1011011000001000010110101110110100100011101110110011010001000111)  
) LUT6_861 (
   .O(gates[523]),
   .I0(InputBits[1339]),
   .I1(InputBits[1303]),
   .I2(InputBits[174]),
   .I3(InputBits[971]),
   .I4(InputBits[1330]),
   .I5(InputBits[1306])
);
LUT6 #(
   .INIT(64'b0000000010111110110000000001010010001011110000100100001111100110)  
) LUT6_862 (
   .O(gates[720]),
   .I0(InputBits[933]),
   .I1(InputBits[1551]),
   .I2(InputBits[1017]),
   .I3(InputBits[219]),
   .I4(InputBits[932]),
   .I5(InputBits[1633])
);
LUT6 #(
   .INIT(64'b0110111011110011110000000011001001010110100000100100001000011001)  
) LUT6_863 (
   .O(gates[1270]),
   .I0(InputBits[1647]),
   .I1(InputBits[841]),
   .I2(InputBits[164]),
   .I3(InputBits[1165]),
   .I4(InputBits[1161]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b1100110001101110111011110011101101111010011011100101110111110011)  
) LUT6_864 (
   .O(gates[460]),
   .I0(InputBits[508]),
   .I1(InputBits[1114]),
   .I2(InputBits[136]),
   .I3(InputBits[448]),
   .I4(InputBits[1714]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0001000010011000100101010010001100011100000111111000000001100011)  
) LUT6_865 (
   .O(gates[723]),
   .I0(InputBits[1077]),
   .I1(InputBits[1123]),
   .I2(InputBits[246]),
   .I3(InputBits[93]),
   .I4(InputBits[1343]),
   .I5(InputBits[1519])
);
LUT6 #(
   .INIT(64'b0001101011110010111100111011100010000111100110001010100110000111)  
) LUT6_866 (
   .O(gates[324]),
   .I0(InputBits[1372]),
   .I1(InputBits[1257]),
   .I2(InputBits[711]),
   .I3(InputBits[1608]),
   .I4(InputBits[1275]),
   .I5(InputBits[1360])
);
LUT6 #(
   .INIT(64'b0111111000010101000000111000000010101111000011111010110111000110)  
) LUT6_867 (
   .O(gates[453]),
   .I0(InputBits[1170]),
   .I1(InputBits[377]),
   .I2(InputBits[1387]),
   .I3(InputBits[961]),
   .I4(InputBits[1061]),
   .I5(InputBits[1079])
);
LUT6 #(
   .INIT(64'b0110000010110110110000100101000101100100011011101001010011110111)  
) LUT6_868 (
   .O(gates[1389]),
   .I0(InputBits[230]),
   .I1(InputBits[1584]),
   .I2(InputBits[983]),
   .I3(InputBits[893]),
   .I4(InputBits[1414]),
   .I5(InputBits[952])
);
LUT6 #(
   .INIT(64'b0100001011110010110110010001110011000111000110111011010100001011)  
) LUT6_869 (
   .O(gates[1460]),
   .I0(InputBits[1166]),
   .I1(InputBits[1496]),
   .I2(InputBits[512]),
   .I3(InputBits[75]),
   .I4(InputBits[996]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0100110111001000001011010100000110110111010110001011111100111000)  
) LUT6_870 (
   .O(gates[244]),
   .I0(InputBits[1554]),
   .I1(InputBits[1630]),
   .I2(InputBits[599]),
   .I3(InputBits[83]),
   .I4(InputBits[589]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0101101001111000000000010111000000001100100001000011110111100001)  
) LUT6_871 (
   .O(gates[1202]),
   .I0(InputBits[255]),
   .I1(InputBits[648]),
   .I2(InputBits[60]),
   .I3(InputBits[1582]),
   .I4(InputBits[1276]),
   .I5(InputBits[1510])
);
LUT6 #(
   .INIT(64'b1011010100000100100101101011101000001000100010100000101110010111)  
) LUT6_872 (
   .O(gates[637]),
   .I0(InputBits[1377]),
   .I1(InputBits[177]),
   .I2(InputBits[518]),
   .I3(InputBits[832]),
   .I4(InputBits[1199]),
   .I5(InputBits[851])
);
LUT6 #(
   .INIT(64'b1001101101100010110110101101000001101111101001011100100000100100)  
) LUT6_873 (
   .O(gates[351]),
   .I0(InputBits[1617]),
   .I1(InputBits[1439]),
   .I2(InputBits[369]),
   .I3(InputBits[1701]),
   .I4(InputBits[1163]),
   .I5(InputBits[1487])
);
LUT6 #(
   .INIT(64'b0001111011100101000000011010110010111111110011111011101101100010)  
) LUT6_874 (
   .O(gates[1040]),
   .I0(InputBits[1037]),
   .I1(InputBits[105]),
   .I2(InputBits[870]),
   .I3(InputBits[148]),
   .I4(InputBits[1652]),
   .I5(InputBits[735])
);
LUT6 #(
   .INIT(64'b1110100010111010001000110001001100011001011010100010011001111110)  
) LUT6_875 (
   .O(gates[595]),
   .I0(InputBits[759]),
   .I1(InputBits[531]),
   .I2(InputBits[661]),
   .I3(InputBits[261]),
   .I4(InputBits[905]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b1111110100000111110101001100101110100101101101010110101100101011)  
) LUT6_876 (
   .O(gates[1138]),
   .I0(InputBits[1288]),
   .I1(InputBits[955]),
   .I2(InputBits[1144]),
   .I3(InputBits[790]),
   .I4(InputBits[903]),
   .I5(InputBits[1032])
);
LUT6 #(
   .INIT(64'b1100110110101111000111110110110110010110110001100100001100011010)  
) LUT6_877 (
   .O(gates[488]),
   .I0(InputBits[1569]),
   .I1(InputBits[53]),
   .I2(InputBits[773]),
   .I3(InputBits[1418]),
   .I4(InputBits[1012]),
   .I5(InputBits[1444])
);
LUT6 #(
   .INIT(64'b1100011011111001100011110000100011101000111001001101011000000111)  
) LUT6_878 (
   .O(gates[752]),
   .I0(InputBits[886]),
   .I1(InputBits[1421]),
   .I2(InputBits[919]),
   .I3(InputBits[1677]),
   .I4(InputBits[1334]),
   .I5(InputBits[859])
);
LUT6 #(
   .INIT(64'b1001000111101001111110110110100101110100010100001100000011010110)  
) LUT6_879 (
   .O(gates[1012]),
   .I0(InputBits[1369]),
   .I1(InputBits[1683]),
   .I2(InputBits[348]),
   .I3(InputBits[719]),
   .I4(InputBits[639]),
   .I5(InputBits[730])
);
LUT6 #(
   .INIT(64'b1110011011010010010101101001100110000110011110000001110111010011)  
) LUT6_880 (
   .O(gates[1232]),
   .I0(InputBits[1603]),
   .I1(InputBits[1537]),
   .I2(InputBits[447]),
   .I3(InputBits[1309]),
   .I4(InputBits[1212]),
   .I5(InputBits[633])
);
LUT6 #(
   .INIT(64'b0111111100100010010010010001001011100111001110101011111110100100)  
) LUT6_881 (
   .O(gates[1498]),
   .I0(InputBits[533]),
   .I1(InputBits[223]),
   .I2(InputBits[112]),
   .I3(InputBits[304]),
   .I4(InputBits[784]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b1101010110001010001111000111100010101111101101110110101111101110)  
) LUT6_882 (
   .O(gates[835]),
   .I0(InputBits[579]),
   .I1(InputBits[1561]),
   .I2(InputBits[1221]),
   .I3(InputBits[804]),
   .I4(InputBits[1684]),
   .I5(InputBits[1346])
);
LUT6 #(
   .INIT(64'b1101011011001101010001110100101001111010011111010000111001110100)  
) LUT6_883 (
   .O(gates[1267]),
   .I0(InputBits[1556]),
   .I1(InputBits[879]),
   .I2(InputBits[490]),
   .I3(InputBits[1594]),
   .I4(InputBits[1027]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b0110111010101100100110110100111011111000101100010100111110100110)  
) LUT6_884 (
   .O(gates[379]),
   .I0(InputBits[478]),
   .I1(InputBits[499]),
   .I2(InputBits[173]),
   .I3(InputBits[1230]),
   .I4(InputBits[1669]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b0010111000101011001011110001010000010011100010001101100011101000)  
) LUT6_885 (
   .O(gates[1032]),
   .I0(InputBits[1121]),
   .I1(InputBits[1352]),
   .I2(InputBits[1315]),
   .I3(InputBits[30]),
   .I4(InputBits[322]),
   .I5(InputBits[1384])
);
LUT6 #(
   .INIT(64'b0000001011011010111110010110110000101001101101001011000001101000)  
) LUT6_886 (
   .O(gates[1386]),
   .I0(InputBits[1304]),
   .I1(InputBits[1150]),
   .I2(InputBits[1638]),
   .I3(InputBits[672]),
   .I4(InputBits[1686]),
   .I5(InputBits[1464])
);
LUT6 #(
   .INIT(64'b0111101010011000000000100110111110011100010100111101001011100001)  
) LUT6_887 (
   .O(gates[113]),
   .I0(InputBits[614]),
   .I1(InputBits[1703]),
   .I2(InputBits[186]),
   .I3(InputBits[212]),
   .I4(InputBits[563]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b0011100110100100100101011011101000010100000110001001001010100101)  
) LUT6_888 (
   .O(gates[1536]),
   .I0(InputBits[682]),
   .I1(InputBits[133]),
   .I2(InputBits[839]),
   .I3(InputBits[1042]),
   .I4(InputBits[775]),
   .I5(InputBits[1294])
);
LUT6 #(
   .INIT(64'b1111000101111101100011001011000111101110111000001010101010001111)  
) LUT6_889 (
   .O(gates[901]),
   .I0(InputBits[316]),
   .I1(InputBits[1099]),
   .I2(InputBits[830]),
   .I3(InputBits[1403]),
   .I4(InputBits[277]),
   .I5(InputBits[1240])
);
LUT6 #(
   .INIT(64'b0100000001010101000111110011010110101010000100100110100000000111)  
) LUT6_890 (
   .O(gates[1035]),
   .I0(InputBits[1149]),
   .I1(InputBits[1592]),
   .I2(InputBits[1621]),
   .I3(InputBits[1705]),
   .I4(InputBits[5]),
   .I5(InputBits[1645])
);
LUT6 #(
   .INIT(64'b1011100010001100000001001100101100101011101000000101010010111110)  
) LUT6_891 (
   .O(gates[152]),
   .I0(InputBits[1481]),
   .I1(InputBits[207]),
   .I2(InputBits[613]),
   .I3(InputBits[1525]),
   .I4(InputBits[506]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b0001011100010111011111101101001000001010011100000100011000101001)  
) LUT6_892 (
   .O(gates[342]),
   .I0(InputBits[1155]),
   .I1(InputBits[949]),
   .I2(InputBits[1243]),
   .I3(InputBits[1397]),
   .I4(InputBits[795]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b1101111001100101001101010111010000101110001011011010101110001110)  
) LUT6_893 (
   .O(gates[452]),
   .I0(InputBits[924]),
   .I1(InputBits[1066]),
   .I2(InputBits[1663]),
   .I3(InputBits[492]),
   .I4(InputBits[25]),
   .I5(InputBits[1719])
);
LUT6 #(
   .INIT(64'b0100101111010101111011101100111010111001000110010100111111010001)  
) LUT6_894 (
   .O(gates[862]),
   .I0(InputBits[1382]),
   .I1(InputBits[864]),
   .I2(InputBits[591]),
   .I3(InputBits[1602]),
   .I4(InputBits[1290]),
   .I5(InputBits[969])
);
LUT6 #(
   .INIT(64'b0110101101110011001101001010100110100111101011000000111010010010)  
) LUT6_895 (
   .O(gates[1419]),
   .I0(InputBits[927]),
   .I1(InputBits[380]),
   .I2(InputBits[1164]),
   .I3(InputBits[1135]),
   .I4(InputBits[259]),
   .I5(InputBits[1172])
);
LUT6 #(
   .INIT(64'b1011000100011101000010111100001111000000001010111001111100011100)  
) LUT6_896 (
   .O(gates[579]),
   .I0(InputBits[650]),
   .I1(InputBits[1411]),
   .I2(InputBits[658]),
   .I3(InputBits[1253]),
   .I4(InputBits[523]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b0100100011101111001101000010111010111111001101111001100101110101)  
) LUT6_897 (
   .O(gates[295]),
   .I0(InputBits[1470]),
   .I1(InputBits[1449]),
   .I2(InputBits[1385]),
   .I3(InputBits[1517]),
   .I4(InputBits[418]),
   .I5(InputBits[1355])
);
LUT6 #(
   .INIT(64'b0001111000011010011010011000010000100011010101011100110011101100)  
) LUT6_898 (
   .O(gates[341]),
   .I0(InputBits[436]),
   .I1(InputBits[1472]),
   .I2(InputBits[197]),
   .I3(InputBits[21]),
   .I4(InputBits[1658]),
   .I5(InputBits[1625])
);
LUT6 #(
   .INIT(64'b0001101010111000101011100000011110010111000010000000010000100001)  
) LUT6_899 (
   .O(gates[1056]),
   .I0(InputBits[747]),
   .I1(InputBits[1319]),
   .I2(InputBits[1126]),
   .I3(InputBits[203]),
   .I4(InputBits[67]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b1000000111000101010110011101100101010101100111101000100010111101)  
) LUT6_900 (
   .O(gates[535]),
   .I0(InputBits[1190]),
   .I1(InputBits[1508]),
   .I2(InputBits[153]),
   .I3(InputBits[665]),
   .I4(InputBits[356]),
   .I5(InputBits[1301])
);
LUT6 #(
   .INIT(64'b1111111011110101000000001101010011110001011001000100111110001100)  
) LUT6_901 (
   .O(gates[77]),
   .I0(InputBits[973]),
   .I1(InputBits[36]),
   .I2(InputBits[122]),
   .I3(InputBits[1181]),
   .I4(InputBits[479]),
   .I5(InputBits[644])
);
LUT6 #(
   .INIT(64'b0010110111110011100101011001101110110001010101000110110110000100)  
) LUT6_902 (
   .O(gates[683]),
   .I0(InputBits[845]),
   .I1(InputBits[703]),
   .I2(InputBits[619]),
   .I3(InputBits[474]),
   .I4(InputBits[794]),
   .I5(InputBits[1447])
);
LUT6 #(
   .INIT(64'b0011010001010000100001111101111000101110101110001000011101001010)  
) LUT6_903 (
   .O(gates[541]),
   .I0(InputBits[1197]),
   .I1(InputBits[1168]),
   .I2(InputBits[1558]),
   .I3(InputBits[438]),
   .I4(InputBits[338]),
   .I5(InputBits[91])
);
LUT6 #(
   .INIT(64'b0000000100000001011100011100110111000001100110000000010001110011)  
) LUT6_904 (
   .O(gates[1215]),
   .I0(InputBits[788]),
   .I1(InputBits[1455]),
   .I2(InputBits[963]),
   .I3(InputBits[1489]),
   .I4(InputBits[553]),
   .I5(InputBits[821])
);
LUT6 #(
   .INIT(64'b1010101010101111001000001110111010111110010001010001101101010001)  
) LUT6_905 (
   .O(gates[64]),
   .I0(InputBits[428]),
   .I1(InputBits[1545]),
   .I2(InputBits[468]),
   .I3(InputBits[422]),
   .I4(InputBits[199]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b0000110011011110010110101101110000001001111101011000110111101101)  
) LUT6_906 (
   .O(gates[1473]),
   .I0(InputBits[270]),
   .I1(InputBits[114]),
   .I2(InputBits[397]),
   .I3(InputBits[538]),
   .I4(InputBits[1475]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0010010011110100101001001111000000101001110001010101000110101010)  
) LUT6_907 (
   .O(gates[765]),
   .I0(InputBits[1298]),
   .I1(InputBits[1040]),
   .I2(InputBits[59]),
   .I3(InputBits[663]),
   .I4(InputBits[761]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b1000000110011110110100001100010111100011000001101100010001001011)  
) LUT6_908 (
   .O(gates[881]),
   .I0(InputBits[404]),
   .I1(InputBits[520]),
   .I2(InputBits[426]),
   .I3(InputBits[1696]),
   .I4(InputBits[990]),
   .I5(InputBits[1206])
);
LUT6 #(
   .INIT(64'b0010110010001100101000101000011010001001000110010111000010110110)  
) LUT6_909 (
   .O(gates[312]),
   .I0(InputBits[1441]),
   .I1(InputBits[319]),
   .I2(InputBits[1650]),
   .I3(InputBits[526]),
   .I4(InputBits[248]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b1011111100001000011000010111100010001110011110100110011111010000)  
) LUT6_910 (
   .O(gates[897]),
   .I0(InputBits[967]),
   .I1(InputBits[753]),
   .I2(InputBits[12]),
   .I3(InputBits[896]),
   .I4(InputBits[221]),
   .I5(InputBits[1010])
);
LUT6 #(
   .INIT(64'b1001110111100011100001000111101010110001000011000011101100111001)  
) LUT6_911 (
   .O(gates[45]),
   .I0(InputBits[603]),
   .I1(InputBits[1492]),
   .I2(InputBits[1021]),
   .I3(InputBits[637]),
   .I4(InputBits[1112]),
   .I5(InputBits[807])
);
LUT6 #(
   .INIT(64'b1100111010101101011011111111111010111100001001011010000010010000)  
) LUT6_912 (
   .O(gates[405]),
   .I0(InputBits[860]),
   .I1(InputBits[1028]),
   .I2(InputBits[1241]),
   .I3(InputBits[1034]),
   .I4(InputBits[440]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b0110000011111011000101000101100110010111011001110001001010000111)  
) LUT6_913 (
   .O(gates[507]),
   .I0(InputBits[1259]),
   .I1(InputBits[801]),
   .I2(InputBits[101]),
   .I3(InputBits[279]),
   .I4(InputBits[587]),
   .I5(InputBits[655])
);
LUT6 #(
   .INIT(64'b0110001100010101011011011001011010001101010100001011100011100010)  
) LUT6_914 (
   .O(gates[237]),
   .I0(InputBits[109]),
   .I1(InputBits[1656]),
   .I2(InputBits[1103]),
   .I3(InputBits[1178]),
   .I4(InputBits[912]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b0100101110111110010000010111011001111001111000110000001111000011)  
) LUT6_915 (
   .O(gates[1002]),
   .I0(InputBits[1225]),
   .I1(InputBits[771]),
   .I2(InputBits[626]),
   .I3(InputBits[389]),
   .I4(InputBits[1534]),
   .I5(InputBits[674])
);
LUT6 #(
   .INIT(64'b0110110101000110111001001001101010000110111001001111101100011101)  
) LUT6_916 (
   .O(gates[1173]),
   .I0(InputBits[27]),
   .I1(InputBits[881]),
   .I2(InputBits[1287]),
   .I3(InputBits[44]),
   .I4(InputBits[1458]),
   .I5(InputBits[751])
);
LUT6 #(
   .INIT(64'b0010001110010110011111100011010111100000101110100101010110001100)  
) LUT6_917 (
   .O(gates[370]),
   .I0(InputBits[1345]),
   .I1(InputBits[1035]),
   .I2(InputBits[828]),
   .I3(InputBits[1559]),
   .I4(InputBits[1097]),
   .I5(InputBits[782])
);
LUT6 #(
   .INIT(64'b1000101110011111100101101100011001011011100100001101001010011001)  
) LUT6_918 (
   .O(gates[309]),
   .I0(InputBits[728]),
   .I1(InputBits[1048]),
   .I2(InputBits[688]),
   .I3(InputBits[1131]),
   .I4(InputBits[852]),
   .I5(InputBits[1327])
);
LUT6 #(
   .INIT(64'b0011001001111110110000111000100011011111001111010000011000100010)  
) LUT6_919 (
   .O(gates[567]),
   .I0(InputBits[1679]),
   .I1(InputBits[107]),
   .I2(InputBits[544]),
   .I3(InputBits[1140]),
   .I4(InputBits[921]),
   .I5(InputBits[1433])
);
LUT6 #(
   .INIT(64'b0111101010111101001010110101000110001011110000111011111100101000)  
) LUT6_920 (
   .O(gates[416]),
   .I0(InputBits[32]),
   .I1(InputBits[366]),
   .I2(InputBits[4]),
   .I3(InputBits[1311]),
   .I4(InputBits[1662]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1110110000001010101010010010100101000110110100010000110010000000)  
) LUT6_921 (
   .O(gates[380]),
   .I0(InputBits[146]),
   .I1(InputBits[305]),
   .I2(InputBits[561]),
   .I3(InputBits[888]),
   .I4(InputBits[695]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b1000110001100001000101110111000001100000011000111110101111010111)  
) LUT6_922 (
   .O(gates[100]),
   .I0(InputBits[346]),
   .I1(InputBits[382]),
   .I2(InputBits[675]),
   .I3(InputBits[330]),
   .I4(InputBits[1210]),
   .I5(InputBits[1350])
);
LUT6 #(
   .INIT(64'b0110111111011100011011011000001111000101001011110001110110000001)  
) LUT6_923 (
   .O(gates[914]),
   .I0(InputBits[262]),
   .I1(InputBits[744]),
   .I2(InputBits[1265]),
   .I3(InputBits[1053]),
   .I4(InputBits[1059]),
   .I5(InputBits[1152])
);
LUT6 #(
   .INIT(64'b1000100100100000010000010000110010111010101101111101100100111000)  
) LUT6_924 (
   .O(gates[300]),
   .I0(InputBits[1262]),
   .I1(InputBits[1499]),
   .I2(InputBits[1068]),
   .I3(InputBits[694]),
   .I4(InputBits[302]),
   .I5(InputBits[868])
);
LUT6 #(
   .INIT(64'b1001111100011000100111111000101101000110000001101110101110000010)  
) LUT6_925 (
   .O(gates[1279]),
   .I0(InputBits[50]),
   .I1(InputBits[352]),
   .I2(InputBits[876]),
   .I3(InputBits[1615]),
   .I4(InputBits[390]),
   .I5(InputBits[1605])
);
LUT6 #(
   .INIT(64'b0000100101000111010111110111110010001100011101101001101011101001)  
) LUT6_926 (
   .O(gates[965]),
   .I0(InputBits[1565]),
   .I1(InputBits[1724]),
   .I2(InputBits[766]),
   .I3(InputBits[433]),
   .I4(InputBits[1580]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b1111111100100101110001101110110001011001110100100010100100110101)  
) LUT6_927 (
   .O(gates[1258]),
   .I0(InputBits[1527]),
   .I1(InputBits[1465]),
   .I2(InputBits[721]),
   .I3(InputBits[1707]),
   .I4(InputBits[19]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b1001001111111011010100000010000000000111100011011100001111101010)  
) LUT6_928 (
   .O(gates[1439]),
   .I0(InputBits[1219]),
   .I1(InputBits[1479]),
   .I2(InputBits[1208]),
   .I3(InputBits[216]),
   .I4(InputBits[1416]),
   .I5(InputBits[1434])
);
LUT6 #(
   .INIT(64'b0101011100100011001000001101000100010110000000001001001111011011)  
) LUT6_929 (
   .O(gates[824]),
   .I0(InputBits[1336]),
   .I1(InputBits[854]),
   .I2(InputBits[1278]),
   .I3(InputBits[169]),
   .I4(InputBits[1089]),
   .I5(InputBits[593])
);
LUT6 #(
   .INIT(64'b1011001011011110101010110100001000110100111100110111010111000110)  
) LUT6_930 (
   .O(gates[286]),
   .I0(InputBits[210]),
   .I1(InputBits[1408]),
   .I2(InputBits[1600]),
   .I3(InputBits[1389]),
   .I4(InputBits[1404]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1010101110011010111111110011111101010101100101110100100010111011)  
) LUT6_931 (
   .O(gates[1395]),
   .I0(InputBits[1589]),
   .I1(InputBits[1095]),
   .I2(InputBits[288]),
   .I3(InputBits[1725]),
   .I4(InputBits[1370]),
   .I5(InputBits[1435])
);
LUT6 #(
   .INIT(64'b1000011000110010111011111001000101111010100011110000010001100011)  
) LUT6_932 (
   .O(gates[120]),
   .I0(InputBits[1071]),
   .I1(InputBits[358]),
   .I2(InputBits[684]),
   .I3(InputBits[1474]),
   .I4(InputBits[1157]),
   .I5(InputBits[837])
);
LUT6 #(
   .INIT(64'b1011001001010111110100111101011001010011001000101111111010000101)  
) LUT6_933 (
   .O(gates[1075]),
   .I0(InputBits[7]),
   .I1(InputBits[324]),
   .I2(InputBits[269]),
   .I3(InputBits[645]),
   .I4(InputBits[726]),
   .I5(InputBits[1362])
);
LUT6 #(
   .INIT(64'b1110111000111000111010011111011111011110111001001111101111010100)  
) LUT6_934 (
   .O(gates[800]),
   .I0(InputBits[2]),
   .I1(InputBits[314]),
   .I2(InputBits[1635]),
   .I3(InputBits[1502]),
   .I4(InputBits[787]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b1010000001101011100010100001110001110001101111110111011010001100)  
) LUT6_935 (
   .O(gates[1148]),
   .I0(InputBits[749]),
   .I1(InputBits[1321]),
   .I2(InputBits[786]),
   .I3(InputBits[580]),
   .I4(InputBits[1249]),
   .I5(InputBits[1292])
);
LUT6 #(
   .INIT(64'b1100001001011110101001001000100001100010111100000011100010001011)  
) LUT6_936 (
   .O(gates[392]),
   .I0(InputBits[1678]),
   .I1(InputBits[1460]),
   .I2(InputBits[365]),
   .I3(InputBits[276]),
   .I4(InputBits[910]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0101111101000111100010001010100000110011010111001011111110100111)  
) LUT6_937 (
   .O(gates[254]),
   .I0(InputBits[1310]),
   .I1(InputBits[143]),
   .I2(InputBits[1227]),
   .I3(InputBits[1437]),
   .I4(InputBits[482]),
   .I5(InputBits[1084])
);
LUT6 #(
   .INIT(64'b1111100001101011100100001001010111010100100101000011011001010110)  
) LUT6_938 (
   .O(gates[1321]),
   .I0(InputBits[900]),
   .I1(InputBits[843]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[1087]),
   .I5(InputBits[799])
);
LUT6 #(
   .INIT(64'b1111000100001010000101000011011001001001001100101000010101100110)  
) LUT6_939 (
   .O(gates[1365]),
   .I0(InputBits[70]),
   .I1(InputBits[281]),
   .I2(InputBits[1431]),
   .I3(InputBits[847]),
   .I4(InputBits[1176]),
   .I5(InputBits[1374])
);
LUT6 #(
   .INIT(64'b0000001100011001001000100011000101001101110010101101111100011110)  
) LUT6_940 (
   .O(gates[1407]),
   .I0(InputBits[740]),
   .I1(InputBits[898]),
   .I2(InputBits[286]),
   .I3(InputBits[327]),
   .I4(InputBits[1272]),
   .I5(InputBits[1183])
);
LUT6 #(
   .INIT(64'b0100011101010100110101100110010011110110000111000010110110011011)  
) LUT6_941 (
   .O(gates[496]),
   .I0(InputBits[1466]),
   .I1(InputBits[1031]),
   .I2(InputBits[1203]),
   .I3(InputBits[1610]),
   .I4(InputBits[978]),
   .I5(InputBits[1215])
);
LUT6 #(
   .INIT(64'b1001110101010110110100000010001011110100011100010010000000001000)  
) LUT6_942 (
   .O(gates[605]),
   .I0(InputBits[1086]),
   .I1(InputBits[1115]),
   .I2(InputBits[1532]),
   .I3(InputBits[1452]),
   .I4(InputBits[29]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b1101000101011010011111110101100101011010011010010011111111011001)  
) LUT6_943 (
   .O(gates[607]),
   .I0(InputBits[22]),
   .I1(InputBits[601]),
   .I2(InputBits[17]),
   .I3(InputBits[1296]),
   .I4(InputBits[1417]),
   .I5(InputBits[1574])
);
LUT6 #(
   .INIT(64'b1111011010010110110111100011101110011100111000101000101001000010)  
) LUT6_944 (
   .O(gates[813]),
   .I0(InputBits[595]),
   .I1(InputBits[451]),
   .I2(InputBits[690]),
   .I3(InputBits[1623]),
   .I4(InputBits[1280]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b1010100111101001001000110000111010100001011001010100010001100001)  
) LUT6_945 (
   .O(gates[42]),
   .I0(InputBits[1314]),
   .I1(InputBits[575]),
   .I2(InputBits[353]),
   .I3(InputBits[170]),
   .I4(InputBits[34]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b0000111001001000011001011101011001000011101111011011000011110110)  
) LUT6_946 (
   .O(gates[759]),
   .I0(InputBits[995]),
   .I1(InputBits[1237]),
   .I2(InputBits[824]),
   .I3(InputBits[1128]),
   .I4(InputBits[1688]),
   .I5(InputBits[1448])
);
LUT6 #(
   .INIT(64'b1111000010100010111100111001110101111111000001001011011100010111)  
) LUT6_947 (
   .O(gates[644]),
   .I0(InputBits[1064]),
   .I1(InputBits[464]),
   .I2(InputBits[115]),
   .I3(InputBits[455]),
   .I4(InputBits[1110]),
   .I5(InputBits[1279])
);
LUT6 #(
   .INIT(64'b0110100100011011000000000000111001111111111001111000111110101100)  
) LUT6_948 (
   .O(gates[851]),
   .I0(InputBits[57]),
   .I1(InputBits[913]),
   .I2(InputBits[1727]),
   .I3(InputBits[193]),
   .I4(InputBits[572]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0011111111111110001011011011001100110001101001011100101010111000)  
) LUT6_949 (
   .O(gates[399]),
   .I0(InputBits[628]),
   .I1(InputBits[667]),
   .I2(InputBits[15]),
   .I3(InputBits[1118]),
   .I4(InputBits[345]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b0111101010001010011010000000000011100001010100100011000000000010)  
) LUT6_950 (
   .O(gates[1228]),
   .I0(InputBits[1023]),
   .I1(InputBits[116]),
   .I2(InputBits[486]),
   .I3(InputBits[507]),
   .I4(InputBits[1338]),
   .I5(InputBits[1596])
);
LUT6 #(
   .INIT(64'b0011101011011001010001010100111010011111000100111101001110010111)  
) LUT6_951 (
   .O(gates[235]),
   .I0(InputBits[1506]),
   .I1(InputBits[1246]),
   .I2(InputBits[8]),
   .I3(InputBits[1536]),
   .I4(InputBits[611]),
   .I5(InputBits[1331])
);
LUT6 #(
   .INIT(64'b1111000100011100010111110000000011011001110010110101100100000111)  
) LUT6_952 (
   .O(gates[1073]),
   .I0(InputBits[988]),
   .I1(InputBits[245]),
   .I2(InputBits[1266]),
   .I3(InputBits[546]),
   .I4(InputBits[162]),
   .I5(InputBits[1507])
);
LUT6 #(
   .INIT(64'b1000001011010010011010101000101101011101111110110101010000100011)  
) LUT6_953 (
   .O(gates[694]),
   .I0(InputBits[1002]),
   .I1(InputBits[1160]),
   .I2(InputBits[550]),
   .I3(InputBits[79]),
   .I4(InputBits[1139]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0000100101001000110110000001000010111010001011011101101110101011)  
) LUT6_954 (
   .O(gates[436]),
   .I0(InputBits[293]),
   .I1(InputBits[621]),
   .I2(InputBits[1236]),
   .I3(InputBits[1159]),
   .I4(InputBits[1102]),
   .I5(InputBits[755])
);
LUT6 #(
   .INIT(64'b0011001000111010110001100101010001010101111100001001100110011101)  
) LUT6_955 (
   .O(gates[1342]),
   .I0(InputBits[312]),
   .I1(InputBits[940]),
   .I2(InputBits[931]),
   .I3(InputBits[1497]),
   .I4(InputBits[767]),
   .I5(InputBits[883])
);
LUT6 #(
   .INIT(64'b1010001000110000011110100011011000011001010010101011111010101010)  
) LUT6_956 (
   .O(gates[94]),
   .I0(InputBits[762]),
   .I1(InputBits[1722]),
   .I2(InputBits[68]),
   .I3(InputBits[1691]),
   .I4(InputBits[950]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b1011111111011110101010000111000110110010000100111001100011100011)  
) LUT6_957 (
   .O(gates[213]),
   .I0(InputBits[1381]),
   .I1(InputBits[654]),
   .I2(InputBits[371]),
   .I3(InputBits[469]),
   .I4(InputBits[819]),
   .I5(InputBits[970])
);
LUT6 #(
   .INIT(64'b1011100100101011001001010010000000100110001011110110101111011100)  
) LUT6_958 (
   .O(gates[816]),
   .I0(InputBits[495]),
   .I1(InputBits[139]),
   .I2(InputBits[343]),
   .I3(InputBits[764]),
   .I4(InputBits[1186]),
   .I5(InputBits[1073])
);
LUT6 #(
   .INIT(64'b1100101100111001101011100100011101010110110111000011110110011000)  
) LUT6_959 (
   .O(gates[1103]),
   .I0(InputBits[915]),
   .I1(InputBits[232]),
   .I2(InputBits[1217]),
   .I3(InputBits[196]),
   .I4(InputBits[696]),
   .I5(InputBits[582])
);
LUT6 #(
   .INIT(64'b1011101000111101101111101111011000010000110000101010011001010100)  
) LUT6_960 (
   .O(gates[1450]),
   .I0(InputBits[1628]),
   .I1(InputBits[1260]),
   .I2(InputBits[1524]),
   .I3(InputBits[1239]),
   .I4(InputBits[566]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0101110111000111110110000000111011011011000010010101011100101100)  
) LUT6_961 (
   .O(gates[568]),
   .I0(InputBits[1515]),
   .I1(InputBits[1153]),
   .I2(InputBits[1007]),
   .I3(InputBits[95]),
   .I4(InputBits[1196]),
   .I5(InputBits[1539])
);
LUT6 #(
   .INIT(64'b0111110111101100010001001000000111000110010111000110101100001001)  
) LUT6_962 (
   .O(gates[296]),
   .I0(InputBits[1234]),
   .I1(InputBits[519]),
   .I2(InputBits[984]),
   .I3(InputBits[1295]),
   .I4(InputBits[992]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0000100110110101001011111001111000001100111110010010100000011110)  
) LUT6_963 (
   .O(gates[265]),
   .I0(InputBits[1224]),
   .I1(InputBits[1693]),
   .I2(InputBits[1364]),
   .I3(InputBits[1398]),
   .I4(InputBits[584]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b0011101000101001000100100011001111011001001010010100000011101001)  
) LUT6_964 (
   .O(gates[1062]),
   .I0(InputBits[228]),
   .I1(InputBits[373]),
   .I2(InputBits[201]),
   .I3(InputBits[700]),
   .I4(InputBits[81]),
   .I5(InputBits[936])
);
LUT6 #(
   .INIT(64'b0010010011110001000101111101000111111010011111100000100111000011)  
) LUT6_965 (
   .O(gates[1129]),
   .I0(InputBits[504]),
   .I1(InputBits[272]),
   .I2(InputBits[959]),
   .I3(InputBits[811]),
   .I4(InputBits[946]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b1101111101000010110111000010100000010110000000111110100111001010)  
) LUT6_966 (
   .O(gates[791]),
   .I0(InputBits[1550]),
   .I1(InputBits[441]),
   .I2(InputBits[1356]),
   .I3(InputBits[715]),
   .I4(InputBits[220]),
   .I5(InputBits[863])
);
LUT6 #(
   .INIT(64'b0111101111111010100101111101001001011000000100111101001000100000)  
) LUT6_967 (
   .O(gates[171]),
   .I0(InputBits[1577]),
   .I1(InputBits[779]),
   .I2(InputBits[975]),
   .I3(InputBits[510]),
   .I4(InputBits[1401]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b1011100011111100000011100011000111111111001000011111001111001100)  
) LUT6_968 (
   .O(gates[1143]),
   .I0(InputBits[1698]),
   .I1(InputBits[834]),
   .I2(InputBits[1009]),
   .I3(InputBits[1690]),
   .I4(InputBits[827]),
   .I5(InputBits[1391])
);
LUT6 #(
   .INIT(64'b0101101100001001100000110010010000111010010111111010001101100010)  
) LUT6_969 (
   .O(gates[1355]),
   .I0(InputBits[1093]),
   .I1(InputBits[1080]),
   .I2(InputBits[175]),
   .I3(InputBits[722]),
   .I4(InputBits[798]),
   .I5(InputBits[296])
);
LUT6 #(
   .INIT(64'b0000001011111010100011001100000100111011001011010001101001110111)  
) LUT6_970 (
   .O(gates[386]),
   .I0(InputBits[1643]),
   .I1(InputBits[1660]),
   .I2(InputBits[1075]),
   .I3(InputBits[604]),
   .I4(InputBits[1504]),
   .I5(InputBits[818])
);
LUT6 #(
   .INIT(64'b0001010101000110010011100001011110101100011111100010100100011110)  
) LUT6_971 (
   .O(gates[916]),
   .I0(InputBits[708]),
   .I1(InputBits[100]),
   .I2(InputBits[388]),
   .I3(InputBits[1708]),
   .I4(InputBits[1318]),
   .I5(InputBits[236])
);
LUT6 #(
   .INIT(64'b1000000110010010110000101010100111010111010001011111100001111111)  
) LUT6_972 (
   .O(gates[1457]),
   .I0(InputBits[87]),
   .I1(InputBits[94]),
   .I2(InputBits[671]),
   .I3(InputBits[1323]),
   .I4(InputBits[625]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b1111100001010101001000110000110101110101010010000000111000000010)  
) LUT6_973 (
   .O(gates[445]),
   .I0(InputBits[1214]),
   .I1(InputBits[1193]),
   .I2(InputBits[243]),
   .I3(InputBits[980]),
   .I4(InputBits[77]),
   .I5(InputBits[857])
);
LUT6 #(
   .INIT(64'b0011110011100001101100100111000100001011010010011010010111110001)  
) LUT6_974 (
   .O(gates[200]),
   .I0(InputBits[132]),
   .I1(InputBits[597]),
   .I2(InputBits[724]),
   .I3(InputBits[278]),
   .I4(InputBits[1587]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0100000010111010000111000010000011001000000001111101011110100101)  
) LUT6_975 (
   .O(gates[1339]),
   .I0(InputBits[1251]),
   .I1(InputBits[1564]),
   .I2(InputBits[1307]),
   .I3(InputBits[9]),
   .I4(InputBits[234]),
   .I5(InputBits[1477])
);
LUT6 #(
   .INIT(64'b0101011111101111001100110101110000000111101011001010101111011110)  
) LUT6_976 (
   .O(gates[1261]),
   .I0(InputBits[685]),
   .I1(InputBits[462]),
   .I2(InputBits[1108]),
   .I3(InputBits[1637]),
   .I4(InputBits[521]),
   .I5(InputBits[1468])
);
LUT6 #(
   .INIT(64'b0110001011001001000100000010110111000000001011101000010001010000)  
) LUT6_977 (
   .O(gates[1352]),
   .I0(InputBits[1329]),
   .I1(InputBits[1106]),
   .I2(InputBits[283]),
   .I3(InputBits[218]),
   .I4(InputBits[1611]),
   .I5(InputBits[1018])
);
LUT6 #(
   .INIT(64'b1111111110100101000111000000000111111010000010010100000111011010)  
) LUT6_978 (
   .O(gates[329]),
   .I0(InputBits[1429]),
   .I1(InputBits[1522]),
   .I2(InputBits[1379]),
   .I3(InputBits[1305]),
   .I4(InputBits[102]),
   .I5(InputBits[1586])
);
LUT6 #(
   .INIT(64'b0110000011010011111000011001000101110101011010001010001101000011)  
) LUT6_979 (
   .O(gates[525]),
   .I0(InputBits[835]),
   .I1(InputBits[1454]),
   .I2(InputBits[630]),
   .I3(InputBits[1162]),
   .I4(InputBits[1025]),
   .I5(InputBits[1572])
);
LUT6 #(
   .INIT(64'b0111010111010100011101000011100011000011101101001111001111100101)  
) LUT6_980 (
   .O(gates[27]),
   .I0(InputBits[796]),
   .I1(InputBits[564]),
   .I2(InputBits[198]),
   .I3(InputBits[1632]),
   .I4(InputBits[570]),
   .I5(InputBits[1133])
);
LUT6 #(
   .INIT(64'b0100011101000101011011010000110000001010111000010011111101010011)  
) LUT6_981 (
   .O(gates[787]),
   .I0(InputBits[292]),
   .I1(InputBits[998]),
   .I2(InputBits[242]),
   .I3(InputBits[1424]),
   .I4(InputBits[359]),
   .I5(InputBits[1715])
);
LUT6 #(
   .INIT(64'b1100111001101100101011110101100101100110101001000000011111111011)  
) LUT6_982 (
   .O(gates[161]),
   .I0(InputBits[891]),
   .I1(InputBits[1484]),
   .I2(InputBits[1014]),
   .I3(InputBits[1406]),
   .I4(InputBits[364]),
   .I5(InputBits[1201])
);
LUT6 #(
   .INIT(64'b1000011110101001100100111100110111100110110001110101111100110111)  
) LUT6_983 (
   .O(gates[582]),
   .I0(InputBits[150]),
   .I1(InputBits[383]),
   .I2(InputBits[1445]),
   .I3(InputBits[540]),
   .I4(InputBits[1672]),
   .I5(InputBits[1046])
);
LUT6 #(
   .INIT(64'b0010101101100100101111001111110000010111001111000010001100101101)  
) LUT6_984 (
   .O(gates[109]),
   .I0(InputBits[1044]),
   .I1(InputBits[1405]),
   .I2(InputBits[1552]),
   .I3(InputBits[1423]),
   .I4(InputBits[31]),
   .I5(InputBits[1016])
);
LUT6 #(
   .INIT(64'b0010010110000111011000100100110100001101100100001010101000011010)  
) LUT6_985 (
   .O(gates[1310]),
   .I0(InputBits[431]),
   .I1(InputBits[1302]),
   .I2(InputBits[1051]),
   .I3(InputBits[367]),
   .I4(InputBits[1493]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b0111100001100110100011000111010110000000001111000110010010101000)  
) LUT6_986 (
   .O(gates[557]),
   .I0(InputBits[258]),
   .I1(InputBits[1393]),
   .I2(InputBits[842]),
   .I3(InputBits[505]),
   .I4(InputBits[1074]),
   .I5(InputBits[113])
);
LUT6 #(
   .INIT(64'b1111111011101001110001110001001111100100010100010000000110110000)  
) LUT6_987 (
   .O(gates[718]),
   .I0(InputBits[160]),
   .I1(InputBits[742]),
   .I2(InputBits[608]),
   .I3(InputBits[659]),
   .I4(InputBits[58]),
   .I5(InputBits[1349])
);
LUT6 #(
   .INIT(64'b0010110000111101000111001000001010110100010001101111111100111110)  
) LUT6_988 (
   .O(gates[1507]),
   .I0(InputBits[548]),
   .I1(InputBits[1394]),
   .I2(InputBits[791]),
   .I3(InputBits[155]),
   .I4(InputBits[640]),
   .I5(InputBits[669])
);
LUT6 #(
   .INIT(64'b1110100010100101001110001011110101000101110111100010010000111100)  
) LUT6_989 (
   .O(gates[1239]),
   .I0(InputBits[557]),
   .I1(InputBits[866]),
   .I2(InputBits[350]),
   .I3(InputBits[666]),
   .I4(InputBits[1282]),
   .I5(InputBits[1000])
);
LUT6 #(
   .INIT(64'b1000111100000001100001000110001111010111011101100101111111000100)  
) LUT6_990 (
   .O(gates[441]),
   .I0(InputBits[1648]),
   .I1(InputBits[1427]),
   .I2(InputBits[20]),
   .I3(InputBits[257]),
   .I4(InputBits[1681]),
   .I5(InputBits[873])
);
LUT6 #(
   .INIT(64'b1000100100101111000001111010100010010000010111010101000101000101)  
) LUT6_991 (
   .O(gates[868]),
   .I0(InputBits[386]),
   .I1(InputBits[214]),
   .I2(InputBits[1271]),
   .I3(InputBits[652]),
   .I4(InputBits[920]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b1010000110111101101110000111001111101011111111111110010111100100)  
) LUT6_992 (
   .O(gates[672]),
   .I0(InputBits[917]),
   .I1(InputBits[118]),
   .I2(InputBits[577]),
   .I3(InputBits[977]),
   .I4(InputBits[1626]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0001001001011010001011010011101110101110000110111100001100100001)  
) LUT6_993 (
   .O(gates[769]),
   .I0(InputBits[1057]),
   .I1(InputBits[166]),
   .I2(InputBits[942]),
   .I3(InputBits[624]),
   .I4(InputBits[617]),
   .I5(InputBits[476])
);
LUT6 #(
   .INIT(64'b0010010100001011010110101100010110101100010111011000101101100100)  
) LUT6_994 (
   .O(gates[1140]),
   .I0(InputBits[1495]),
   .I1(InputBits[717]),
   .I2(InputBits[334]),
   .I3(InputBits[1137]),
   .I4(InputBits[698]),
   .I5(InputBits[1091])
);
LUT6 #(
   .INIT(64'b1111001000010110100010110000010000011110011110001100100011100111)  
) LUT6_995 (
   .O(gates[1181]),
   .I0(InputBits[878]),
   .I1(InputBits[41]),
   .I2(InputBits[1232]),
   .I3(InputBits[250]),
   .I4(InputBits[1671]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b1011000100001001001000011000100000100010000110100101011110010100)  
) LUT6_996 (
   .O(gates[275]),
   .I0(InputBits[172]),
   .I1(InputBits[1367]),
   .I2(InputBits[542]),
   .I3(InputBits[1142]),
   .I4(InputBits[1269]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b0101010110110100111111010110001000110110001010111100001001000100)  
) LUT6_997 (
   .O(gates[983]),
   .I0(InputBits[1184]),
   .I1(InputBits[181]),
   .I2(InputBits[14]),
   .I3(InputBits[623]),
   .I4(InputBits[460]),
   .I5(InputBits[1354])
);
LUT6 #(
   .INIT(64'b0010000001101110101101001111001101010100100001001111001110001010)  
) LUT6_998 (
   .O(gates[803]),
   .I0(InputBits[1653]),
   .I1(InputBits[987]),
   .I2(InputBits[423]),
   .I3(InputBits[568]),
   .I4(InputBits[809]),
   .I5(InputBits[734])
);
LUT6 #(
   .INIT(64'b1101011001000101100001100100001000100011011010101111001011100101)  
) LUT6_999 (
   .O(gates[197]),
   .I0(InputBits[1005]),
   .I1(InputBits[85]),
   .I2(InputBits[1728]),
   .I3(InputBits[757]),
   .I4(InputBits[1154]),
   .I5(InputBits[1512])
);
LUT6 #(
   .INIT(64'b0010111000100000110011110101110101000001111111101111000100010111)  
) LUT6_1000 (
   .O(gates[853]),
   .I0(InputBits[1541]),
   .I1(InputBits[1120]),
   .I2(InputBits[1147]),
   .I3(InputBits[1175]),
   .I4(InputBits[1700]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0011010010101011000100001110001001111111111001001101100100011010)  
) LUT6_1001 (
   .O(gates[751]),
   .I0(InputBits[1038]),
   .I1(InputBits[1641]),
   .I2(InputBits[1575]),
   .I3(InputBits[466]),
   .I4(InputBits[805]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1110101111100101011110111000010000001001001110111110110110100111)  
) LUT6_1002 (
   .O(gates[60]),
   .I0(InputBits[1365]),
   .I1(InputBits[141]),
   .I2(InputBits[1613]),
   .I3(InputBits[848]),
   .I4(InputBits[483]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b1001100001011010111000101001110001001011101100100100100111010111)  
) LUT6_1003 (
   .O(gates[1500]),
   .I0(InputBits[1568]),
   .I1(InputBits[706]),
   .I2(InputBits[493]),
   .I3(InputBits[1555]),
   .I4(InputBits[536]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b0100111111101101011001111001001000100100011000101011110000110100)  
) LUT6_1004 (
   .O(gates[1245]),
   .I0(InputBits[777]),
   .I1(InputBits[416]),
   .I2(InputBits[1375]),
   .I3(InputBits[803]),
   .I4(InputBits[943]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b0100111100001010001100100100100110001110100101000000110111001011)  
) LUT6_1005 (
   .O(gates[1400]),
   .I0(InputBits[189]),
   .I1(InputBits[692]),
   .I2(InputBits[1619]),
   .I3(InputBits[1562]),
   .I4(InputBits[1312]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1001001001110111011111000011000000101001010101011011110100111010)  
) LUT6_1006 (
   .O(gates[691]),
   .I0(InputBits[1316]),
   .I1(InputBits[308]),
   .I2(InputBits[1720]),
   .I3(InputBits[1358]),
   .I4(InputBits[908]),
   .I5(InputBits[745])
);
LUT6 #(
   .INIT(64'b0100101010010010110110000000110101101011110110111000111100101100)  
) LUT6_1007 (
   .O(gates[1067]),
   .I0(InputBits[925]),
   .I1(InputBits[938]),
   .I2(InputBits[92]),
   .I3(InputBits[341]),
   .I4(InputBits[1340]),
   .I5(InputBits[825])
);
LUT6 #(
   .INIT(64'b1011001010110010010110100011001011101010011011011010111010100111)  
) LUT6_1008 (
   .O(gates[1388]),
   .I0(InputBits[813]),
   .I1(InputBits[131]),
   .I2(InputBits[400]),
   .I3(InputBits[1710]),
   .I4(InputBits[1222]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0010011111010011011111100111100010101000100111000010000110000100)  
) LUT6_1009 (
   .O(gates[346]),
   .I0(InputBits[1229]),
   .I1(InputBits[119]),
   .I2(InputBits[1639]),
   .I3(InputBits[679]),
   .I4(InputBits[104]),
   .I5(InputBits[1191])
);
LUT6 #(
   .INIT(64'b0010111101111100110001001100011011101000001000101001011111101110)  
) LUT6_1010 (
   .O(gates[911]),
   .I0(InputBits[240]),
   .I1(InputBits[1482]),
   .I2(InputBits[673]),
   .I3(InputBits[515]),
   .I4(InputBits[1245]),
   .I5(InputBits[618])
);
LUT6 #(
   .INIT(64'b0000011101101101111011100011100110110010100101001010011111010101)  
) LUT6_1011 (
   .O(gates[1295]),
   .I0(InputBits[213]),
   .I1(InputBits[1194]),
   .I2(InputBits[968]),
   .I3(InputBits[1718]),
   .I4(InputBits[840]),
   .I5(InputBits[810])
);
LUT6 #(
   .INIT(64'b1001010001110011110011001000110101101011000001111101111011100111)  
) LUT6_1012 (
   .O(gates[427]),
   .I0(InputBits[134]),
   .I1(InputBits[306]),
   .I2(InputBits[752]),
   .I3(InputBits[434]),
   .I4(InputBits[1270]),
   .I5(InputBits[1151])
);
LUT6 #(
   .INIT(64'b1101111001111110001101011010101110001001011101011111000010000111)  
) LUT6_1013 (
   .O(gates[1111]),
   .I0(InputBits[606]),
   .I1(InputBits[1342]),
   .I2(InputBits[605]),
   .I3(InputBits[578]),
   .I4(InputBits[99]),
   .I5(InputBits[895])
);
LUT6 #(
   .INIT(64'b1000101111111111000011011110110000000010010000110000110101110110)  
) LUT6_1014 (
   .O(gates[677]),
   .I0(InputBits[1713]),
   .I1(InputBits[1461]),
   .I2(InputBits[315]),
   .I3(InputBits[994]),
   .I4(InputBits[681]),
   .I5(InputBits[1674])
);
LUT6 #(
   .INIT(64'b0000101110000010011111010001010101111010000011110010101101010101)  
) LUT6_1015 (
   .O(gates[907]),
   .I0(InputBits[1291]),
   .I1(InputBits[911]),
   .I2(InputBits[1591]),
   .I3(InputBits[1300]),
   .I4(InputBits[1188]),
   .I5(InputBits[18])
);
LUT6 #(
   .INIT(64'b1001011000100111110000000100101001011001010011101000110110001111)  
) LUT6_1016 (
   .O(gates[82]),
   .I0(InputBits[1721]),
   .I1(InputBits[1453]),
   .I2(InputBits[465]),
   .I3(InputBits[590]),
   .I4(InputBits[1020]),
   .I5(InputBits[444])
);
LUT6 #(
   .INIT(64'b0000011001110110101111001100110000101000001000111110111110100000)  
) LUT6_1017 (
   .O(gates[650]),
   .I0(InputBits[649]),
   .I1(InputBits[1067]),
   .I2(InputBits[1469]),
   .I3(InputBits[1244]),
   .I4(InputBits[237]),
   .I5(InputBits[1335])
);
LUT6 #(
   .INIT(64'b0101000110100110101111110011011011000100110001011110001101001101)  
) LUT6_1018 (
   .O(gates[1154]),
   .I0(InputBits[217]),
   .I1(InputBits[769]),
   .I2(InputBits[662]),
   .I3(InputBits[778]),
   .I4(InputBits[1119]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0111111001001011001001000110011011001101000111011111000100110110)  
) LUT6_1019 (
   .O(gates[590]),
   .I0(InputBits[1601]),
   .I1(InputBits[1173]),
   .I2(InputBits[497]),
   .I3(InputBits[321]),
   .I4(InputBits[1313]),
   .I5(InputBits[1412])
);
LUT6 #(
   .INIT(64'b0101110011001100001010110010111101001010101000111001100110110110)  
) LUT6_1020 (
   .O(gates[1210]),
   .I0(InputBits[204]),
   .I1(InputBits[562]),
   .I2(InputBits[419]),
   .I3(InputBits[477]),
   .I4(InputBits[379]),
   .I5(InputBits[981])
);
LUT6 #(
   .INIT(64'b1000111111100001110000111100001100111001110011100101011100110100)  
) LUT6_1021 (
   .O(gates[895]),
   .I0(InputBits[948]),
   .I1(InputBits[646]),
   .I2(InputBits[361]),
   .I3(InputBits[928]),
   .I4(InputBits[1471]),
   .I5(InputBits[167])
);
LUT6 #(
   .INIT(64'b0110000000000001000001000100010000100000010111110111100001011010)  
) LUT6_1022 (
   .O(gates[69]),
   .I0(InputBits[1252]),
   .I1(InputBits[748]),
   .I2(InputBits[1514]),
   .I3(InputBits[137]),
   .I4(InputBits[1125]),
   .I5(InputBits[704])
);
LUT6 #(
   .INIT(64'b1000100100111010010011011000000001100000101000011111110111111010)  
) LUT6_1023 (
   .O(gates[1157]),
   .I0(InputBits[1122]),
   .I1(InputBits[1402]),
   .I2(InputBits[290]),
   .I3(InputBits[123]),
   .I4(InputBits[1509]),
   .I5(InputBits[657])
);
LUT6 #(
   .INIT(64'b0111110111111011110010010010100111011100100111111000010001101011)  
) LUT6_1024 (
   .O(gates[664]),
   .I0(InputBits[331]),
   .I1(InputBits[1528]),
   .I2(InputBits[266]),
   .I3(InputBits[417]),
   .I4(InputBits[437]),
   .I5(InputBits[1518])
);
LUT6 #(
   .INIT(64'b0111000011010100000110011111111111111001101101100100101011010010)  
) LUT6_1025 (
   .O(gates[1470]),
   .I0(InputBits[923]),
   .I1(InputBits[287]),
   .I2(InputBits[785]),
   .I3(InputBits[588]),
   .I4(InputBits[710]),
   .I5(InputBits[822])
);
LUT6 #(
   .INIT(64'b1011111110001011000101010011110001101011011100110000101110000010)  
) LUT6_1026 (
   .O(gates[224]),
   .I0(InputBits[894]),
   .I1(InputBits[90]),
   .I2(InputBits[574]),
   .I3(InputBits[945]),
   .I4(InputBits[1607]),
   .I5(InputBits[511])
);
LUT6 #(
   .INIT(64'b0010010100011110010001110001010000001011000001011111010001100100)  
) LUT6_1027 (
   .O(gates[617]),
   .I0(InputBits[1665]),
   .I1(InputBits[1283]),
   .I2(InputBits[200]),
   .I3(InputBits[1256]),
   .I4(InputBits[299]),
   .I5(InputBits[1371])
);
LUT6 #(
   .INIT(64'b0100010100111100101000100110100100111110100010000100001000111101)  
) LUT6_1028 (
   .O(gates[79]),
   .I0(InputBits[1124]),
   .I1(InputBits[1344]),
   .I2(InputBits[1386]),
   .I3(InputBits[1490]),
   .I4(InputBits[627]),
   .I5(InputBits[52])
);
LUT6 #(
   .INIT(64'b0111100000000010011001101100110111110111111001011111101001100000)  
) LUT6_1029 (
   .O(gates[1420]),
   .I0(InputBits[84]),
   .I1(InputBits[636]),
   .I2(InputBits[1062]),
   .I3(InputBits[1376]),
   .I4(InputBits[339]),
   .I5(InputBits[63])
);
LUT6 #(
   .INIT(64'b1010010111110101111101111000111011000111011110111101111010010011)  
) LUT6_1030 (
   .O(gates[352]),
   .I0(InputBits[1583]),
   .I1(InputBits[1581]),
   .I2(InputBits[1328]),
   .I3(InputBits[634]),
   .I4(InputBits[732]),
   .I5(InputBits[985])
);
LUT6 #(
   .INIT(64'b0010101110101010101001111100111111011010101011110010001000001110)  
) LUT6_1031 (
   .O(gates[1006]),
   .I0(InputBits[705]),
   .I1(InputBits[1553]),
   .I2(InputBits[729]),
   .I3(InputBits[1440]),
   .I4(InputBits[157]),
   .I5(InputBits[789])
);
LUT6 #(
   .INIT(64'b0111111110100101111100010101011100111110110011000001101000010010)  
) LUT6_1032 (
   .O(gates[126]),
   .I0(InputBits[1198]),
   .I1(InputBits[997]),
   .I2(InputBits[966]),
   .I3(InputBits[73]),
   .I4(InputBits[906]),
   .I5(InputBits[1631])
);
LUT6 #(
   .INIT(64'b0011011011010100010110010111110110000101111001011010110001010001)  
) LUT6_1033 (
   .O(gates[251]),
   .I0(InputBits[1664]),
   .I1(InputBits[880]),
   .I2(InputBits[1029]),
   .I3(InputBits[408]),
   .I4(InputBits[1167]),
   .I5(InputBits[816])
);
LUT6 #(
   .INIT(64'b0100000110110011001000111111011110111010100000100101111110000101)  
) LUT6_1034 (
   .O(gates[1034]),
   .I0(InputBits[179]),
   .I1(InputBits[964]),
   .I2(InputBits[530]),
   .I3(InputBits[1368]),
   .I4(InputBits[1055]),
   .I5(InputBits[178])
);
LUT6 #(
   .INIT(64'b0001001100110000110011111110111111000111110000110000100100010000)  
) LUT6_1035 (
   .O(gates[426]),
   .I0(InputBits[1675]),
   .I1(InputBits[1395]),
   .I2(InputBits[558]),
   .I3(InputBits[1560]),
   .I4(InputBits[1657]),
   .I5(InputBits[598])
);
LUT6 #(
   .INIT(64'b1001100111001101101111110101101110101111011111101111111101110111)  
) LUT6_1036 (
   .O(gates[369]),
   .I0(InputBits[1651]),
   .I1(InputBits[1419]),
   .I2(InputBits[524]),
   .I3(InputBits[850]),
   .I4(InputBits[1013]),
   .I5(InputBits[871])
);
LUT6 #(
   .INIT(64'b0000001001101000000110001000100001100101010100101101101111000110)  
) LUT6_1037 (
   .O(gates[996]),
   .I0(InputBits[677]),
   .I1(InputBits[831]),
   .I2(InputBits[758]),
   .I3(InputBits[1286]),
   .I4(InputBits[1570]),
   .I5(InputBits[877])
);
LUT6 #(
   .INIT(64'b1100110001111010000001011100000111101010110110101110000110101011)  
) LUT6_1038 (
   .O(gates[1533]),
   .I0(InputBits[687]),
   .I1(InputBits[1274]),
   .I2(InputBits[887]),
   .I3(InputBits[699]),
   .I4(InputBits[432]),
   .I5(InputBits[224])
);
LUT6 #(
   .INIT(64'b1001000001111000011000110101011101101111000110000000001111110111)  
) LUT6_1039 (
   .O(gates[1548]),
   .I0(InputBits[1432]),
   .I1(InputBits[13]),
   .I2(InputBits[1026]),
   .I3(InputBits[252]),
   .I4(InputBits[144]),
   .I5(InputBits[1347])
);
LUT6 #(
   .INIT(64'b0111111101101001110000110011001010101101001000001010111101001101)  
) LUT6_1040 (
   .O(gates[1435]),
   .I0(InputBits[459]),
   .I1(InputBits[1047]),
   .I2(InputBits[922]),
   .I3(InputBits[265]),
   .I4(InputBits[1538]),
   .I5(InputBits[953])
);
LUT6 #(
   .INIT(64'b1101010100100001000101010101011000101101101100001101111100011011)  
) LUT6_1041 (
   .O(gates[651]),
   .I0(InputBits[741]),
   .I1(InputBits[736]),
   .I2(InputBits[632]),
   .I3(InputBits[376]),
   .I4(InputBits[1036]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1001011010101010011101001010000100010100011001010010001011101100)  
) LUT6_1042 (
   .O(gates[279]),
   .I0(InputBits[555]),
   .I1(InputBits[1289]),
   .I2(InputBits[902]),
   .I3(InputBits[247]),
   .I4(InputBits[413]),
   .I5(InputBits[1220])
);
LUT6 #(
   .INIT(64'b0111101110111011111111011110011100100011010101111000111111100111)  
) LUT6_1043 (
   .O(gates[176]),
   .I0(InputBits[1476]),
   .I1(InputBits[1456]),
   .I2(InputBits[689]),
   .I3(InputBits[1308]),
   .I4(InputBits[1593]),
   .I5(InputBits[1113])
);
LUT6 #(
   .INIT(64'b1101001001111000011100101101110011101000111111110001100010101111)  
) LUT6_1044 (
   .O(gates[956]),
   .I0(InputBits[1543]),
   .I1(InputBits[1604]),
   .I2(InputBits[1695]),
   .I3(InputBits[718]),
   .I4(InputBits[856]),
   .I5(InputBits[1557])
);
LUT6 #(
   .INIT(64'b1011011011000110100001001000110010111111110111101101011011000111)  
) LUT6_1045 (
   .O(gates[498]),
   .I0(InputBits[1614]),
   .I1(InputBits[145]),
   .I2(InputBits[1293]),
   .I3(InputBits[676]),
   .I4(InputBits[1054]),
   .I5(InputBits[406])
);
LUT6 #(
   .INIT(64'b0100011000011001000100110001001111010110000001110111110010001110)  
) LUT6_1046 (
   .O(gates[483]),
   .I0(InputBits[1540]),
   .I1(InputBits[1676]),
   .I2(InputBits[488]),
   .I3(InputBits[1706]),
   .I4(InputBits[576]),
   .I5(InputBits[1132])
);
LUT6 #(
   .INIT(64'b1111101010100110011111111010101011001010110000000111011001110111)  
) LUT6_1047 (
   .O(gates[629]),
   .I0(InputBits[783]),
   .I1(InputBits[457]),
   .I2(InputBits[66]),
   .I3(InputBits[1415]),
   .I4(InputBits[347]),
   .I5(InputBits[776])
);
LUT6 #(
   .INIT(64'b0000100001011001010111110000000001001001110100001111111111001111)  
) LUT6_1048 (
   .O(gates[947]),
   .I0(InputBits[6]),
   .I1(InputBits[1646]),
   .I2(InputBits[1702]),
   .I3(InputBits[311]),
   .I4(InputBits[329]),
   .I5(InputBits[565])
);
LUT6 #(
   .INIT(64'b1011111010100101011111001011100100001101110010110010111101111011)  
) LUT6_1049 (
   .O(gates[256]),
   .I0(InputBits[446]),
   .I1(InputBits[1661]),
   .I2(InputBits[560]),
   .I3(InputBits[303]),
   .I4(InputBits[763]),
   .I5(InputBits[592])
);
LUT6 #(
   .INIT(64'b1110100000101110010101110001110100101010010100010110110101001100)  
) LUT6_1050 (
   .O(gates[372]),
   .I0(InputBits[26]),
   .I1(InputBits[1096]),
   .I2(InputBits[49]),
   .I3(InputBits[1171]),
   .I4(InputBits[1480]),
   .I5(InputBits[1209])
);
LUT6 #(
   .INIT(64'b1110010111111111000110101000101100110001101001000101010000010000)  
) LUT6_1051 (
   .O(gates[1487]),
   .I0(InputBits[1242]),
   .I1(InputBits[1]),
   .I2(InputBits[254]),
   .I3(InputBits[480]),
   .I4(InputBits[1189]),
   .I5(InputBits[653])
);
LUT6 #(
   .INIT(64'b0000001000010111000100011111000000010101110011001010011100010001)  
) LUT6_1052 (
   .O(gates[1540]),
   .I0(InputBits[176]),
   .I1(InputBits[1004]),
   .I2(InputBits[1644]),
   .I3(InputBits[211]),
   .I4(InputBits[191]),
   .I5(InputBits[1060])
);
LUT6 #(
   .INIT(64'b1110010000111001010000011011010111110100000110011011110111011001)  
) LUT6_1053 (
   .O(gates[920]),
   .I0(InputBits[612]),
   .I1(InputBits[425]),
   .I2(InputBits[581]),
   .I3(InputBits[720]),
   .I4(InputBits[1130]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1000011110000010111101010010010010111100100011000000000010000011)  
) LUT6_1054 (
   .O(gates[1330]),
   .I0(InputBits[1598]),
   .I1(InputBits[1579]),
   .I2(InputBits[1530]),
   .I3(InputBits[1473]),
   .I4(InputBits[1616]),
   .I5(InputBits[1277])
);
LUT6 #(
   .INIT(64'b1001111010010010010111000100000011111111011010110100110001001000)  
) LUT6_1055 (
   .O(gates[1284]),
   .I0(InputBits[517]),
   .I1(InputBits[1726]),
   .I2(InputBits[1694]),
   .I3(InputBits[1566]),
   .I4(InputBits[647]),
   .I5(InputBits[1716])
);
LUT6 #(
   .INIT(64'b0011101011011110101111110010001100001010010100101110100011110001)  
) LUT6_1056 (
   .O(gates[428]),
   .I0(InputBits[683]),
   .I1(InputBits[313]),
   .I2(InputBits[1599]),
   .I3(InputBits[1069]),
   .I4(InputBits[208]),
   .I5(InputBits[1410])
);
LUT6 #(
   .INIT(64'b0010101011111100111110000101111111111001011111101011010110011101)  
) LUT6_1057 (
   .O(gates[887]),
   .I0(InputBits[355]),
   .I1(InputBits[235]),
   .I2(InputBits[323]),
   .I3(InputBits[1207]),
   .I4(InputBits[1521]),
   .I5(InputBits[833])
);
LUT6 #(
   .INIT(64'b1011111111110011111010111011101011010101001000001001111101010000)  
) LUT6_1058 (
   .O(gates[99]),
   .I0(InputBits[1383]),
   .I1(InputBits[709]),
   .I2(InputBits[135]),
   .I3(InputBits[1409]),
   .I4(InputBits[1709]),
   .I5(InputBits[1156])
);
LUT6 #(
   .INIT(64'b0101001100011111101111110000100101011101101011100011100000110100)  
) LUT6_1059 (
   .O(gates[1160]),
   .I0(InputBits[545]),
   .I1(InputBits[427]),
   .I2(InputBits[947]),
   .I3(InputBits[1363]),
   .I4(InputBits[838]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1011000110101101100101110111010000110001011010001010110000100010)  
) LUT6_1060 (
   .O(gates[72]),
   .I0(InputBits[1248]),
   .I1(InputBits[1320]),
   .I2(InputBits[1667]),
   .I3(InputBits[1450]),
   .I4(InputBits[285]),
   .I5(InputBits[853])
);
LUT6 #(
   .INIT(64'b0111000001100111010100011010101111001100001100110111110011001100)  
) LUT6_1061 (
   .O(gates[869]),
   .I0(InputBits[514]),
   .I1(InputBits[1590]),
   .I2(InputBits[268]),
   .I3(InputBits[500]),
   .I4(InputBits[712]),
   .I5(InputBits[982])
);
LUT6 #(
   .INIT(64'b1110011101001001001001100010011101001101011111101110110110100000)  
) LUT6_1062 (
   .O(gates[500]),
   .I0(InputBits[1396]),
   .I1(InputBits[1255]),
   .I2(InputBits[1649]),
   .I3(InputBits[473]),
   .I4(InputBits[106]),
   .I5(InputBits[1520])
);
LUT6 #(
   .INIT(64'b0111101000110110011001100011011000101000111001010101111101111110)  
) LUT6_1063 (
   .O(gates[1496]),
   .I0(InputBits[750]),
   .I1(InputBits[1486]),
   .I2(InputBits[51]),
   .I3(InputBits[509]),
   .I4(InputBits[37]),
   .I5(InputBits[378])
);
LUT6 #(
   .INIT(64'b1001011101011100010000011011101101011101101110100100010001101011)  
) LUT6_1064 (
   .O(gates[1221]),
   .I0(InputBits[202]),
   .I1(InputBits[467]),
   .I2(InputBits[127]),
   .I3(InputBits[525]),
   .I4(InputBits[1226]),
   .I5(InputBits[1442])
);
LUT6 #(
   .INIT(64'b0111010000011001000000001001100000101000110010001001000111101010)  
) LUT6_1065 (
   .O(gates[1200]),
   .I0(InputBits[861]),
   .I1(InputBits[552]),
   .I2(InputBits[142]),
   .I3(InputBits[43]),
   .I4(InputBits[656]),
   .I5(InputBits[727])
);
LUT6 #(
   .INIT(64'b1101001111010111100001001001101101000010101101010100010011101011)  
) LUT6_1066 (
   .O(gates[790]),
   .I0(InputBits[215]),
   .I1(InputBits[1205]),
   .I2(InputBits[301]),
   .I3(InputBits[974]),
   .I4(InputBits[1180]),
   .I5(InputBits[249])
);
LUT6 #(
   .INIT(64'b1000001010001111100010001011111001110101010011011001100001111101)  
) LUT6_1067 (
   .O(gates[533]),
   .I0(InputBits[760]),
   .I1(InputBits[802]),
   .I2(InputBits[929]),
   .I3(InputBits[702]),
   .I4(InputBits[889]),
   .I5(InputBits[1104])
);
LUT6 #(
   .INIT(64'b1110111110000000100111100101101010100111010100010011001110100101)  
) LUT6_1068 (
   .O(gates[918]),
   .I0(InputBits[1430]),
   .I1(InputBits[793]),
   .I2(InputBits[691]),
   .I3(InputBits[1090]),
   .I4(InputBits[439]),
   .I5(InputBits[1697])
);
LUT6 #(
   .INIT(64'b1110101110000111100101011100110010101010101000000110000100101110)  
) LUT6_1069 (
   .O(gates[1413]),
   .I0(InputBits[1078]),
   .I1(InputBits[1655]),
   .I2(InputBits[71]),
   .I3(InputBits[1618]),
   .I4(InputBits[664]),
   .I5(InputBits[586])
);
LUT6 #(
   .INIT(64'b0010011100000111010100110110101010110010001010000010011111000111)  
) LUT6_1070 (
   .O(gates[1122]),
   .I0(InputBits[904]),
   .I1(InputBits[909]),
   .I2(InputBits[642]),
   .I3(InputBits[161]),
   .I4(InputBits[1299]),
   .I5(InputBits[226])
);
LUT6 #(
   .INIT(64'b1010011001011010101010110010101110100000011100001100001010110111)  
) LUT6_1071 (
   .O(gates[1275]),
   .I0(InputBits[108]),
   .I1(InputBits[1333]),
   .I2(InputBits[128]),
   .I3(InputBits[602]),
   .I4(InputBits[56]),
   .I5(InputBits[858])
);
LUT6 #(
   .INIT(64'b1000001010110100101101111001111000011000100110110101011110101001)  
) LUT6_1072 (
   .O(gates[1108]),
   .I0(InputBits[1011]),
   .I1(InputBits[1491]),
   .I2(InputBits[280]),
   .I3(InputBits[11]),
   .I4(InputBits[829]),
   .I5(InputBits[1326])
);
LUT6 #(
   .INIT(64'b1010010111000100101011111100000001011001100010010000111000100111)  
) LUT6_1073 (
   .O(gates[1053]),
   .I0(InputBits[260]),
   .I1(InputBits[1082]),
   .I2(InputBits[534]),
   .I3(InputBits[532]),
   .I4(InputBits[1546]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0001111010000101100011010100011101111110110011011001101011011001)  
) LUT6_1074 (
   .O(gates[414]),
   .I0(InputBits[629]),
   .I1(InputBits[743]),
   .I2(InputBits[1606]),
   .I3(InputBits[1463]),
   .I4(InputBits[808]),
   .I5(InputBits[781])
);
LUT6 #(
   .INIT(64'b0010110100001100011000011101101011111110000111101101101010011010)  
) LUT6_1075 (
   .O(gates[462]),
   .I0(InputBits[1353]),
   .I1(InputBits[738]),
   .I2(InputBits[152]),
   .I3(InputBits[956]),
   .I4(InputBits[1548]),
   .I5(InputBits[1049])
);
LUT6 #(
   .INIT(64'b0010001111100100111000101100111110111010111111110100010111101111)  
) LUT6_1076 (
   .O(gates[1014]),
   .I0(InputBits[1533]),
   .I1(InputBits[337]),
   .I2(InputBits[635]),
   .I3(InputBits[222]),
   .I4(InputBits[489]),
   .I5(InputBits[991])
);
LUT6 #(
   .INIT(64'b0011000101011111011100111010110011100110011010001000000000010010)  
) LUT6_1077 (
   .O(gates[843]),
   .I0(InputBits[1258]),
   .I1(InputBits[939]),
   .I2(InputBits[1169]),
   .I3(InputBits[962]),
   .I4(InputBits[1022]),
   .I5(InputBits[1111])
);
LUT6 #(
   .INIT(64'b1010001111111001010000110111001110001111111101100010101101010000)  
) LUT6_1078 (
   .O(gates[1491]),
   .I0(InputBits[1457]),
   .I1(InputBits[774]),
   .I2(InputBits[1179]),
   .I3(InputBits[410]),
   .I4(InputBits[45]),
   .I5(InputBits[1685])
);
LUT6 #(
   .INIT(64'b0000100000100100110101000001000111111110001100111000111001100110)  
) LUT6_1079 (
   .O(gates[1362]),
   .I0(InputBits[185]),
   .I1(InputBits[1425]),
   .I2(InputBits[1098]),
   .I3(InputBits[1195]),
   .I4(InputBits[1101]),
   .I5(InputBits[972])
);
LUT6 #(
   .INIT(64'b0110110001110001111001010010001011011110111101010000110001101000)  
) LUT6_1080 (
   .O(gates[1209]),
   .I0(InputBits[993]),
   .I1(InputBits[527]),
   .I2(InputBits[295]),
   .I3(InputBits[1501]),
   .I4(InputBits[1058]),
   .I5(InputBits[1138])
);
LUT6 #(
   .INIT(64'b1010110111111110101111111100111011011111010101100110101001111100)  
) LUT6_1081 (
   .O(gates[632]),
   .I0(InputBits[409]),
   .I1(InputBits[1547]),
   .I2(InputBits[1692]),
   .I3(InputBits[1070]),
   .I4(InputBits[1158]),
   .I5(InputBits[1263])
);
LUT6 #(
   .INIT(64'b1101111011000100000100010111111100110001001111101101011011010011)  
) LUT6_1082 (
   .O(gates[263]),
   .I0(InputBits[869]),
   .I1(InputBits[916]),
   .I2(InputBits[64]),
   .I3(InputBits[1711]),
   .I4(InputBits[551]),
   .I5(InputBits[1141])
);
LUT6 #(
   .INIT(64'b0001111011110111100101100101110111000101100000111111100000000000)  
) LUT6_1083 (
   .O(gates[1371]),
   .I0(InputBits[1325]),
   .I1(InputBits[756]),
   .I2(InputBits[1523]),
   .I3(InputBits[643]),
   .I4(InputBits[138]),
   .I5(InputBits[1001])
);
LUT6 #(
   .INIT(64'b0010000001110110100001110011111001101111011100110010111110111010)  
) LUT6_1084 (
   .O(gates[991]),
   .I0(InputBits[1392]),
   .I1(InputBits[251]),
   .I2(InputBits[733]),
   .I3(InputBits[183]),
   .I4(InputBits[231]),
   .I5(InputBits[470])
);
LUT6 #(
   .INIT(64'b1000110000001000000110001010000011100100100100110010001101011101)  
) LUT6_1085 (
   .O(gates[394]),
   .I0(InputBits[294]),
   .I1(InputBits[1399]),
   .I2(InputBits[765]),
   .I3(InputBits[1094]),
   .I4(InputBits[1185]),
   .I5(InputBits[885])
);
LUT6 #(
   .INIT(64'b1111011100001111011011011100110110110101010101111011001000110011)  
) LUT6_1086 (
   .O(gates[514]),
   .I0(InputBits[585]),
   .I1(InputBits[1233]),
   .I2(InputBits[716]),
   .I3(InputBits[1670]),
   .I4(InputBits[812]),
   .I5(InputBits[1218])
);
LUT6 #(
   .INIT(64'b0000001001100100011101111000111001011001110010011011101010001100)  
) LUT6_1087 (
   .O(gates[610]),
   .I0(InputBits[1500]),
   .I1(InputBits[1704]),
   .I2(InputBits[445]),
   .I3(InputBits[882]),
   .I4(InputBits[976]),
   .I5(InputBits[890])
);
LUT6 #(
   .INIT(64'b1011000110011011001000001100100011101010100100000001000101011000)  
) LUT6_1088 (
   .O(gates[725]),
   .I0(InputBits[1576]),
   .I1(InputBits[1134]),
   .I2(InputBits[1485]),
   .I3(InputBits[874]),
   .I4(InputBits[1516]),
   .I5(InputBits[1235])
);
LUT6 #(
   .INIT(64'b0000010110000001100000010101001111111010111011100110000111101101)  
) LUT6_1089 (
   .O(gates[931]),
   .I0(InputBits[1717]),
   .I1(InputBits[384]),
   .I2(InputBits[855]),
   .I3(InputBits[424]),
   .I4(InputBits[1542]),
   .I5(InputBits[344])
);
LUT6 #(
   .INIT(64'b0001100101010110110110001111001111001010001000011101001010100000)  
) LUT6_1090 (
   .O(gates[513]),
   .I0(InputBits[1511]),
   .I1(InputBits[374]),
   .I2(InputBits[930]),
   .I3(InputBits[182]),
   .I4(InputBits[393]),
   .I5(InputBits[1588])
);
LUT6 #(
   .INIT(64'b1110111011110100101010011110101011010101111011010001110101110100)  
) LUT6_1091 (
   .O(gates[615]),
   .I0(InputBits[403]),
   .I1(InputBits[407]),
   .I2(InputBits[1578]),
   .I3(InputBits[1006]),
   .I4(InputBits[54]),
   .I5(InputBits[415])
);
LUT6 #(
   .INIT(64'b1011000001111111100111010011000100011100010111010000000001100101)  
) LUT6_1092 (
   .O(gates[50]),
   .I0(InputBits[836]),
   .I1(InputBits[225]),
   .I2(InputBits[1668]),
   .I3(InputBits[1689]),
   .I4(InputBits[567]),
   .I5(InputBits[1264])
);
LUT6 #(
   .INIT(64'b0110011011100100011111110000010001000101000100000011111000101111)  
) LUT6_1093 (
   .O(gates[476]),
   .I0(InputBits[309]),
   .I1(InputBits[725]),
   .I2(InputBits[1659]),
   .I3(InputBits[48]),
   .I4(InputBits[875]),
   .I5(InputBits[678])
);
LUT6 #(
   .INIT(64'b0111101000100100101010111101100101110001001111001000111010011001)  
) LUT6_1094 (
   .O(gates[1198]),
   .I0(InputBits[1388]),
   .I1(InputBits[326]),
   .I2(InputBits[1041]),
   .I3(InputBits[826]),
   .I4(InputBits[707]),
   .I5(InputBits[1216])
);
LUT6 #(
   .INIT(64'b0000000001101000110110101000111110110100010101100100001010000111)  
) LUT6_1095 (
   .O(gates[1519]),
   .I0(InputBits[820]),
   .I1(InputBits[381]),
   .I2(InputBits[701]),
   .I3(InputBits[1204]),
   .I4(InputBits[494]),
   .I5(InputBits[103])
);
LUT6 #(
   .INIT(64'b0011100000011110010010001000001100110110111101101000101111001001)  
) LUT6_1096 (
   .O(gates[1409]),
   .I0(InputBits[1357]),
   .I1(InputBits[1642]),
   .I2(InputBits[88]),
   .I3(InputBits[957]),
   .I4(InputBits[10]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1110100001111110001110101110000101000111011100000111000000001111)  
) LUT6_1097 (
   .O(gates[797]),
   .I0(InputBits[502]),
   .I1(InputBits[241]),
   .I2(InputBits[80]),
   .I3(InputBits[806]),
   .I4(InputBits[1443]),
   .I5(InputBits[620])
);
LUT6 #(
   .INIT(64'b0010110110100011111101010010101101000110001110111010101000000100)  
) LUT6_1098 (
   .O(gates[1077]),
   .I0(InputBits[1083]),
   .I1(InputBits[317]),
   .I2(InputBits[935]),
   .I3(InputBits[1008]),
   .I4(InputBits[503]),
   .I5(InputBits[1531])
);
LUT6 #(
   .INIT(64'b0100010101000101101011000100101001010100001011100101010110101001)  
) LUT6_1099 (
   .O(gates[1136]),
   .I0(InputBits[78]),
   .I1(InputBits[1088]),
   .I2(InputBits[1322]),
   .I3(InputBits[1380]),
   .I4(InputBits[387]),
   .I5(InputBits[958])
);
LUT6 #(
   .INIT(64'b1110110100101111000000100001000111110001111111010010010000100111)  
) LUT6_1100 (
   .O(gates[1175]),
   .I0(InputBits[487]),
   .I1(InputBits[450]),
   .I2(InputBits[151]),
   .I3(InputBits[284]),
   .I4(InputBits[1273]),
   .I5(InputBits[233])
);
LUT6 #(
   .INIT(64'b1011001010110010110001110110001110100110010011111110100101011000)  
) LUT6_1101 (
   .O(gates[293]),
   .I0(InputBits[631]),
   .I1(InputBits[1285]),
   .I2(InputBits[47]),
   .I3(InputBits[452]),
   .I4(InputBits[405]),
   .I5(InputBits[368])
);
LUT6 #(
   .INIT(64'b1000110101010101100001000001111011000110101100000010011110010110)  
) LUT6_1102 (
   .O(gates[1272]),
   .I0(InputBits[800]),
   .I1(InputBits[1228]),
   .I2(InputBits[357]),
   .I3(InputBits[609]),
   .I4(InputBits[737]),
   .I5(InputBits[442])
);
LUT6 #(
   .INIT(64'b1101000010000110011011001101001011010001111001010000000100011111)  
) LUT6_1103 (
   .O(gates[1299]),
   .I0(InputBits[1467]),
   .I1(InputBits[125]),
   .I2(InputBits[398]),
   .I3(InputBits[1324]),
   .I4(InputBits[1202]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1000000000100110011100010110110100100000010110000110011111100001)  
) LUT6_1104 (
   .O(gates[1236]),
   .I0(InputBits[899]),
   .I1(InputBits[522]),
   .I2(InputBits[481]),
   .I3(InputBits[484]),
   .I4(InputBits[192]),
   .I5(InputBits[187])
);
LUT6 #(
   .INIT(64'b0010001100010011100010110101010111010111000001110111011100110010)  
) LUT6_1105 (
   .O(gates[967]),
   .I0(InputBits[1573]),
   .I1(InputBits[1030]),
   .I2(InputBits[69]),
   .I3(InputBits[244]),
   .I4(InputBits[1337]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0100101110011111011001011111010000100010110111000101011111000000)  
) LUT6_1106 (
   .O(gates[322]),
   .I0(InputBits[140]),
   .I1(InputBits[979]),
   .I2(InputBits[823]),
   .I3(InputBits[1428]),
   .I4(InputBits[149]),
   .I5(InputBits[1459])
);
LUT6 #(
   .INIT(64'b0000110000110100110111100100001101110011110010110110101100001111)  
) LUT6_1107 (
   .O(gates[645]),
   .I0(InputBits[1529]),
   .I1(InputBits[1332]),
   .I2(InputBits[194]),
   .I3(InputBits[897]),
   .I4(InputBits[573]),
   .I5(InputBits[668])
);
LUT6 #(
   .INIT(64'b1011010100001000011000010001100100110011010011111110011110001000)  
) LUT6_1108 (
   .O(gates[1326]),
   .I0(InputBits[1146]),
   .I1(InputBits[1129]),
   .I2(InputBits[1597]),
   .I3(InputBits[1015]),
   .I4(InputBits[385]),
   .I5(InputBits[754])
);
LUT6 #(
   .INIT(64'b1110110000000011110100111111101000111010101110001110011000010000)  
) LUT6_1109 (
   .O(gates[469]),
   .I0(InputBits[86]),
   .I1(InputBits[360]),
   .I2(InputBits[1407]),
   .I3(InputBits[1109]),
   .I4(InputBits[1182]),
   .I5(InputBits[1629])
);
LUT6 #(
   .INIT(64'b0001000010001010000010011101101100001111000100111011111010101001)  
) LUT6_1110 (
   .O(gates[635]),
   .I0(InputBits[513]),
   .I1(InputBits[171]),
   .I2(InputBits[1003]),
   .I3(InputBits[1348]),
   .I4(InputBits[1117]),
   .I5(InputBits[610])
);
LUT6 #(
   .INIT(64'b0110100010000111101011111011010100010110010110010110001110000010)  
) LUT6_1111 (
   .O(gates[575]),
   .I0(InputBits[263]),
   .I1(InputBits[792]),
   .I2(InputBits[539]),
   .I3(InputBits[282]),
   .I4(InputBits[159]),
   .I5(InputBits[463])
);
LUT6 #(
   .INIT(64'b1101111110100100011000101000001110010111111000000000011110001010)  
) LUT6_1112 (
   .O(gates[1088]),
   .I0(InputBits[351]),
   .I1(InputBits[1231]),
   .I2(InputBits[1535]),
   .I3(InputBits[117]),
   .I4(InputBits[1422]),
   .I5(InputBits[1680])
);
LUT6 #(
   .INIT(64'b1100101001011111001000010011100110101100010101011010011110111110)  
) LUT6_1113 (
   .O(gates[1382]),
   .I0(InputBits[768]),
   .I1(InputBits[770]),
   .I2(InputBits[130]),
   .I3(InputBits[456]),
   .I4(InputBits[336]),
   .I5(InputBits[1494])
);
LUT6 #(
   .INIT(64'b0011001011001110101010110011010110101011000000011110110000100101)  
) LUT6_1114 (
   .O(gates[1176]),
   .I0(InputBits[1267]),
   .I1(InputBits[1213]),
   .I2(InputBits[713]),
   .I3(InputBits[1478]),
   .I4(InputBits[772]),
   .I5(InputBits[714])
);
LUT6 #(
   .INIT(64'b0110100111100011111010001101010101011001000010111000001111100011)  
) LUT6_1115 (
   .O(gates[1452]),
   .I0(InputBits[1624]),
   .I1(InputBits[1634]),
   .I2(InputBits[1359]),
   .I3(InputBits[989]),
   .I4(InputBits[1351]),
   .I5(InputBits[986])
);
LUT6 #(
   .INIT(64'b0000101010000101010010001011111111101110110111101000110111101111)  
) LUT6_1116 (
   .O(gates[1039]),
   .I0(InputBits[1666]),
   .I1(InputBits[1177]),
   .I2(InputBits[1297]),
   .I3(InputBits[600]),
   .I4(InputBits[38]),
   .I5(InputBits[844])
);
LUT6 #(
   .INIT(64'b0111010001001010111000111100000110110110111001111001010101000001)  
) LUT6_1117 (
   .O(gates[979]),
   .I0(InputBits[156]),
   .I1(InputBits[1436]),
   .I2(InputBits[1052]),
   .I3(InputBits[1281]),
   .I4(InputBits[547]),
   .I5(InputBits[1024])
);
LUT6 #(
   .INIT(64'b0101110111001111111001010110011100110001101010111010101111100000)  
) LUT6_1118 (
   .O(gates[709]),
   .I0(InputBits[1687]),
   .I1(InputBits[461]),
   .I2(InputBits[1627]),
   .I3(InputBits[1513]),
   .I4(InputBits[165]),
   .I5(InputBits[180])
);
LUT6 #(
   .INIT(64'b0010010000111101101111110100111001011010101101000101101101101111)  
) LUT6_1119 (
   .O(gates[1005]),
   .I0(InputBits[1498]),
   .I1(InputBits[651]),
   .I2(InputBits[622]),
   .I3(InputBits[333]),
   .I4(InputBits[941]),
   .I5(InputBits[475])
);
LUT6 #(
   .INIT(64'b0010111011011000011000011100001010100110010110101011010111111010)  
) LUT6_1120 (
   .O(gates[28]),
   .I0(InputBits[1712]),
   .I1(InputBits[731]),
   .I2(InputBits[814]),
   .I3(InputBits[375]),
   .I4(InputBits[1092]),
   .I5(InputBits[40])
);
LUT6 #(
   .INIT(64'b0010010111000001100011001111011100100100100000010101000100100001)  
) LUT6_1121 (
   .O(gates[40]),
   .I0(InputBits[1261]),
   .I1(InputBits[195]),
   .I2(InputBits[253]),
   .I3(InputBits[184]),
   .I4(InputBits[1247]),
   .I5(InputBits[55])
);
LUT6 #(
   .INIT(64'b1100110011000000001011100101011100101110110010110000001101011110)  
) LUT6_1122 (
   .O(gates[310]),
   .I0(InputBits[496]),
   .I1(InputBits[1127]),
   .I2(InputBits[1268]),
   .I3(InputBits[1446]),
   .I4(InputBits[934]),
   .I5(InputBits[849])
);
LUT6 #(
   .INIT(64'b1100010111111010111011001111100101001100011110011001110010001010)  
) LUT6_1123 (
   .O(gates[192]),
   .I0(InputBits[1100]),
   .I1(InputBits[1622]),
   .I2(InputBits[954]),
   .I3(InputBits[1148]),
   .I4(InputBits[1400]),
   .I5(InputBits[616])
);
LUT6 #(
   .INIT(64'b0001010011111010000100010110010100010100010001100011001111110011)  
) LUT6_1124 (
   .O(gates[589]),
   .I0(InputBits[1056]),
   .I1(InputBits[411]),
   .I2(InputBits[454]),
   .I3(InputBits[110]),
   .I4(InputBits[354]),
   .I5(InputBits[1072])
);
LUT6 #(
   .INIT(64'b1001111110000000000111000001000001111011111000001010010000100000)  
) LUT6_1125 (
   .O(gates[1337]),
   .I0(InputBits[227]),
   .I1(InputBits[884]),
   .I2(InputBits[1143]),
   .I3(InputBits[697]),
   .I4(InputBits[1187]),
   .I5(InputBits[951])
);
LUT6 #(
   .INIT(64'b0110111110111010011001010001101110100001011110000110101010011101)  
) LUT6_1126 (
   .O(gates[699]),
   .I0(InputBits[529]),
   .I1(InputBits[918]),
   .I2(InputBits[1043]),
   .I3(InputBits[1654]),
   .I4(InputBits[1567]),
   .I5(InputBits[615])
);
LUT6 #(
   .INIT(64'b0000101001110101011011101011101100011000010111100001010101110101)  
) LUT6_1127 (
   .O(gates[215]),
   .I0(InputBits[1341]),
   .I1(InputBits[780]),
   .I2(InputBits[867]),
   .I3(InputBits[1366]),
   .I4(InputBits[435]),
   .I5(InputBits[35])
);
LUT6 #(
   .INIT(64'b0000101101001000000001000010000000101001100000110010100010010101)  
) LUT6_1128 (
   .O(gates[687]),
   .I0(InputBits[1699]),
   .I1(InputBits[97]),
   .I2(InputBits[846]),
   .I3(InputBits[1640]),
   .I4(InputBits[937]),
   .I5(InputBits[907])
);
LUT6 #(
   .INIT(64'b1110011011010101101010111010011100000010000111110000100110000001)  
) LUT6_1129 (
   .O(gates[1115]),
   .I0(InputBits[498]),
   .I1(InputBits[1378]),
   .I2(InputBits[554]),
   .I3(InputBits[154]),
   .I4(InputBits[746]),
   .I5(InputBits[472])
);
LUT6 #(
   .INIT(64'b0000100101110110000011001100110101100010001001001111100000011001)  
) LUT6_1130 (
   .O(gates[960]),
   .I0(InputBits[926]),
   .I1(InputBits[914]),
   .I2(InputBits[1317]),
   .I3(InputBits[190]),
   .I4(InputBits[1039]),
   .I5(InputBits[556])
);
LUT6 #(
   .INIT(64'b1011100011110101100100001101100010101010100101100001111000100110)  
) LUT6_1131 (
   .O(gates[818]),
   .I0(InputBits[535]),
   .I1(InputBits[307]),
   .I2(InputBits[797]),
   .I3(InputBits[569]),
   .I4(InputBits[342]),
   .I5(InputBits[1105])
);
LUT6 #(
   .INIT(64'b1101010001111101000100111100111110100001010101011001010011010101)  
) LUT6_1132 (
   .O(gates[150]),
   .I0(InputBits[297]),
   .I1(InputBits[1136]),
   .I2(InputBits[817]),
   .I3(InputBits[1503]),
   .I4(InputBits[401]),
   .I5(InputBits[1390])
);
LUT6 #(
   .INIT(64'b0000011010111110000101111000011000100010000111110100110101111001)  
) LUT6_1133 (
   .O(gates[1038]),
   .I0(InputBits[693]),
   .I1(InputBits[1223]),
   .I2(InputBits[680]),
   .I3(InputBits[1620]),
   .I4(InputBits[1526]),
   .I5(InputBits[1254])
);
LUT6 #(
   .INIT(64'b0010111000001011110010111001011010010011011011101001100110011011)  
) LUT6_1134 (
   .O(gates[245]),
   .I0(InputBits[1544]),
   .I1(InputBits[1723]),
   .I2(InputBits[1076]),
   .I3(InputBits[723]),
   .I4(InputBits[872]),
   .I5(InputBits[396])
);
LUT6 #(
   .INIT(64'b0111110111000010011011000000100011000011100011001011110000111100)  
) LUT6_1135 (
   .O(gates[543]),
   .I0(InputBits[82]),
   .I1(InputBits[1211]),
   .I2(InputBits[1373]),
   .I3(InputBits[239]),
   .I4(InputBits[638]),
   .I5(InputBits[1081])
);
LUT6 #(
   .INIT(64'b0010100101111111011010011101000000011001111100111110001100111111)  
) LUT6_1136 (
   .O(gates[267]),
   .I0(InputBits[537]),
   .I1(InputBits[1413]),
   .I2(InputBits[944]),
   .I3(InputBits[901]),
   .I4(InputBits[1636]),
   .I5(InputBits[1250])
);
LUT6 #(
   .INIT(64'b1000101101010011000001010110011111111100000001010011111000110001)  
) LUT6_1137 (
   .O(gates[826]),
   .I0(InputBits[541]),
   .I1(InputBits[229]),
   .I2(InputBits[1284]),
   .I3(InputBits[124]),
   .I4(InputBits[594]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b1011100010011111110110101011001000010111010111000110011001110010)  
) LUT6_1138 (
   .O(gates[354]),
   .I0(InputBits[1462]),
   .I1(InputBits[1085]),
   .I2(InputBits[65]),
   .I3(InputBits[1145]),
   .I4(InputBits[686]),
   .I5(InputBits[1549])
);
LUT6 #(
   .INIT(64'b1100110000100011110100101001001000110100011000101110100010110000)  
) LUT6_1139 (
   .O(gates[1437]),
   .I0(InputBits[1420]),
   .I1(InputBits[1505]),
   .I2(InputBits[1612]),
   .I3(InputBits[1192]),
   .I4(InputBits[328]),
   .I5(InputBits[607])
);
LUT6 #(
   .INIT(64'b1000110101000010111101101100110101111111011110000110011011001010)  
) LUT6_1140 (
   .O(gates[1344]),
   .I0(InputBits[815]),
   .I1(InputBits[291]),
   .I2(InputBits[660]),
   .I3(InputBits[1116]),
   .I4(InputBits[370]),
   .I5(InputBits[999])
);
LUT6 #(
   .INIT(64'b1001110101111001011011000110110000011000110111001111100001100001)  
) LUT6_1141 (
   .O(gates[1064]),
   .I0(InputBits[1019]),
   .I1(InputBits[1361]),
   .I2(InputBits[1571]),
   .I3(InputBits[1045]),
   .I4(InputBits[960]),
   .I5(InputBits[61])
);
LUT6 #(
   .INIT(64'b1001010011101010010011001001000110001010000111011110000001101011)  
) LUT6_1142 (
   .O(gates[757]),
   .I0(InputBits[28]),
   .I1(InputBits[862]),
   .I2(InputBits[76]),
   .I3(InputBits[273]),
   .I4(InputBits[1050]),
   .I5(InputBits[1065])
);
LUT6 #(
   .INIT(64'b1100101100010010100010000010111011101000001110000001000010010001)  
) LUT6_1143 (
   .O(gates[332]),
   .I0(InputBits[739]),
   .I1(InputBits[1451]),
   .I2(InputBits[583]),
   .I3(InputBits[965]),
   .I4(InputBits[892]),
   .I5(InputBits[670])
);
LUT6 #(
   .INIT(64'b0110111100001000111101001000011101110000001111011100010011000011)  
) LUT6_1144 (
   .O(gates[9]),
   .I0(InputBits[23]),
   .I1(InputBits[1673]),
   .I2(InputBits[1585]),
   .I3(InputBits[1488]),
   .I4(InputBits[1063]),
   .I5(InputBits[1426])
);
LUT6 #(
   .INIT(64'b0111110100001110010111000111010101101110011010111101011110011011)  
) LUT6_1145 (
   .O(gates[1099]),
   .I0(InputBits[1483]),
   .I1(InputBits[596]),
   .I2(InputBits[1238]),
   .I3(InputBits[274]),
   .I4(InputBits[362]),
   .I5(InputBits[1033])
);
LUT6 #(
   .INIT(64'b1101110100110110011101011001100100110010010111101010101000011001)  
) LUT6_1146 (
   .O(gates[1217]),
   .I0(InputBits[1438]),
   .I1(InputBits[349]),
   .I2(InputBits[206]),
   .I3(InputBits[74]),
   .I4(InputBits[363]),
   .I5(InputBits[1200])
);
LUT6 #(
   .INIT(64'b1001111000000101011110100000010111110010100110101110111011101101)  
) LUT6_1147 (
   .O(gates[745]),
   .I0(InputBits[641]),
   .I1(InputBits[147]),
   .I2(InputBits[1682]),
   .I3(InputBits[1563]),
   .I4(InputBits[158]),
   .I5(InputBits[1595])
);
LUT6 #(
   .INIT(64'b1001001010011110110110101111001110110011001101110011100001110010)  
) LUT6_1148 (
   .O(gates[34]),
   .I0(InputBits[1107]),
   .I1(InputBits[865]),
   .I2(InputBits[1174]),
   .I3(InputBits[549]),
   .I4(InputBits[1609]),
   .I5(InputBits[571])
);
LUT6 #(
   .INIT(64'b0111110101010011100010101111111001001001110001100100001101010100)  
) LUT6_1149 (
   .O(gates[603]),
   .I0(InputBits[1339]),
   .I1(InputBits[1303]),
   .I2(InputBits[174]),
   .I3(InputBits[971]),
   .I4(InputBits[1330]),
   .I5(InputBits[1306])
);
LUT6 #(
   .INIT(64'b0100010011000010101101010010110111100011011100110110000101110001)  
) LUT6_1150 (
   .O(gates[90]),
   .I0(InputBits[933]),
   .I1(InputBits[1551]),
   .I2(InputBits[1017]),
   .I3(InputBits[219]),
   .I4(InputBits[932]),
   .I5(InputBits[1633])
);
LUT6 #(
   .INIT(64'b1110010111001001011001000010101110001101111101011101001001100101)  
) LUT6_1151 (
   .O(gates[620]),
   .I0(InputBits[1647]),
   .I1(InputBits[841]),
   .I2(InputBits[164]),
   .I3(InputBits[1165]),
   .I4(InputBits[1161]),
   .I5(InputBits[430])
);
LUT6 #(
   .INIT(64'b1010101100110101101100110111110101010010001000110101000101011001)  
) LUT6_1152 (
   .O(gates[565]),
   .I0(InputBits[508]),
   .I1(InputBits[1114]),
   .I2(InputBits[136]),
   .I3(InputBits[448]),
   .I4(InputBits[1714]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1010010100111010111011111101100001000010100111110010100001100111)  
) LUT6_1153 (
   .O(gates[1410]),
   .I0(InputBits[1077]),
   .I1(InputBits[1123]),
   .I2(InputBits[246]),
   .I3(InputBits[93]),
   .I4(InputBits[1343]),
   .I5(InputBits[1519])
);
LUT6 #(
   .INIT(64'b1011001101101111010111100001000101000110011110100011011011011100)  
) LUT6_1154 (
   .O(gates[1346]),
   .I0(InputBits[1372]),
   .I1(InputBits[1257]),
   .I2(InputBits[711]),
   .I3(InputBits[1608]),
   .I4(InputBits[1275]),
   .I5(InputBits[1360])
);
LUT6 #(
   .INIT(64'b1110011000110011100001100011100010010100100101010000011111100000)  
) LUT6_1155 (
   .O(gates[1434]),
   .I0(InputBits[1170]),
   .I1(InputBits[377]),
   .I2(InputBits[1387]),
   .I3(InputBits[961]),
   .I4(InputBits[1061]),
   .I5(InputBits[1079])
);
LUT6 #(
   .INIT(64'b0100100100101110000001011000000101100101001100011100011111110111)  
) LUT6_1156 (
   .O(gates[850]),
   .I0(InputBits[230]),
   .I1(InputBits[1584]),
   .I2(InputBits[983]),
   .I3(InputBits[893]),
   .I4(InputBits[1414]),
   .I5(InputBits[952])
);
LUT6 #(
   .INIT(64'b0110001001100001111010100111101000100101111011011011101010100001)  
) LUT6_1157 (
   .O(gates[1547]),
   .I0(InputBits[1166]),
   .I1(InputBits[1496]),
   .I2(InputBits[512]),
   .I3(InputBits[75]),
   .I4(InputBits[996]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0110111101011110111010110001001110110101101010001001011100001101)  
) LUT6_1158 (
   .O(gates[891]),
   .I0(InputBits[1554]),
   .I1(InputBits[1630]),
   .I2(InputBits[599]),
   .I3(InputBits[83]),
   .I4(InputBits[589]),
   .I5(InputBits[414])
);
LUT6 #(
   .INIT(64'b0000110000111001100011101011010100010000011111101101010001100111)  
) LUT6_1159 (
   .O(gates[1045]),
   .I0(InputBits[255]),
   .I1(InputBits[648]),
   .I2(InputBits[60]),
   .I3(InputBits[1582]),
   .I4(InputBits[1276]),
   .I5(InputBits[1510])
);
LUT6 #(
   .INIT(64'b1111110000101100100101011111110110001011000101011100111110110101)  
) LUT6_1160 (
   .O(gates[937]),
   .I0(InputBits[1377]),
   .I1(InputBits[177]),
   .I2(InputBits[518]),
   .I3(InputBits[832]),
   .I4(InputBits[1199]),
   .I5(InputBits[851])
);
LUT6 #(
   .INIT(64'b1001001001011011100101110100110010011101001000111101100011000010)  
) LUT6_1161 (
   .O(gates[1004]),
   .I0(InputBits[1617]),
   .I1(InputBits[1439]),
   .I2(InputBits[369]),
   .I3(InputBits[1701]),
   .I4(InputBits[1163]),
   .I5(InputBits[1487])
);
LUT6 #(
   .INIT(64'b1011100010000000001101001101101100110011010110001110101001010100)  
) LUT6_1162 (
   .O(gates[730]),
   .I0(InputBits[1037]),
   .I1(InputBits[105]),
   .I2(InputBits[870]),
   .I3(InputBits[148]),
   .I4(InputBits[1652]),
   .I5(InputBits[735])
);
LUT6 #(
   .INIT(64'b1010111111111100110010010000110011010100110101100010111101001000)  
) LUT6_1163 (
   .O(gates[16]),
   .I0(InputBits[759]),
   .I1(InputBits[531]),
   .I2(InputBits[661]),
   .I3(InputBits[261]),
   .I4(InputBits[905]),
   .I5(InputBits[399])
);
LUT6 #(
   .INIT(64'b1000011001111010110100111010001110001111101010000111001101100000)  
) LUT6_1164 (
   .O(gates[921]),
   .I0(InputBits[1288]),
   .I1(InputBits[955]),
   .I2(InputBits[1144]),
   .I3(InputBits[790]),
   .I4(InputBits[903]),
   .I5(InputBits[1032])
);
LUT6 #(
   .INIT(64'b1010110101010011110110011010001100010011001111111101111110101101)  
) LUT6_1165 (
   .O(gates[1360]),
   .I0(InputBits[1569]),
   .I1(InputBits[53]),
   .I2(InputBits[773]),
   .I3(InputBits[1418]),
   .I4(InputBits[1012]),
   .I5(InputBits[1444])
);
LUT6 #(
   .INIT(64'b1001000110110011011100001100010010100101001001000010011010010101)  
) LUT6_1166 (
   .O(gates[1013]),
   .I0(InputBits[886]),
   .I1(InputBits[1421]),
   .I2(InputBits[919]),
   .I3(InputBits[1677]),
   .I4(InputBits[1334]),
   .I5(InputBits[859])
);
LUT6 #(
   .INIT(64'b0000010000101010001111010111001101101010001011000001000100000100)  
) LUT6_1167 (
   .O(gates[1069]),
   .I0(InputBits[1369]),
   .I1(InputBits[1683]),
   .I2(InputBits[348]),
   .I3(InputBits[719]),
   .I4(InputBits[639]),
   .I5(InputBits[730])
);
LUT6 #(
   .INIT(64'b0100101001000010001101101100010101111010100110100011011110100100)  
) LUT6_1168 (
   .O(gates[233]),
   .I0(InputBits[1603]),
   .I1(InputBits[1537]),
   .I2(InputBits[447]),
   .I3(InputBits[1309]),
   .I4(InputBits[1212]),
   .I5(InputBits[633])
);
LUT6 #(
   .INIT(64'b1101011011100110110011101110000011001110001110101110110001010110)  
) LUT6_1169 (
   .O(gates[1224]),
   .I0(InputBits[533]),
   .I1(InputBits[223]),
   .I2(InputBits[112]),
   .I3(InputBits[304]),
   .I4(InputBits[784]),
   .I5(InputBits[559])
);
LUT6 #(
   .INIT(64'b0100011011100100111110110010001100001011111111100100010100110001)  
) LUT6_1170 (
   .O(gates[1490]),
   .I0(InputBits[579]),
   .I1(InputBits[1561]),
   .I2(InputBits[1221]),
   .I3(InputBits[804]),
   .I4(InputBits[1684]),
   .I5(InputBits[1346])
);
LUT6 #(
   .INIT(64'b1110110100010010011001001010000111000001100001100000010100001100)  
) LUT6_1171 (
   .O(gates[368]),
   .I0(InputBits[1556]),
   .I1(InputBits[879]),
   .I2(InputBits[490]),
   .I3(InputBits[1594]),
   .I4(InputBits[1027]),
   .I5(InputBits[205])
);
LUT6 #(
   .INIT(64'b0110001010001000101010010011010101110011111011001001110010100011)  
) LUT6_1172 (
   .O(gates[316]),
   .I0(InputBits[478]),
   .I1(InputBits[499]),
   .I2(InputBits[173]),
   .I3(InputBits[1230]),
   .I4(InputBits[1669]),
   .I5(InputBits[332])
);
LUT6 #(
   .INIT(64'b1111010000100110010100000011100010011111111001100000001100000110)  
) LUT6_1173 (
   .O(gates[994]),
   .I0(InputBits[1121]),
   .I1(InputBits[1352]),
   .I2(InputBits[1315]),
   .I3(InputBits[30]),
   .I4(InputBits[322]),
   .I5(InputBits[1384])
);
LUT6 #(
   .INIT(64'b1011111011001011010100011000111110110111111111010000110010011110)  
) LUT6_1174 (
   .O(gates[611]),
   .I0(InputBits[1304]),
   .I1(InputBits[1150]),
   .I2(InputBits[1638]),
   .I3(InputBits[672]),
   .I4(InputBits[1686]),
   .I5(InputBits[1464])
);
LUT6 #(
   .INIT(64'b1101011110010001000001010010100001101100101010000110000110111101)  
) LUT6_1175 (
   .O(gates[1370]),
   .I0(InputBits[614]),
   .I1(InputBits[1703]),
   .I2(InputBits[186]),
   .I3(InputBits[212]),
   .I4(InputBits[563]),
   .I5(InputBits[98])
);
LUT6 #(
   .INIT(64'b1000001001110111001011100100100010010001100010100000111100111001)  
) LUT6_1176 (
   .O(gates[849]),
   .I0(InputBits[682]),
   .I1(InputBits[133]),
   .I2(InputBits[839]),
   .I3(InputBits[1042]),
   .I4(InputBits[775]),
   .I5(InputBits[1294])
);
LUT6 #(
   .INIT(64'b0100001010010001111010111011111111000000011001000100011011101010)  
) LUT6_1177 (
   .O(gates[11]),
   .I0(InputBits[316]),
   .I1(InputBits[1099]),
   .I2(InputBits[830]),
   .I3(InputBits[1403]),
   .I4(InputBits[277]),
   .I5(InputBits[1240])
);
LUT6 #(
   .INIT(64'b0010010010011010100110000010011111111111001010111110100010100111)  
) LUT6_1178 (
   .O(gates[492]),
   .I0(InputBits[1149]),
   .I1(InputBits[1592]),
   .I2(InputBits[1621]),
   .I3(InputBits[1705]),
   .I4(InputBits[5]),
   .I5(InputBits[1645])
);
LUT6 #(
   .INIT(64'b0011001010011001011100010001101110111000000110111010111110000010)  
) LUT6_1179 (
   .O(gates[208]),
   .I0(InputBits[1481]),
   .I1(InputBits[207]),
   .I2(InputBits[613]),
   .I3(InputBits[1525]),
   .I4(InputBits[506]),
   .I5(InputBits[289])
);
LUT6 #(
   .INIT(64'b1110101011000111000001010000000110101011100101001110100110100100)  
) LUT6_1180 (
   .O(gates[842]),
   .I0(InputBits[1155]),
   .I1(InputBits[949]),
   .I2(InputBits[1243]),
   .I3(InputBits[1397]),
   .I4(InputBits[795]),
   .I5(InputBits[168])
);
LUT6 #(
   .INIT(64'b1001101010100010110010011011110111101111110101000101000011100100)  
) LUT6_1181 (
   .O(gates[511]),
   .I0(InputBits[924]),
   .I1(InputBits[1066]),
   .I2(InputBits[1663]),
   .I3(InputBits[492]),
   .I4(InputBits[25]),
   .I5(InputBits[1719])
);
LUT6 #(
   .INIT(64'b1101000011010100110011011010000100101100010111011011101010000101)  
) LUT6_1182 (
   .O(gates[1523]),
   .I0(InputBits[1382]),
   .I1(InputBits[864]),
   .I2(InputBits[591]),
   .I3(InputBits[1602]),
   .I4(InputBits[1290]),
   .I5(InputBits[969])
);
LUT6 #(
   .INIT(64'b0101010111000011010101100100101010010101011100001000010000001100)  
) LUT6_1183 (
   .O(gates[93]),
   .I0(InputBits[927]),
   .I1(InputBits[380]),
   .I2(InputBits[1164]),
   .I3(InputBits[1135]),
   .I4(InputBits[259]),
   .I5(InputBits[1172])
);
LUT6 #(
   .INIT(64'b0101101110010111001001101111011001000001010011111001111100101011)  
) LUT6_1184 (
   .O(gates[899]),
   .I0(InputBits[650]),
   .I1(InputBits[1411]),
   .I2(InputBits[658]),
   .I3(InputBits[1253]),
   .I4(InputBits[523]),
   .I5(InputBits[420])
);
LUT6 #(
   .INIT(64'b0111110110110001101111111111111110010110101100100100011000000010)  
) LUT6_1185 (
   .O(gates[292]),
   .I0(InputBits[1470]),
   .I1(InputBits[1449]),
   .I2(InputBits[1385]),
   .I3(InputBits[1517]),
   .I4(InputBits[418]),
   .I5(InputBits[1355])
);
LUT6 #(
   .INIT(64'b0001000001001000110101000001001000111011000110000000001110010011)  
) LUT6_1186 (
   .O(gates[291]),
   .I0(InputBits[436]),
   .I1(InputBits[1472]),
   .I2(InputBits[197]),
   .I3(InputBits[21]),
   .I4(InputBits[1658]),
   .I5(InputBits[1625])
);
LUT6 #(
   .INIT(64'b1011100100011111101110100000010100110000110101001000111100011101)  
) LUT6_1187 (
   .O(gates[374]),
   .I0(InputBits[747]),
   .I1(InputBits[1319]),
   .I2(InputBits[1126]),
   .I3(InputBits[203]),
   .I4(InputBits[67]),
   .I5(InputBits[267])
);
LUT6 #(
   .INIT(64'b0111100000111010110100011010101110101111011001001010110000001111)  
) LUT6_1188 (
   .O(gates[114]),
   .I0(InputBits[1190]),
   .I1(InputBits[1508]),
   .I2(InputBits[153]),
   .I3(InputBits[665]),
   .I4(InputBits[356]),
   .I5(InputBits[1301])
);
LUT6 #(
   .INIT(64'b1010101010001100110100001010110101100110100111100111111101101110)  
) LUT6_1189 (
   .O(gates[199]),
   .I0(InputBits[973]),
   .I1(InputBits[36]),
   .I2(InputBits[122]),
   .I3(InputBits[1181]),
   .I4(InputBits[479]),
   .I5(InputBits[644])
);
LUT6 #(
   .INIT(64'b0110101001000001010110100001100101111010011000100110010110011001)  
) LUT6_1190 (
   .O(gates[429]),
   .I0(InputBits[845]),
   .I1(InputBits[703]),
   .I2(InputBits[619]),
   .I3(InputBits[474]),
   .I4(InputBits[794]),
   .I5(InputBits[1447])
);
LUT6 #(
   .INIT(64'b1001101010100100100110100011101111001001100001111101010110110110)  
) LUT6_1191 (
   .O(gates[1306]),
   .I0(InputBits[1197]),
   .I1(InputBits[1168]),
   .I2(InputBits[1558]),
   .I3(InputBits[438]),
   .I4(InputBits[338]),
   .I5(InputBits[91])
);
LUT6 #(
   .INIT(64'b1001010110111101110001001011100011001011100100110110000000101011)  
) LUT6_1192 (
   .O(gates[1328]),
   .I0(InputBits[788]),
   .I1(InputBits[1455]),
   .I2(InputBits[963]),
   .I3(InputBits[1489]),
   .I4(InputBits[553]),
   .I5(InputBits[821])
);
LUT6 #(
   .INIT(64'b0000000001111111011100100000010011100101010001010010110011011010)  
) LUT6_1193 (
   .O(gates[1091]),
   .I0(InputBits[428]),
   .I1(InputBits[1545]),
   .I2(InputBits[468]),
   .I3(InputBits[422]),
   .I4(InputBits[199]),
   .I5(InputBits[72])
);
LUT6 #(
   .INIT(64'b1101001101010011101101000110111100101010110111001011010011100011)  
) LUT6_1194 (
   .O(gates[73]),
   .I0(InputBits[270]),
   .I1(InputBits[114]),
   .I2(InputBits[397]),
   .I3(InputBits[538]),
   .I4(InputBits[1475]),
   .I5(InputBits[372])
);
LUT6 #(
   .INIT(64'b0001111011100100000011011010110111010011010110110011110011000000)  
) LUT6_1195 (
   .O(gates[409]),
   .I0(InputBits[1298]),
   .I1(InputBits[1040]),
   .I2(InputBits[59]),
   .I3(InputBits[663]),
   .I4(InputBits[761]),
   .I5(InputBits[188])
);
LUT6 #(
   .INIT(64'b0101001111010111110101011101101100000111000010100010111011010000)  
) LUT6_1196 (
   .O(gates[67]),
   .I0(InputBits[404]),
   .I1(InputBits[520]),
   .I2(InputBits[426]),
   .I3(InputBits[1696]),
   .I4(InputBits[990]),
   .I5(InputBits[1206])
);
LUT6 #(
   .INIT(64'b1010000100101101001000100010010101101000010011001110010001100010)  
) LUT6_1197 (
   .O(gates[812]),
   .I0(InputBits[1441]),
   .I1(InputBits[319]),
   .I2(InputBits[1650]),
   .I3(InputBits[526]),
   .I4(InputBits[248]),
   .I5(InputBits[300])
);
LUT6 #(
   .INIT(64'b1100110000000011101011001100111110101100010100001100010110110011)  
) LUT6_1198 (
   .O(gates[241]),
   .I0(InputBits[967]),
   .I1(InputBits[753]),
   .I2(InputBits[12]),
   .I3(InputBits[896]),
   .I4(InputBits[221]),
   .I5(InputBits[1010])
);
LUT6 #(
   .INIT(64'b1001010111111101010000001001101000110000011010010100001010100000)  
) LUT6_1199 (
   .O(gates[795]),
   .I0(InputBits[603]),
   .I1(InputBits[1492]),
   .I2(InputBits[1021]),
   .I3(InputBits[637]),
   .I4(InputBits[1112]),
   .I5(InputBits[807])
);
LUT6 #(
   .INIT(64'b0011111000010100011001100100111000101101110000110001101101010001)  
) LUT6_1200 (
   .O(gates[489]),
   .I0(InputBits[860]),
   .I1(InputBits[1028]),
   .I2(InputBits[1241]),
   .I3(InputBits[1034]),
   .I4(InputBits[440]),
   .I5(InputBits[46])
);
LUT6 #(
   .INIT(64'b0000011010110010100100111111001101111010011101100001110001011110)  
) LUT6_1201 (
   .O(gates[585]),
   .I0(InputBits[1259]),
   .I1(InputBits[801]),
   .I2(InputBits[101]),
   .I3(InputBits[279]),
   .I4(InputBits[587]),
   .I5(InputBits[655])
);
LUT6 #(
   .INIT(64'b1110110100110110001111000000110111100101100100010000110100000001)  
) LUT6_1202 (
   .O(gates[794]),
   .I0(InputBits[109]),
   .I1(InputBits[1656]),
   .I2(InputBits[1103]),
   .I3(InputBits[1178]),
   .I4(InputBits[912]),
   .I5(InputBits[129])
);
LUT6 #(
   .INIT(64'b0001000101100110000100000110010100111011101001101001100011010101)  
) LUT6_1203 (
   .O(gates[327]),
   .I0(InputBits[1225]),
   .I1(InputBits[771]),
   .I2(InputBits[626]),
   .I3(InputBits[389]),
   .I4(InputBits[1534]),
   .I5(InputBits[674])
);
LUT6 #(
   .INIT(64'b0010011001111000111110011100011110101000110000110000101001100001)  
) LUT6_1204 (
   .O(gates[1392]),
   .I0(InputBits[27]),
   .I1(InputBits[881]),
   .I2(InputBits[1287]),
   .I3(InputBits[44]),
   .I4(InputBits[1458]),
   .I5(InputBits[751])
);
LUT6 #(
   .INIT(64'b0010010000100010101000000101111110100101011001010111010110000010)  
) LUT6_1205 (
   .O(gates[1080]),
   .I0(InputBits[1345]),
   .I1(InputBits[1035]),
   .I2(InputBits[828]),
   .I3(InputBits[1559]),
   .I4(InputBits[1097]),
   .I5(InputBits[782])
);
LUT6 #(
   .INIT(64'b1111111001010100111010100000111001101000010111011001100010001011)  
) LUT6_1206 (
   .O(gates[944]),
   .I0(InputBits[728]),
   .I1(InputBits[1048]),
   .I2(InputBits[688]),
   .I3(InputBits[1131]),
   .I4(InputBits[852]),
   .I5(InputBits[1327])
);
LUT6 #(
   .INIT(64'b0010100111111000011100101010111011001010110000101100101101001000)  
) LUT6_1207 (
   .O(gates[1281]),
   .I0(InputBits[1679]),
   .I1(InputBits[107]),
   .I2(InputBits[544]),
   .I3(InputBits[1140]),
   .I4(InputBits[921]),
   .I5(InputBits[1433])
);
LUT6 #(
   .INIT(64'b0100011100111100001100001000011000010101010011100000010010000010)  
) LUT6_1208 (
   .O(gates[1113]),
   .I0(InputBits[32]),
   .I1(InputBits[366]),
   .I2(InputBits[4]),
   .I3(InputBits[1311]),
   .I4(InputBits[1662]),
   .I5(InputBits[238])
);
LUT6 #(
   .INIT(64'b1111001011100111110010010111010101110110010110000010001000011011)  
) LUT6_1209 (
   .O(gates[732]),
   .I0(InputBits[146]),
   .I1(InputBits[305]),
   .I2(InputBits[561]),
   .I3(InputBits[888]),
   .I4(InputBits[695]),
   .I5(InputBits[458])
);
LUT6 #(
   .INIT(64'b1001011010010011011111111011010000000011010001011001000110111100)  
) LUT6_1210 (
   .O(gates[674]),
   .I0(InputBits[346]),
   .I1(InputBits[382]),
   .I2(InputBits[675]),
   .I3(InputBits[330]),
   .I4(InputBits[1210]),
   .I5(InputBits[1350])
);
LUT6 #(
   .INIT(64'b0000101001111001111110010010101000101011001101001000110111011100)  
) LUT6_1211 (
   .O(gates[1317]),
   .I0(InputBits[262]),
   .I1(InputBits[744]),
   .I2(InputBits[1265]),
   .I3(InputBits[1053]),
   .I4(InputBits[1059]),
   .I5(InputBits[1152])
);
LUT6 #(
   .INIT(64'b1011011101110001110010000101110011110010101111111110111011101001)  
) LUT6_1212 (
   .O(gates[280]),
   .I0(InputBits[1262]),
   .I1(InputBits[1499]),
   .I2(InputBits[1068]),
   .I3(InputBits[694]),
   .I4(InputBits[302]),
   .I5(InputBits[868])
);
LUT6 #(
   .INIT(64'b1011101001000010110110011000001111111001111101101101101111000010)  
) LUT6_1213 (
   .O(gates[957]),
   .I0(InputBits[50]),
   .I1(InputBits[352]),
   .I2(InputBits[876]),
   .I3(InputBits[1615]),
   .I4(InputBits[390]),
   .I5(InputBits[1605])
);
LUT6 #(
   .INIT(64'b0001010010110111110111001000001011110000001010110110111101010111)  
) LUT6_1214 (
   .O(gates[273]),
   .I0(InputBits[1565]),
   .I1(InputBits[1724]),
   .I2(InputBits[766]),
   .I3(InputBits[433]),
   .I4(InputBits[1580]),
   .I5(InputBits[391])
);
LUT6 #(
   .INIT(64'b0010110001011011010100000010011111000000011010110101000101101101)  
) LUT6_1215 (
   .O(gates[471]),
   .I0(InputBits[1527]),
   .I1(InputBits[1465]),
   .I2(InputBits[721]),
   .I3(InputBits[1707]),
   .I4(InputBits[19]),
   .I5(InputBits[24])
);
LUT6 #(
   .INIT(64'b0010010100001101101011001100001000001000011001101010001010100001)  
) LUT6_1216 (
   .O(gates[622]),
   .I0(InputBits[1219]),
   .I1(InputBits[1479]),
   .I2(InputBits[1208]),
   .I3(InputBits[216]),
   .I4(InputBits[1416]),
   .I5(InputBits[1434])
);
LUT6 #(
   .INIT(64'b1011001100111011111000010001001000100111100011110110111010110110)  
) LUT6_1217 (
   .O(gates[1503]),
   .I0(InputBits[1336]),
   .I1(InputBits[854]),
   .I2(InputBits[1278]),
   .I3(InputBits[169]),
   .I4(InputBits[1089]),
   .I5(InputBits[593])
);
LUT6 #(
   .INIT(64'b0011111100010110111000001010111100000001101110010001100100011000)  
) LUT6_1218 (
   .O(gates[970]),
   .I0(InputBits[210]),
   .I1(InputBits[1408]),
   .I2(InputBits[1600]),
   .I3(InputBits[1389]),
   .I4(InputBits[1404]),
   .I5(InputBits[62])
);
LUT6 #(
   .INIT(64'b1000010111010011100001010100000101001100011011100100000011011100)  
) LUT6_1219 (
   .O(gates[1509]),
   .I0(InputBits[1589]),
   .I1(InputBits[1095]),
   .I2(InputBits[288]),
   .I3(InputBits[1725]),
   .I4(InputBits[1370]),
   .I5(InputBits[1435])
);
LUT6 #(
   .INIT(64'b1111111101111101010111001000110100101001111001000010011110101011)  
) LUT6_1220 (
   .O(gates[1416]),
   .I0(InputBits[1071]),
   .I1(InputBits[358]),
   .I2(InputBits[684]),
   .I3(InputBits[1474]),
   .I4(InputBits[1157]),
   .I5(InputBits[837])
);
LUT6 #(
   .INIT(64'b0011111011001110010100101000011001001111001111010001010000001101)  
) LUT6_1221 (
   .O(gates[24]),
   .I0(InputBits[7]),
   .I1(InputBits[324]),
   .I2(InputBits[269]),
   .I3(InputBits[645]),
   .I4(InputBits[726]),
   .I5(InputBits[1362])
);
LUT6 #(
   .INIT(64'b0111011001011000010110010010001011101011111001111010000101000111)  
) LUT6_1222 (
   .O(gates[104]),
   .I0(InputBits[2]),
   .I1(InputBits[314]),
   .I2(InputBits[1635]),
   .I3(InputBits[1502]),
   .I4(InputBits[787]),
   .I5(InputBits[501])
);
LUT6 #(
   .INIT(64'b1100000100111110001100010101000100011000010001010110111100111000)  
) LUT6_1223 (
   .O(gates[1325]),
   .I0(InputBits[749]),
   .I1(InputBits[1321]),
   .I2(InputBits[786]),
   .I3(InputBits[580]),
   .I4(InputBits[1249]),
   .I5(InputBits[1292])
);
LUT6 #(
   .INIT(64'b0111101101011101001000000010011000000110011011110101101000000000)  
) LUT6_1224 (
   .O(gates[131]),
   .I0(InputBits[1678]),
   .I1(InputBits[1460]),
   .I2(InputBits[365]),
   .I3(InputBits[276]),
   .I4(InputBits[910]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0010101001010111100101101111110101100111010110000110000001011011)  
) LUT6_1225 (
   .O(gates[502]),
   .I0(InputBits[1310]),
   .I1(InputBits[143]),
   .I2(InputBits[1227]),
   .I3(InputBits[1437]),
   .I4(InputBits[482]),
   .I5(InputBits[1084])
);
LUT6 #(
   .INIT(64'b1101100001000010110011000111100001101010101001111101110110000001)  
) LUT6_1226 (
   .O(gates[314]),
   .I0(InputBits[900]),
   .I1(InputBits[843]),
   .I2(InputBits[335]),
   .I3(InputBits[126]),
   .I4(InputBits[1087]),
   .I5(InputBits[799])
);
LUT6 #(
   .INIT(64'b0000111011000111100110011000111001110111011110000101110011010011)  
) LUT6_1227 (
   .O(gates[1286]),
   .I0(InputBits[70]),
   .I1(InputBits[281]),
   .I2(InputBits[1431]),
   .I3(InputBits[847]),
   .I4(InputBits[1176]),
   .I5(InputBits[1374])
);
LUT6 #(
   .INIT(64'b0001110011110110110100010011000000110001011000011001001100011001)  
) LUT6_1228 (
   .O(gates[1237]),
   .I0(InputBits[740]),
   .I1(InputBits[898]),
   .I2(InputBits[286]),
   .I3(InputBits[327]),
   .I4(InputBits[1272]),
   .I5(InputBits[1183])
);
LUT6 #(
   .INIT(64'b0101000101101101101110111011101100010110110011101110101111100001)  
) LUT6_1229 (
   .O(gates[1513]),
   .I0(InputBits[1466]),
   .I1(InputBits[1031]),
   .I2(InputBits[1203]),
   .I3(InputBits[1610]),
   .I4(InputBits[978]),
   .I5(InputBits[1215])
);
LUT6 #(
   .INIT(64'b0010001100101010010011100111111011111101001011000010010010000100)  
) LUT6_1230 (
   .O(gates[1502]),
   .I0(InputBits[1086]),
   .I1(InputBits[1115]),
   .I2(InputBits[1532]),
   .I3(InputBits[1452]),
   .I4(InputBits[29]),
   .I5(InputBits[120])
);
LUT6 #(
   .INIT(64'b1010001011011011010001111100110110000100111100100111011000111110)  
) LUT6_1231 (
   .O(gates[1264]),
   .I0(InputBits[22]),
   .I1(InputBits[601]),
   .I2(InputBits[17]),
   .I3(InputBits[1296]),
   .I4(InputBits[1417]),
   .I5(InputBits[1574])
);
LUT6 #(
   .INIT(64'b0101100100101101011001011111110110110010000011011010110011111100)  
) LUT6_1232 (
   .O(gates[355]),
   .I0(InputBits[595]),
   .I1(InputBits[451]),
   .I2(InputBits[690]),
   .I3(InputBits[1623]),
   .I4(InputBits[1280]),
   .I5(InputBits[209])
);
LUT6 #(
   .INIT(64'b0000101000010001010101001101011100000001111010110001000001011010)  
) LUT6_1233 (
   .O(gates[553]),
   .I0(InputBits[1314]),
   .I1(InputBits[575]),
   .I2(InputBits[353]),
   .I3(InputBits[170]),
   .I4(InputBits[34]),
   .I5(InputBits[163])
);
LUT6 #(
   .INIT(64'b0101100011111100000000000001101010100110101000010101010011000011)  
) LUT6_1234 (
   .O(gates[159]),
   .I0(InputBits[995]),
   .I1(InputBits[1237]),
   .I2(InputBits[824]),
   .I3(InputBits[1128]),
   .I4(InputBits[1688]),
   .I5(InputBits[1448])
);
LUT6 #(
   .INIT(64'b1011010110100101101011101010101011111010011111000010101001100111)  
) LUT6_1235 (
   .O(gates[747]),
   .I0(InputBits[1064]),
   .I1(InputBits[464]),
   .I2(InputBits[115]),
   .I3(InputBits[455]),
   .I4(InputBits[1110]),
   .I5(InputBits[1279])
);
LUT6 #(
   .INIT(64'b1101000111110010101111100001011011011000011100000011110010100010)  
) LUT6_1236 (
   .O(gates[1252]),
   .I0(InputBits[57]),
   .I1(InputBits[913]),
   .I2(InputBits[1727]),
   .I3(InputBits[193]),
   .I4(InputBits[572]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1010000010111111101000010111100001110100010100101110011000000111)  
) LUT6_1237 (
   .O(gates[555]),
   .I0(InputBits[628]),
   .I1(InputBits[667]),
   .I2(InputBits[15]),
   .I3(InputBits[1118]),
   .I4(InputBits[345]),
   .I5(InputBits[429])
);
LUT6 #(
   .INIT(64'b1000000011010100111011111010110100101001110001011110100011110111)  
) LUT6_1238 (
   .O(gates[47]),
   .I0(InputBits[1023]),
   .I1(InputBits[116]),
   .I2(InputBits[486]),
   .I3(InputBits[507]),
   .I4(InputBits[1338]),
   .I5(InputBits[1596])
);
LUT6 #(
   .INIT(64'b1101100111111100111001000010101111001111011000000000001101010110)  
) LUT6_1239 (
   .O(gates[1037]),
   .I0(InputBits[1506]),
   .I1(InputBits[1246]),
   .I2(InputBits[8]),
   .I3(InputBits[1536]),
   .I4(InputBits[611]),
   .I5(InputBits[1331])
);
LUT6 #(
   .INIT(64'b0110100101000000000101111000101110101100110111001001110010010000)  
) LUT6_1240 (
   .O(gates[1427]),
   .I0(InputBits[988]),
   .I1(InputBits[245]),
   .I2(InputBits[1266]),
   .I3(InputBits[546]),
   .I4(InputBits[162]),
   .I5(InputBits[1507])
);
LUT6 #(
   .INIT(64'b0111000100111100111110100100000010000000111101101100100011001010)  
) LUT6_1241 (
   .O(gates[1484]),
   .I0(InputBits[1002]),
   .I1(InputBits[1160]),
   .I2(InputBits[550]),
   .I3(InputBits[79]),
   .I4(InputBits[1139]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100110100011100101011100000110000010100100111111110111011111010)  
) LUT6_1242 (
   .O(gates[37]),
   .I0(InputBits[293]),
   .I1(InputBits[621]),
   .I2(InputBits[1236]),
   .I3(InputBits[1159]),
   .I4(InputBits[1102]),
   .I5(InputBits[755])
);
LUT6 #(
   .INIT(64'b0110101111001100111101101100011100010110010101111001010110111011)  
) LUT6_1243 (
   .O(gates[1017]),
   .I0(InputBits[312]),
   .I1(InputBits[940]),
   .I2(InputBits[931]),
   .I3(InputBits[1497]),
   .I4(InputBits[767]),
   .I5(InputBits[883])
);
LUT6 #(
   .INIT(64'b0001001110101000111000110110100011010101100001010010001100011000)  
) LUT6_1244 (
   .O(gates[855]),
   .I0(InputBits[762]),
   .I1(InputBits[1722]),
   .I2(InputBits[68]),
   .I3(InputBits[1691]),
   .I4(InputBits[950]),
   .I5(InputBits[111])
);
LUT6 #(
   .INIT(64'b1100011110110111011000010000111111000011011001011000001001000010)  
) LUT6_1245 (
   .O(gates[270]),
   .I0(InputBits[1381]),
   .I1(InputBits[654]),
   .I2(InputBits[371]),
   .I3(InputBits[469]),
   .I4(InputBits[819]),
   .I5(InputBits[970])
);
LUT6 #(
   .INIT(64'b1001111001010010101100011010010111000101100101000110110010010001)  
) LUT6_1246 (
   .O(gates[195]),
   .I0(InputBits[495]),
   .I1(InputBits[139]),
   .I2(InputBits[343]),
   .I3(InputBits[764]),
   .I4(InputBits[1186]),
   .I5(InputBits[1073])
);
LUT6 #(
   .INIT(64'b1100100001101001101110101010010101110100010010010101001101011011)  
) LUT6_1247 (
   .O(gates[1057]),
   .I0(InputBits[915]),
   .I1(InputBits[232]),
   .I2(InputBits[1217]),
   .I3(InputBits[196]),
   .I4(InputBits[696]),
   .I5(InputBits[582])
);
LUT6 #(
   .INIT(64'b0000101101101110110000000101000101100011001101010010101101111100)  
) LUT6_1248 (
   .O(gates[538]),
   .I0(InputBits[1628]),
   .I1(InputBits[1260]),
   .I2(InputBits[1524]),
   .I3(InputBits[1239]),
   .I4(InputBits[566]),
   .I5(InputBits[421])
);
LUT6 #(
   .INIT(64'b0011001000000010001010010001011010000110010000111111101011011101)  
) LUT6_1249 (
   .O(gates[679]),
   .I0(InputBits[1515]),
   .I1(InputBits[1153]),
   .I2(InputBits[1007]),
   .I3(InputBits[95]),
   .I4(InputBits[1196]),
   .I5(InputBits[1539])
);
LUT6 #(
   .INIT(64'b1001010101110011101101110001110000000101100111001111110110000101)  
) LUT6_1250 (
   .O(gates[680]),
   .I0(InputBits[1234]),
   .I1(InputBits[519]),
   .I2(InputBits[984]),
   .I3(InputBits[1295]),
   .I4(InputBits[992]),
   .I5(InputBits[412])
);
LUT6 #(
   .INIT(64'b0100101110011001011001000001001110111000110011011000010011101111)  
) LUT6_1251 (
   .O(gates[831]),
   .I0(InputBits[1224]),
   .I1(InputBits[1693]),
   .I2(InputBits[1364]),
   .I3(InputBits[1398]),
   .I4(InputBits[584]),
   .I5(InputBits[310])
);
LUT6 #(
   .INIT(64'b1011110010100011111100010101111010010111001111000101000110010010)  
) LUT6_1252 (
   .O(gates[521]),
   .I0(InputBits[228]),
   .I1(InputBits[373]),
   .I2(InputBits[201]),
   .I3(InputBits[700]),
   .I4(InputBits[81]),
   .I5(InputBits[936])
);
LUT6 #(
   .INIT(64'b0000010111011111111100100111000111111101100010011010101110111101)  
) LUT6_1253 (
   .O(gates[1147]),
   .I0(InputBits[504]),
   .I1(InputBits[272]),
   .I2(InputBits[959]),
   .I3(InputBits[811]),
   .I4(InputBits[946]),
   .I5(InputBits[392])
);
LUT6 #(
   .INIT(64'b1010011101100101011101111001011110011110101011000010000001101001)  
) LUT6_1254 (
   .O(gates[1332]),
   .I0(InputBits[1550]),
   .I1(InputBits[441]),
   .I2(InputBits[1356]),
   .I3(InputBits[715]),
   .I4(InputBits[220]),
   .I5(InputBits[863])
);
LUT6 #(
   .INIT(64'b0010101110101100011110001100111110011101100000101011101101000011)  
) LUT6_1255 (
   .O(gates[162]),
   .I0(InputBits[1577]),
   .I1(InputBits[779]),
   .I2(InputBits[975]),
   .I3(InputBits[510]),
   .I4(InputBits[1401]),
   .I5(InputBits[89])
);
LUT6 #(
   .INIT(64'b1100101111101111101010011000000101011111100111111101111000001101)  
) LUT6_1256 (
   .O(gates[1241]),
   .I0(InputBits[1698]),
   .I1(InputBits[834]),
   .I2(InputBits[1009]),
   .I3(InputBits[1690]),
   .I4(InputBits[827]),
   .I5(InputBits[1391])
);
LUT6 #(
   .INIT(64'b1100100100110110001011110101110110010011100101101011111001100001)  
) LUT6_1257 (
   .O(gates[433]),
   .I0(InputBits[1093]),
   .I1(InputBits[1080]),
   .I2(InputBits[175]),
   .I3(InputBits[722]),
   .I4(InputBits[798]),
   .I5(InputBits[296])
);
LUT6 #(
   .INIT(64'b1011111110110110010111000101101101101000000110011100011001110000)  
) LUT6_1258 (
   .O(gates[880]),
   .I0(InputBits[1643]),
   .I1(InputBits[1660]),
   .I2(InputBits[1075]),
   .I3(InputBits[604]),
   .I4(InputBits[1504]),
   .I5(InputBits[818])
);
LUT6 #(
   .INIT(64'b1100011111001010010100111010110100111110011010011111011011111100)  
) LUT6_1259 (
   .O(gates[1441]),
   .I0(InputBits[708]),
   .I1(InputBits[100]),
   .I2(InputBits[388]),
   .I3(InputBits[1708]),
   .I4(InputBits[1318]),
   .I5(InputBits[236])
);
LUT6 #(
   .INIT(64'b1001000111110001001110110111101101001000010000101100011010010001)  
) LUT6_1260 (
   .O(gates[647]),
   .I0(InputBits[87]),
   .I1(InputBits[94]),
   .I2(InputBits[671]),
   .I3(InputBits[1323]),
   .I4(InputBits[625]),
   .I5(InputBits[516])
);
LUT6 #(
   .INIT(64'b0100000001000000110011000110001101101000001111101000010000001000)  
) LUT6_1261 (
   .O(gates[1399]),
   .I0(InputBits[1214]),
   .I1(InputBits[1193]),
   .I2(InputBits[243]),
   .I3(InputBits[980]),
   .I4(InputBits[77]),
   .I5(InputBits[857])
);
LUT6 #(
   .INIT(64'b0111100010010001011011001101110110011101110100101101001010101011)  
) LUT6_1262 (
   .O(gates[1206]),
   .I0(InputBits[132]),
   .I1(InputBits[597]),
   .I2(InputBits[724]),
   .I3(InputBits[278]),
   .I4(InputBits[1587]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1010111011111011001101101110011110111001010101100110100010011001)  
) LUT6_1263 (
   .O(gates[334]),
   .I0(InputBits[1251]),
   .I1(InputBits[1564]),
   .I2(InputBits[1307]),
   .I3(InputBits[9]),
   .I4(InputBits[234]),
   .I5(InputBits[1477])
);
LUT6 #(
   .INIT(64'b0100010111011011110000101100110110100001010011111100010100011010)  
) LUT6_1264 (
   .O(gates[986]),
   .I0(InputBits[685]),
   .I1(InputBits[462]),
   .I2(InputBits[1108]),
   .I3(InputBits[1637]),
   .I4(InputBits[521]),
   .I5(InputBits[1468])
);
LUT6 #(
   .INIT(64'b1100001101100110000101010000000000000000000000001101000000011100)  
) LUT6_1265 (
   .O(gates[786]),
   .I0(InputBits[1329]),
   .I1(InputBits[1106]),
   .I2(InputBits[283]),
   .I3(InputBits[218]),
   .I4(InputBits[1611]),
   .I5(InputBits[1018])
);
LUT6 #(
   .INIT(64'b0011011111001101000110101011111111110110111001011100101010000000)  
) LUT6_1266 (
   .O(gates[1117]),
   .I0(InputBits[1429]),
   .I1(InputBits[1522]),
   .I2(InputBits[1379]),
   .I3(InputBits[1305]),
   .I4(InputBits[102]),
   .I5(InputBits[1586])
);
LUT6 #(
   .INIT(64'b0001100001010100100001111110111101011111110110000100110011011100)  
) LUT6_1267 (
   .O(gates[740]),
   .I0(InputBits[835]),
   .I1(InputBits[1454]),
   .I2(InputBits[630]),
   .I3(InputBits[1162]),
   .I4(InputBits[1025]),
   .I5(InputBits[1572])
);
LUT6 #(
   .INIT(64'b0101011000111000100010001100011000110011101010000111101110000000)  
) LUT6_1268 (
   .O(gates[1008]),
   .I0(InputBits[796]),
   .I1(InputBits[564]),
   .I2(InputBits[198]),
   .I3(InputBits[1632]),
   .I4(InputBits[570]),
   .I5(InputBits[1133])
);
LUT6 #(
   .INIT(64'b0100011100000010111101101001011110110011100100100110111010011110)  
) LUT6_1269 (
   .O(gates[1027]),
   .I0(InputBits[292]),
   .I1(InputBits[998]),
   .I2(InputBits[242]),
   .I3(InputBits[1424]),
   .I4(InputBits[359]),
   .I5(InputBits[1715])
);
LUT6 #(
   .INIT(64'b1010000100110011010010110000111010101111111001100001110011110101)  
) LUT6_1270 (
   .O(gates[103]),
   .I0(InputBits[891]),
   .I1(InputBits[1484]),
   .I2(InputBits[1014]),
   .I3(InputBits[1406]),
   .I4(InputBits[364]),
   .I5(InputBits[1201])
);
LUT6 #(
   .INIT(64'b1011000110111000010110000101110100110101101001101101000110000000)  
) LUT6_1271 (
   .O(gates[201]),
   .I0(InputBits[150]),
   .I1(InputBits[383]),
   .I2(InputBits[1445]),
   .I3(InputBits[540]),
   .I4(InputBits[1672]),
   .I5(InputBits[1046])
);
LUT6 #(
   .INIT(64'b1101011000101101010001010010011111101011111010101110111001011010)  
) LUT6_1272 (
   .O(gates[871]),
   .I0(InputBits[1044]),
   .I1(InputBits[1405]),
   .I2(InputBits[1552]),
   .I3(InputBits[1423]),
   .I4(InputBits[31]),
   .I5(InputBits[1016])
);
LUT6 #(
   .INIT(64'b0001111001100001010000000010111011110000000011111110010010001010)  
) LUT6_1273 (
   .O(gates[1401]),
   .I0(InputBits[431]),
   .I1(InputBits[1302]),
   .I2(InputBits[1051]),
   .I3(InputBits[367]),
   .I4(InputBits[1493]),
   .I5(InputBits[449])
);
LUT6 #(
   .INIT(64'b1100001010010011101000011010101010000100100000000010110101110001)  
) LUT6_1274 (
   .O(gates[423]),
   .I0(InputBits[258]),
   .I1(InputBits[1393]),
   .I2(InputBits[842]),
   .I3(InputBits[505]),
   .I4(InputBits[1074]),
   .I5(InputBits[113])
);
LUT6 #(
   .INIT(64'b0010110010010010111100001101011001111001011000100000111111111101)  
) LUT6_1275 (
   .O(gates[719]),
   .I0(InputBits[160]),
   .I1(InputBits[742]),
   .I2(InputBits[608]),
   .I3(InputBits[659]),
   .I4(InputBits[58]),
   .I5(InputBits[1349])
);
LUT6 #(
   .INIT(64'b1010101100000101111000110010011101011110100001000111001011110110)  
) LUT6_1276 (
   .O(gates[1139]),
   .I0(InputBits[548]),
   .I1(InputBits[1394]),
   .I2(InputBits[791]),
   .I3(InputBits[155]),
   .I4(InputBits[640]),
   .I5(InputBits[669])
);
LUT6 #(
   .INIT(64'b0111011001001110010011011011000100011001101001010000010111000011)  
) LUT6_1277 (
   .O(gates[1319]),
   .I0(InputBits[557]),
   .I1(InputBits[866]),
   .I2(InputBits[350]),
   .I3(InputBits[666]),
   .I4(InputBits[1282]),
   .I5(InputBits[1000])
);
LUT6 #(
   .INIT(64'b0100110001110010010101100000010000111001011000011110011001110101)  
) LUT6_1278 (
   .O(gates[1529]),
   .I0(InputBits[1648]),
   .I1(InputBits[1427]),
   .I2(InputBits[20]),
   .I3(InputBits[257]),
   .I4(InputBits[1681]),
   .I5(InputBits[873])
);
LUT6 #(
   .INIT(64'b1110110010000110000001011110111000111111101011110001111100101010)  
) LUT6_1279 (
   .O(gates[902]),
   .I0(InputBits[386]),
   .I1(InputBits[214]),
   .I2(InputBits[1271]),
   .I3(InputBits[652]),
   .I4(InputBits[920]),
   .I5(InputBits[320])
);
LUT6 #(
   .INIT(64'b0010100101100110010101001010001100110110100110110110100000011100)  
) LUT6_1280 (
   .O(gates[1222]),
   .I0(InputBits[917]),
   .I1(InputBits[118]),
   .I2(InputBits[577]),
   .I3(InputBits[977]),
   .I4(InputBits[1626]),
   .I5(InputBits[318])
);
LUT6 #(
   .INIT(64'b0011010100100110110000100001111001001110100111001011110011001011)  
) LUT6_1281 (
   .O(gates[827]),
   .I0(InputBits[1057]),
   .I1(InputBits[166]),
   .I2(InputBits[942]),
   .I3(InputBits[624]),
   .I4(InputBits[617]),
   .I5(InputBits[476])
);
LUT6 #(
   .INIT(64'b0101001110001101011001101010101111101001000010001010000110100001)  
) LUT6_1282 (
   .O(gates[266]),
   .I0(InputBits[1495]),
   .I1(InputBits[717]),
   .I2(InputBits[334]),
   .I3(InputBits[1137]),
   .I4(InputBits[698]),
   .I5(InputBits[1091])
);
LUT6 #(
   .INIT(64'b1110100111110110011010100111011101001011110010001110011000000110)  
) LUT6_1283 (
   .O(gates[1353]),
   .I0(InputBits[878]),
   .I1(InputBits[41]),
   .I2(InputBits[1232]),
   .I3(InputBits[250]),
   .I4(InputBits[1671]),
   .I5(InputBits[528])
);
LUT6 #(
   .INIT(64'b0000101111110100101011000001110101000101111010100000011111010111)  
) LUT6_1284 (
   .O(gates[174]),
   .I0(InputBits[172]),
   .I1(InputBits[1367]),
   .I2(InputBits[542]),
   .I3(InputBits[1142]),
   .I4(InputBits[1269]),
   .I5(InputBits[96])
);
LUT6 #(
   .INIT(64'b1101111011010001001000011010011001000010000010010101001011101101)  
) LUT6_1285 (
   .O(gates[820]),
   .I0(InputBits[1184]),
   .I1(InputBits[181]),
   .I2(InputBits[14]),
   .I3(InputBits[623]),
   .I4(InputBits[460]),
   .I5(InputBits[1354])
);
LUT6 #(
   .INIT(64'b1000010001000110000111001010110011000011011010100011100000010110)  
) LUT6_1286 (
   .O(gates[422]),
   .I0(InputBits[1653]),
   .I1(InputBits[987]),
   .I2(InputBits[423]),
   .I3(InputBits[568]),
   .I4(InputBits[809]),
   .I5(InputBits[734])
);
LUT6 #(
   .INIT(64'b0010101100110011001110110010001000111000010000110001110111111101)  
) LUT6_1287 (
   .O(gates[905]),
   .I0(InputBits[1005]),
   .I1(InputBits[85]),
   .I2(InputBits[1728]),
   .I3(InputBits[757]),
   .I4(InputBits[1154]),
   .I5(InputBits[1512])
);
LUT6 #(
   .INIT(64'b1111010110011010000110111011110101001101111011111110100011101000)  
) LUT6_1288 (
   .O(gates[1219]),
   .I0(InputBits[1541]),
   .I1(InputBits[1120]),
   .I2(InputBits[1147]),
   .I3(InputBits[1175]),
   .I4(InputBits[1700]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1010110100110100010111100011101010101111011010001110011111010010)  
) LUT6_1289 (
   .O(gates[1194]),
   .I0(InputBits[1038]),
   .I1(InputBits[1641]),
   .I2(InputBits[1575]),
   .I3(InputBits[466]),
   .I4(InputBits[805]),
   .I5(InputBits[340])
);
LUT6 #(
   .INIT(64'b1111001111000111010111001100101011010101000100100011001110011101)  
) LUT6_1290 (
   .O(gates[1552]),
   .I0(InputBits[1365]),
   .I1(InputBits[141]),
   .I2(InputBits[1613]),
   .I3(InputBits[848]),
   .I4(InputBits[483]),
   .I5(InputBits[325])
);
LUT6 #(
   .INIT(64'b0000001101011010101111110011010010000010110011100100011001110001)  
) LUT6_1291 (
   .O(gates[97]),
   .I0(InputBits[1568]),
   .I1(InputBits[706]),
   .I2(InputBits[493]),
   .I3(InputBits[1555]),
   .I4(InputBits[536]),
   .I5(InputBits[443])
);
LUT6 #(
   .INIT(64'b1010001010011011100001100011100000000101101010101010001000011010)  
) LUT6_1292 (
   .O(gates[41]),
   .I0(InputBits[777]),
   .I1(InputBits[416]),
   .I2(InputBits[1375]),
   .I3(InputBits[803]),
   .I4(InputBits[943]),
   .I5(InputBits[394])
);
LUT6 #(
   .INIT(64'b0011101010111000001000110101110111100100111110101011010011111000)  
) LUT6_1293 (
   .O(gates[668]),
   .I0(InputBits[189]),
   .I1(InputBits[692]),
   .I2(InputBits[1619]),
   .I3(InputBits[1562]),
   .I4(InputBits[1312]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0100101111101000100100000110111010110010001001111001100100111111)  
) LUT6_1294 (
   .O(gates[52]),
   .I0(InputBits[1316]),
   .I1(InputBits[308]),
   .I2(InputBits[1720]),
   .I3(InputBits[1358]),
   .I4(InputBits[908]),
   .I5(InputBits[745])
);
LUT6 #(
   .INIT(64'b1100100111100110110000000001101111110001010101010000001000000101)  
) LUT6_1295 (
   .O(gates[688]),
   .I0(InputBits[925]),
   .I1(InputBits[938]),
   .I2(InputBits[92]),
   .I3(InputBits[341]),
   .I4(InputBits[1340]),
   .I5(InputBits[825])
);
LUT6 #(
   .INIT(64'b1111110000010101101111100011100110000000101100111010101010011110)  
) LUT6_1296 (
   .O(gates[750]),
   .I0(InputBits[813]),
   .I1(InputBits[131]),
   .I2(InputBits[400]),
   .I3(InputBits[1710]),
   .I4(InputBits[1222]),
   .I5(InputBits[33])
);
LUT6 #(
   .INIT(64'b0011001111100010010111010000011000010110100111111010101011111001)  
) LUT6_1297 (
   .O(gates[302]),
   .I0(gatesReg[127]),
   .I1(gatesReg[1049]),
   .I2(gatesReg[71]),
   .I3(gatesReg[1481]),
   .I4(gatesReg[882]),
   .I5(gatesReg[1050])
);
LUT6 #(
   .INIT(64'b1011100011001001110110101011101001011011111001110000111011000110)  
) LUT6_1298 (
   .O(gates[1451]),
   .I0(gatesReg[1488]),
   .I1(gatesReg[560]),
   .I2(gatesReg[1178]),
   .I3(gatesReg[898]),
   .I4(gatesReg[798]),
   .I5(gatesReg[1031])
);
LUT6 #(
   .INIT(64'b1001101011000111110100100000011100011011111110010001100000101000)  
) LUT6_1299 (
   .O(gates[1126]),
   .I0(gatesReg[1387]),
   .I1(gatesReg[512]),
   .I2(gatesReg[463]),
   .I3(gatesReg[1273]),
   .I4(gatesReg[517]),
   .I5(gatesReg[458])
);
LUT6 #(
   .INIT(64'b0011010000000101001100100100100000011110100111100100100101100000)  
) LUT6_1300 (
   .O(gates[774]),
   .I0(gatesReg[451]),
   .I1(gatesReg[454]),
   .I2(gatesReg[1364]),
   .I3(gatesReg[1408]),
   .I4(gatesReg[1250]),
   .I5(gatesReg[1363])
);
LUT6 #(
   .INIT(64'b1011001011110100101011100101011010100011000000110011010110111101)  
) LUT6_1301 (
   .O(gates[1453]),
   .I0(gatesReg[722]),
   .I1(gatesReg[634]),
   .I2(gatesReg[1109]),
   .I3(gatesReg[578]),
   .I4(gatesReg[695]),
   .I5(gatesReg[978])
);
LUT6 #(
   .INIT(64'b0000001000101100101110101001111100110011110011000011100111011011)  
) LUT6_1302 (
   .O(gates[866]),
   .I0(gatesReg[728]),
   .I1(gatesReg[1244]),
   .I2(gatesReg[742]),
   .I3(gatesReg[325]),
   .I4(gatesReg[378]),
   .I5(gatesReg[29])
);
LUT6 #(
   .INIT(64'b0000100000001110110101101001111001010100101010100110011101001001)  
) LUT6_1303 (
   .O(gates[910]),
   .I0(gatesReg[889]),
   .I1(gatesReg[350]),
   .I2(gatesReg[1233]),
   .I3(gatesReg[540]),
   .I4(gatesReg[58]),
   .I5(gatesReg[1162])
);
LUT6 #(
   .INIT(64'b0111011011000111011110000000101110111001110010101010111000011111)  
) LUT6_1304 (
   .O(gates[1341]),
   .I0(gatesReg[153]),
   .I1(gatesReg[684]),
   .I2(gatesReg[211]),
   .I3(gatesReg[861]),
   .I4(gatesReg[337]),
   .I5(gatesReg[101])
);
LUT6 #(
   .INIT(64'b1000000011010101000011000000110110111010101000110100000101011100)  
) LUT6_1305 (
   .O(gates[693]),
   .I0(gatesReg[1546]),
   .I1(gatesReg[340]),
   .I2(gatesReg[76]),
   .I3(gatesReg[311]),
   .I4(gatesReg[982]),
   .I5(gatesReg[571])
);
LUT6 #(
   .INIT(64'b1011011001111110101000110000010100001100011010100010110011010000)  
) LUT6_1306 (
   .O(gates[770]),
   .I0(gatesReg[1214]),
   .I1(gatesReg[1190]),
   .I2(gatesReg[825]),
   .I3(gatesReg[389]),
   .I4(gatesReg[917]),
   .I5(gatesReg[495])
);
LUT6 #(
   .INIT(64'b0111000000110000010001111111100011011000101000111000110100011101)  
) LUT6_1307 (
   .O(gates[593]),
   .I0(gatesReg[1345]),
   .I1(gatesReg[1171]),
   .I2(gatesReg[966]),
   .I3(gatesReg[1123]),
   .I4(gatesReg[1322]),
   .I5(gatesReg[992])
);
LUT6 #(
   .INIT(64'b1001001111111001100011001110001001100101110011010000001010110101)  
) LUT6_1308 (
   .O(gates[188]),
   .I0(gatesReg[758]),
   .I1(gatesReg[236]),
   .I2(gatesReg[706]),
   .I3(gatesReg[218]),
   .I4(gatesReg[1172]),
   .I5(gatesReg[14])
);
LUT6 #(
   .INIT(64'b0111001000111000101011011001010011010000111100000010000110000001)  
) LUT6_1309 (
   .O(gates[402]),
   .I0(gatesReg[1259]),
   .I1(gatesReg[834]),
   .I2(gatesReg[285]),
   .I3(gatesReg[234]),
   .I4(gatesReg[594]),
   .I5(gatesReg[1216])
);
LUT6 #(
   .INIT(64'b1101111110110100011000110010110000000011110110001000100010010001)  
) LUT6_1310 (
   .O(gates[1534]),
   .I0(gatesReg[1438]),
   .I1(gatesReg[1135]),
   .I2(gatesReg[1203]),
   .I3(gatesReg[96]),
   .I4(gatesReg[1068]),
   .I5(gatesReg[486])
);
LUT6 #(
   .INIT(64'b0011000111011101011110111110000010100010000010011110000101110110)  
) LUT6_1311 (
   .O(gates[641]),
   .I0(gatesReg[1354]),
   .I1(gatesReg[160]),
   .I2(gatesReg[569]),
   .I3(gatesReg[8]),
   .I4(gatesReg[98]),
   .I5(gatesReg[1278])
);
LUT6 #(
   .INIT(64'b0001100000100111011000010000100011000010011101100100000110001101)  
) LUT6_1312 (
   .O(gates[1097]),
   .I0(gatesReg[1048]),
   .I1(gatesReg[1000]),
   .I2(gatesReg[1381]),
   .I3(gatesReg[1061]),
   .I4(gatesReg[43]),
   .I5(gatesReg[686])
);
LUT6 #(
   .INIT(64'b1000111001011100000101001101100010010000101101010000010101011010)  
) LUT6_1313 (
   .O(gates[893]),
   .I0(gatesReg[1396]),
   .I1(gatesReg[391]),
   .I2(gatesReg[193]),
   .I3(gatesReg[943]),
   .I4(gatesReg[288]),
   .I5(gatesReg[1555])
);
LUT6 #(
   .INIT(64'b0010010100000111101010110001100000000001001010100101101100000101)  
) LUT6_1314 (
   .O(gates[838]),
   .I0(gatesReg[119]),
   .I1(gatesReg[586]),
   .I2(gatesReg[180]),
   .I3(gatesReg[1375]),
   .I4(gatesReg[410]),
   .I5(gatesReg[246])
);
LUT6 #(
   .INIT(64'b0001001100101111110111000000010010100010000011011101100100011110)  
) LUT6_1315 (
   .O(gates[616]),
   .I0(gatesReg[690]),
   .I1(gatesReg[999]),
   .I2(gatesReg[61]),
   .I3(gatesReg[1168]),
   .I4(gatesReg[1180]),
   .I5(gatesReg[1185])
);
LUT6 #(
   .INIT(64'b0110001010110101000110011000110000110111101101100000010011001010)  
) LUT6_1316 (
   .O(gates[640]),
   .I0(gatesReg[430]),
   .I1(gatesReg[447]),
   .I2(gatesReg[1446]),
   .I3(gatesReg[536]),
   .I4(gatesReg[1130]),
   .I5(gatesReg[1315])
);
LUT6 #(
   .INIT(64'b0011100111110001111100001111000010110111100111010011100010010110)  
) LUT6_1317 (
   .O(gates[1121]),
   .I0(gatesReg[415]),
   .I1(gatesReg[1266]),
   .I2(gatesReg[189]),
   .I3(gatesReg[1292]),
   .I4(gatesReg[1356]),
   .I5(gatesReg[480])
);
LUT6 #(
   .INIT(64'b1010011011011110011011111000101000101111110110010010000101010001)  
) LUT6_1318 (
   .O(gates[870]),
   .I0(gatesReg[438]),
   .I1(gatesReg[1153]),
   .I2(gatesReg[107]),
   .I3(gatesReg[87]),
   .I4(gatesReg[1022]),
   .I5(gatesReg[1458])
);
LUT6 #(
   .INIT(64'b0001100101101011001111000010110100101100011111110010111111000010)  
) LUT6_1319 (
   .O(gates[804]),
   .I0(gatesReg[444]),
   .I1(gatesReg[508]),
   .I2(gatesReg[953]),
   .I3(gatesReg[1336]),
   .I4(gatesReg[221]),
   .I5(gatesReg[39])
);
LUT6 #(
   .INIT(64'b0111110100111100011101110101110011100001110011011011000011111100)  
) LUT6_1320 (
   .O(gates[83]),
   .I0(gatesReg[1424]),
   .I1(gatesReg[1089]),
   .I2(gatesReg[558]),
   .I3(gatesReg[417]),
   .I4(gatesReg[12]),
   .I5(gatesReg[1554])
);
LUT6 #(
   .INIT(64'b0000100011111101100100011001110101111010001010111100010101001111)  
) LUT6_1321 (
   .O(gates[1384]),
   .I0(gatesReg[784]),
   .I1(gatesReg[260]),
   .I2(gatesReg[573]),
   .I3(gatesReg[1084]),
   .I4(gatesReg[1530]),
   .I5(gatesReg[762])
);
LUT6 #(
   .INIT(64'b0010110100110100100101011110111010001111101010111100000010001101)  
) LUT6_1322 (
   .O(gates[896]),
   .I0(gatesReg[1144]),
   .I1(gatesReg[638]),
   .I2(gatesReg[734]),
   .I3(gatesReg[875]),
   .I4(gatesReg[1522]),
   .I5(gatesReg[1])
);
LUT6 #(
   .INIT(64'b0001011110110111101101100011100010100010101000001011010011111100)  
) LUT6_1323 (
   .O(gates[1468]),
   .I0(gatesReg[506]),
   .I1(gatesReg[136]),
   .I2(gatesReg[116]),
   .I3(gatesReg[1197]),
   .I4(gatesReg[144]),
   .I5(gatesReg[661])
);
LUT6 #(
   .INIT(64'b1011001110001011001111001010100101001100111111011001101010101010)  
) LUT6_1324 (
   .O(gates[1385]),
   .I0(gatesReg[1440]),
   .I1(gatesReg[381]),
   .I2(gatesReg[1471]),
   .I3(gatesReg[581]),
   .I4(gatesReg[308]),
   .I5(gatesReg[906])
);
LUT6 #(
   .INIT(64'b0011111101110011000110000011001000000010001010000111101101010100)  
) LUT6_1325 (
   .O(gates[1464]),
   .I0(gatesReg[1349]),
   .I1(gatesReg[177]),
   .I2(gatesReg[678]),
   .I3(gatesReg[1517]),
   .I4(gatesReg[373]),
   .I5(gatesReg[773])
);
LUT6 #(
   .INIT(64'b1111100011010011111001101110000010001110100111011111101110110101)  
) LUT6_1326 (
   .O(gates[1494]),
   .I0(gatesReg[1247]),
   .I1(gatesReg[205]),
   .I2(gatesReg[22]),
   .I3(gatesReg[927]),
   .I4(gatesReg[1309]),
   .I5(gatesReg[301])
);
LUT6 #(
   .INIT(64'b1011100010100100001110000001001101011000111100111100111111101000)  
) LUT6_1327 (
   .O(gates[962]),
   .I0(gatesReg[51]),
   .I1(gatesReg[1260]),
   .I2(gatesReg[456]),
   .I3(gatesReg[652]),
   .I4(gatesReg[874]),
   .I5(gatesReg[975])
);
LUT6 #(
   .INIT(64'b0100010101100110010111010001001001110011010111111001101100011110)  
) LUT6_1328 (
   .O(gates[1085]),
   .I0(gatesReg[493]),
   .I1(gatesReg[1033]),
   .I2(gatesReg[1436]),
   .I3(gatesReg[1539]),
   .I4(gatesReg[1320]),
   .I5(gatesReg[796])
);
LUT6 #(
   .INIT(64'b0010000011110011011001100111001000000110011001010001011101010101)  
) LUT6_1329 (
   .O(gates[755]),
   .I0(gatesReg[1026]),
   .I1(gatesReg[366]),
   .I2(gatesReg[844]),
   .I3(gatesReg[1541]),
   .I4(gatesReg[1390]),
   .I5(gatesReg[272])
);
LUT6 #(
   .INIT(64'b0011011111110100110111001001000011010010001100011110000100010001)  
) LUT6_1330 (
   .O(gates[777]),
   .I0(gatesReg[775]),
   .I1(gatesReg[1469]),
   .I2(gatesReg[1499]),
   .I3(gatesReg[746]),
   .I4(gatesReg[400]),
   .I5(gatesReg[534])
);
LUT6 #(
   .INIT(64'b0110000011010000101000110110011011100100011111000001001101101101)  
) LUT6_1331 (
   .O(gates[143]),
   .I0(gatesReg[919]),
   .I1(gatesReg[744]),
   .I2(gatesReg[1268]),
   .I3(gatesReg[20]),
   .I4(gatesReg[888]),
   .I5(gatesReg[633])
);
LUT6 #(
   .INIT(64'b1001111101000101010011110000101100101000011000100111001001000110)  
) LUT6_1332 (
   .O(gates[464]),
   .I0(gatesReg[1372]),
   .I1(gatesReg[1011]),
   .I2(gatesReg[151]),
   .I3(gatesReg[468]),
   .I4(gatesReg[1161]),
   .I5(gatesReg[1285])
);
LUT6 #(
   .INIT(64'b0100101000011011011011001101000000101000011001111110110100001110)  
) LUT6_1333 (
   .O(gates[1403]),
   .I0(gatesReg[1019]),
   .I1(gatesReg[700]),
   .I2(gatesReg[287]),
   .I3(gatesReg[78]),
   .I4(gatesReg[475]),
   .I5(gatesReg[1380])
);
LUT6 #(
   .INIT(64'b0010000110101011101001111011101111000001110010100000000010011111)  
) LUT6_1334 (
   .O(gates[6]),
   .I0(gatesReg[413]),
   .I1(gatesReg[990]),
   .I2(gatesReg[294]),
   .I3(gatesReg[349]),
   .I4(gatesReg[932]),
   .I5(gatesReg[1442])
);
LUT6 #(
   .INIT(64'b0111111110000000011010100010001101011001100111000001101000011111)  
) LUT6_1335 (
   .O(gates[1051]),
   .I0(gatesReg[764]),
   .I1(gatesReg[1549]),
   .I2(gatesReg[1525]),
   .I3(gatesReg[515]),
   .I4(gatesReg[1242]),
   .I5(gatesReg[1107])
);
LUT6 #(
   .INIT(64'b1101001100011101110101100100000011100010100110001101000100011111)  
) LUT6_1336 (
   .O(gates[562]),
   .I0(gatesReg[1208]),
   .I1(gatesReg[138]),
   .I2(gatesReg[606]),
   .I3(gatesReg[1383]),
   .I4(gatesReg[137]),
   .I5(gatesReg[1414])
);
LUT6 #(
   .INIT(64'b1111010111001000111010100110011010101110110110010101011000110110)  
) LUT6_1337 (
   .O(gates[1497]),
   .I0(gatesReg[724]),
   .I1(gatesReg[1201]),
   .I2(gatesReg[432]),
   .I3(gatesReg[666]),
   .I4(gatesReg[519]),
   .I5(gatesReg[1074])
);
LUT6 #(
   .INIT(64'b1010011100010010101010011000101101011001011100011011000100110000)  
) LUT6_1338 (
   .O(gates[1304]),
   .I0(gatesReg[860]),
   .I1(gatesReg[1195]),
   .I2(gatesReg[1063]),
   .I3(gatesReg[17]),
   .I4(gatesReg[1327]),
   .I5(gatesReg[1274])
);
LUT6 #(
   .INIT(64'b0110011110001011100110111011010110001011010011100111110001000110)  
) LUT6_1339 (
   .O(gates[183]),
   .I0(gatesReg[708]),
   .I1(gatesReg[110]),
   .I2(gatesReg[333]),
   .I3(gatesReg[710]),
   .I4(gatesReg[323]),
   .I5(gatesReg[856])
);
LUT6 #(
   .INIT(64'b1111100110101110111101000100001000000001011011010110111001110000)  
) LUT6_1340 (
   .O(gates[497]),
   .I0(gatesReg[112]),
   .I1(gatesReg[545]),
   .I2(gatesReg[191]),
   .I3(gatesReg[187]),
   .I4(gatesReg[588]),
   .I5(gatesReg[646])
);
LUT6 #(
   .INIT(64'b1100111101011101010110000011011110001111001100110101101000000010)  
) LUT6_1341 (
   .O(gates[1102]),
   .I0(gatesReg[756]),
   .I1(gatesReg[446]),
   .I2(gatesReg[262]),
   .I3(gatesReg[1283]),
   .I4(gatesReg[1220]),
   .I5(gatesReg[212])
);
LUT6 #(
   .INIT(64'b0010100011000010110010010010111101101110010011111111101011101110)  
) LUT6_1342 (
   .O(gates[518]),
   .I0(gatesReg[1331]),
   .I1(gatesReg[1149]),
   .I2(gatesReg[542]),
   .I3(gatesReg[1305]),
   .I4(gatesReg[961]),
   .I5(gatesReg[1288])
);
LUT6 #(
   .INIT(64'b1100100100110001000110000100111110100100010011001111001001101110)  
) LUT6_1343 (
   .O(gates[1478]),
   .I0(gatesReg[1087]),
   .I1(gatesReg[810]),
   .I2(gatesReg[574]),
   .I3(gatesReg[1238]),
   .I4(gatesReg[170]),
   .I5(gatesReg[33])
);
LUT6 #(
   .INIT(64'b1110001110001111000011000101101001001110101000110101111101101100)  
) LUT6_1344 (
   .O(gates[439]),
   .I0(gatesReg[660]),
   .I1(gatesReg[7]),
   .I2(gatesReg[227]),
   .I3(gatesReg[26]),
   .I4(gatesReg[977]),
   .I5(gatesReg[566])
);
LUT6 #(
   .INIT(64'b0110010101010011101111111011011001000111011011111001111101001110)  
) LUT6_1345 (
   .O(gates[1211]),
   .I0(gatesReg[526]),
   .I1(gatesReg[806]),
   .I2(gatesReg[264]),
   .I3(gatesReg[255]),
   .I4(gatesReg[359]),
   .I5(gatesReg[182])
);
LUT6 #(
   .INIT(64'b1010110110110110101101010000001011111010111111001010100010000001)  
) LUT6_1346 (
   .O(gates[362]),
   .I0(gatesReg[1229]),
   .I1(gatesReg[108]),
   .I2(gatesReg[604]),
   .I3(gatesReg[1001]),
   .I4(gatesReg[556]),
   .I5(gatesReg[717])
);
LUT6 #(
   .INIT(64'b1100101010100010110011101110000100001001000010011101010100110000)  
) LUT6_1347 (
   .O(gates[1379]),
   .I0(gatesReg[232]),
   .I1(gatesReg[477]),
   .I2(gatesReg[815]),
   .I3(gatesReg[671]),
   .I4(gatesReg[1338]),
   .I5(gatesReg[1511])
);
LUT6 #(
   .INIT(64'b0011110101101011001101000100111011110101110000010001101110101101)  
) LUT6_1348 (
   .O(gates[169]),
   .I0(gatesReg[1182]),
   .I1(gatesReg[225]),
   .I2(gatesReg[330]),
   .I3(gatesReg[142]),
   .I4(gatesReg[1447]),
   .I5(gatesReg[207])
);
LUT6 #(
   .INIT(64'b1110100000011010100110111111110101010010110111101001110001010010)  
) LUT6_1349 (
   .O(gates[411]),
   .I0(gatesReg[1510]),
   .I1(gatesReg[167]),
   .I2(gatesReg[48]),
   .I3(gatesReg[360]),
   .I4(gatesReg[692]),
   .I5(gatesReg[663])
);
LUT6 #(
   .INIT(64'b0001000101101100100010001001010010011100111100010110000010100101)  
) LUT6_1350 (
   .O(gates[1542]),
   .I0(gatesReg[854]),
   .I1(gatesReg[969]),
   .I2(gatesReg[1174]),
   .I3(gatesReg[1076]),
   .I4(gatesReg[510]),
   .I5(gatesReg[766])
);
LUT6 #(
   .INIT(64'b1001010101111001111001011100101111110111000110001101000011001110)  
) LUT6_1351 (
   .O(gates[705]),
   .I0(gatesReg[393]),
   .I1(gatesReg[449]),
   .I2(gatesReg[1501]),
   .I3(gatesReg[658]),
   .I4(gatesReg[274]),
   .I5(gatesReg[549])
);
LUT6 #(
   .INIT(64'b0001001000001011100110010100011010101111001110110111101100111011)  
) LUT6_1352 (
   .O(gates[478]),
   .I0(gatesReg[659]),
   .I1(gatesReg[877]),
   .I2(gatesReg[1508]),
   .I3(gatesReg[1141]),
   .I4(gatesReg[1128]),
   .I5(gatesReg[682])
);
LUT6 #(
   .INIT(64'b1001110101111100100010000000010100111011010101111100000000000001)  
) LUT6_1353 (
   .O(gates[398]),
   .I0(gatesReg[353]),
   .I1(gatesReg[375]),
   .I2(gatesReg[984]),
   .I3(gatesReg[1155]),
   .I4(gatesReg[946]),
   .I5(gatesReg[1485])
);
LUT6 #(
   .INIT(64'b1011010110100000111101101110000000001011100100110111100011000010)  
) LUT6_1354 (
   .O(gates[384]),
   .I0(gatesReg[788]),
   .I1(gatesReg[128]),
   .I2(gatesReg[1520]),
   .I3(gatesReg[303]),
   .I4(gatesReg[250]),
   .I5(gatesReg[1361])
);
LUT6 #(
   .INIT(64'b1111101010000000100101001011001011101101011001000011011101011011)  
) LUT6_1355 (
   .O(gates[836]),
   .I0(gatesReg[614]),
   .I1(gatesReg[501]),
   .I2(gatesReg[1313]),
   .I3(gatesReg[278]),
   .I4(gatesReg[490]),
   .I5(gatesReg[155])
);
LUT6 #(
   .INIT(64'b0111111001001010010101101000110111101111001101001100001001001010)  
) LUT6_1356 (
   .O(gates[942]),
   .I0(gatesReg[130]),
   .I1(gatesReg[53]),
   .I2(gatesReg[387]),
   .I3(gatesReg[1373]),
   .I4(gatesReg[1465]),
   .I5(gatesReg[1302])
);
LUT6 #(
   .INIT(64'b0110101010011000011001100001110111011001010011100010011111000010)  
) LUT6_1357 (
   .O(gates[955]),
   .I0(gatesReg[1112]),
   .I1(gatesReg[626]),
   .I2(gatesReg[1397]),
   .I3(gatesReg[1294]),
   .I4(gatesReg[941]),
   .I5(gatesReg[461])
);
LUT6 #(
   .INIT(64'b1001111000011110100010111011000110111010011110111111110110100110)  
) LUT6_1358 (
   .O(gates[1376]),
   .I0(gatesReg[583]),
   .I1(gatesReg[1426]),
   .I2(gatesReg[257]),
   .I3(gatesReg[1358]),
   .I4(gatesReg[782]),
   .I5(gatesReg[951])
);
LUT6 #(
   .INIT(64'b1001100001000011100100000010010100001001100011101110100101010110)  
) LUT6_1359 (
   .O(gates[407]),
   .I0(gatesReg[85]),
   .I1(gatesReg[809]),
   .I2(gatesReg[1156]),
   .I3(gatesReg[425]),
   .I4(gatesReg[1486]),
   .I5(gatesReg[591])
);
LUT6 #(
   .INIT(64'b1011100110011010111110110100101010101101011110101110000110010000)  
) LUT6_1360 (
   .O(gates[18]),
   .I0(gatesReg[832]),
   .I1(gatesReg[736]),
   .I2(gatesReg[539]),
   .I3(gatesReg[781]),
   .I4(gatesReg[828]),
   .I5(gatesReg[276])
);
LUT6 #(
   .INIT(64'b1100101001110010110001101010000110110110000010011111110000110110)  
) LUT6_1361 (
   .O(gates[376]),
   .I0(gatesReg[102]),
   .I1(gatesReg[520]),
   .I2(gatesReg[532]),
   .I3(gatesReg[1218]),
   .I4(gatesReg[1193]),
   .I5(gatesReg[55])
);
LUT6 #(
   .INIT(64'b1001111011010111011011110100010010110001100101110111100101110101)  
) LUT6_1362 (
   .O(gates[912]),
   .I0(gatesReg[1404]),
   .I1(gatesReg[1543]),
   .I2(gatesReg[57]),
   .I3(gatesReg[259]),
   .I4(gatesReg[424]),
   .I5(gatesReg[872])
);
LUT6 #(
   .INIT(64'b1000111011000011101000100100100110000110111110100101010001101010)  
) LUT6_1363 (
   .O(gates[785]),
   .I0(gatesReg[163]),
   .I1(gatesReg[1106]),
   .I2(gatesReg[1402]),
   .I3(gatesReg[395]),
   .I4(gatesReg[1146]),
   .I5(gatesReg[89])
);
LUT6 #(
   .INIT(64'b1100100111011011101010000010011110111111001100100111100101000111)  
) LUT6_1364 (
   .O(gates[1432]),
   .I0(gatesReg[175]),
   .I1(gatesReg[1531]),
   .I2(gatesReg[584]),
   .I3(gatesReg[988]),
   .I4(gatesReg[35]),
   .I5(gatesReg[1550])
);
LUT6 #(
   .INIT(64'b0010101001001010011010001010001010001100000010011001011110101010)  
) LUT6_1365 (
   .O(gates[599]),
   .I0(gatesReg[1421]),
   .I1(gatesReg[1454]),
   .I2(gatesReg[347]),
   .I3(gatesReg[1333]),
   .I4(gatesReg[665]),
   .I5(gatesReg[434])
);
LUT6 #(
   .INIT(64'b1111011010100110010010111010100101000001011000110111010110110011)  
) LUT6_1366 (
   .O(gates[1167]),
   .I0(gatesReg[1184]),
   .I1(gatesReg[1476]),
   .I2(gatesReg[865]),
   .I3(gatesReg[1207]),
   .I4(gatesReg[904]),
   .I5(gatesReg[442])
);
LUT6 #(
   .INIT(64'b0100100000000101011111110110000111110101100110000100000001110100)  
) LUT6_1367 (
   .O(gates[587]),
   .I0(gatesReg[930]),
   .I1(gatesReg[649]),
   .I2(gatesReg[689]),
   .I3(gatesReg[886]),
   .I4(gatesReg[1318]),
   .I5(gatesReg[642])
);
LUT6 #(
   .INIT(64'b0001101010010110101111111000110111101000011010000110000011101110)  
) LUT6_1368 (
   .O(gates[1393]),
   .I0(gatesReg[648]),
   .I1(gatesReg[1116]),
   .I2(gatesReg[1329]),
   .I3(gatesReg[1028]),
   .I4(gatesReg[198]),
   .I5(gatesReg[1098])
);
LUT6 #(
   .INIT(64'b0101101110010010001110011111011010111101110101011010000110011001)  
) LUT6_1369 (
   .O(gates[609]),
   .I0(gatesReg[1059]),
   .I1(gatesReg[727]),
   .I2(gatesReg[939]),
   .I3(gatesReg[320]),
   .I4(gatesReg[811]),
   .I5(gatesReg[913])
);
LUT6 #(
   .INIT(64'b0001111111110000110111011001011100101001000010000011111101000000)  
) LUT6_1370 (
   .O(gates[1235]),
   .I0(gatesReg[202]),
   .I1(gatesReg[249]),
   .I2(gatesReg[465]),
   .I3(gatesReg[361]),
   .I4(gatesReg[184]),
   .I5(gatesReg[819])
);
LUT6 #(
   .INIT(64'b0111001010010011101101011001100100011000101010001110011110100000)  
) LUT6_1371 (
   .O(gates[190]),
   .I0(gatesReg[1177]),
   .I1(gatesReg[1189]),
   .I2(gatesReg[776]),
   .I3(gatesReg[1127]),
   .I4(gatesReg[1537]),
   .I5(gatesReg[894])
);
LUT6 #(
   .INIT(64'b0011010011110000010010001010011001100111101000101110110010100111)  
) LUT6_1372 (
   .O(gates[95]),
   .I0(gatesReg[858]),
   .I1(gatesReg[1298]),
   .I2(gatesReg[140]),
   .I3(gatesReg[1459]),
   .I4(gatesReg[1269]),
   .I5(gatesReg[181])
);
LUT6 #(
   .INIT(64'b0001001111101001110001010101000000000010001001011000011001110110)  
) LUT6_1373 (
   .O(gates[298]),
   .I0(gatesReg[412]),
   .I1(gatesReg[954]),
   .I2(gatesReg[385]),
   .I3(gatesReg[1479]),
   .I4(gatesReg[1359]),
   .I5(gatesReg[307])
);
LUT6 #(
   .INIT(64'b0100010101100000000000110111110111001100010001001011101011111101)  
) LUT6_1374 (
   .O(gates[923]),
   .I0(gatesReg[801]),
   .I1(gatesReg[985]),
   .I2(gatesReg[1463]),
   .I3(gatesReg[154]),
   .I4(gatesReg[830]),
   .I5(gatesReg[971])
);
LUT6 #(
   .INIT(64'b1100100001101000011100100011000111100001101100100101010100110011)  
) LUT6_1375 (
   .O(gates[601]),
   .I0(gatesReg[1467]),
   .I1(gatesReg[754]),
   .I2(gatesReg[479]),
   .I3(gatesReg[847]),
   .I4(gatesReg[1101]),
   .I5(gatesReg[1166])
);
LUT6 #(
   .INIT(64'b1011011011001001001000010100010110000100111011011001010000110110)  
) LUT6_1376 (
   .O(gates[822]),
   .I0(gatesReg[704]),
   .I1(gatesReg[326]),
   .I2(gatesReg[1378]),
   .I3(gatesReg[1003]),
   .I4(gatesReg[1462]),
   .I5(gatesReg[1165])
);
LUT6 #(
   .INIT(64'b0010100110001111110001101101001001100001011000101110101010101000)  
) LUT6_1377 (
   .O(gates[231]),
   .I0(gatesReg[1054]),
   .I1(gatesReg[681]),
   .I2(gatesReg[619]),
   .I3(gatesReg[335]),
   .I4(gatesReg[1029]),
   .I5(gatesReg[5])
);
LUT6 #(
   .INIT(64'b1011111000011110100000000111101001010111001110000110000010011011)  
) LUT6_1378 (
   .O(gates[243]),
   .I0(gatesReg[698]),
   .I1(gatesReg[621]),
   .I2(gatesReg[524]),
   .I3(gatesReg[554]),
   .I4(gatesReg[552]),
   .I5(gatesReg[598])
);
LUT6 #(
   .INIT(64'b1010111000101000010011011101001001011100010111111010011010001010)  
) LUT6_1379 (
   .O(gates[779]),
   .I0(gatesReg[780]),
   .I1(gatesReg[1433]),
   .I2(gatesReg[74]),
   .I3(gatesReg[240]),
   .I4(gatesReg[890]),
   .I5(gatesReg[440])
);
LUT6 #(
   .INIT(64'b1110001110101010010110000111110100000101111110001101110011110001)  
) LUT6_1380 (
   .O(gates[551]),
   .I0(gatesReg[230]),
   .I1(gatesReg[115]),
   .I2(gatesReg[1289]),
   .I3(gatesReg[299]),
   .I4(gatesReg[377]),
   .I5(gatesReg[1282])
);
LUT6 #(
   .INIT(64'b0111001011001100110000101010011001100011111000001000101001110011)  
) LUT6_1381 (
   .O(gates[148]),
   .I0(gatesReg[922]),
   .I1(gatesReg[602]),
   .I2(gatesReg[841]),
   .I3(gatesReg[1311]),
   .I4(gatesReg[1044]),
   .I5(gatesReg[1072])
);
LUT6 #(
   .INIT(64'b1110110010010110100000110110000000111111001111000010001110001110)  
) LUT6_1382 (
   .O(gates[343]),
   .I0(gatesReg[1394]),
   .I1(gatesReg[612]),
   .I2(gatesReg[1350]),
   .I3(gatesReg[936]),
   .I4(gatesReg[1391]),
   .I5(gatesReg[1277])
);
LUT6 #(
   .INIT(64'b1100001110110110100110111010101010111110001111111100111101000010)  
) LUT6_1383 (
   .O(gates[504]),
   .I0(gatesReg[91]),
   .I1(gatesReg[1086]),
   .I2(gatesReg[1240]),
   .I3(gatesReg[467]),
   .I4(gatesReg[701]),
   .I5(gatesReg[474])
);
LUT6 #(
   .INIT(64'b0110111110011110101110000000011101010001011101100011001110101011)  
) LUT6_1384 (
   .O(gates[753]),
   .I0(gatesReg[481]),
   .I1(gatesReg[867]),
   .I2(gatesReg[214]),
   .I3(gatesReg[564]),
   .I4(gatesReg[817]),
   .I5(gatesReg[563])
);
LUT6 #(
   .INIT(64'b1011010111111000100110000001110011111010011011001110101110001110)  
) LUT6_1385 (
   .O(gates[1343]),
   .I0(gatesReg[731]),
   .I1(gatesReg[657]),
   .I2(gatesReg[229]),
   .I3(gatesReg[768]),
   .I4(gatesReg[1092]),
   .I5(gatesReg[673])
);
LUT6 #(
   .INIT(64'b0011011100111011011000111010101011001001000110001101010111010011)  
) LUT6_1386 (
   .O(gates[697]),
   .I0(gatesReg[503]),
   .I1(gatesReg[68]),
   .I2(gatesReg[1483]),
   .I3(gatesReg[315]),
   .I4(gatesReg[338]),
   .I5(gatesReg[1347])
);
LUT6 #(
   .INIT(64'b1010001001100111111001010101011001000111001000101001110010011111)  
) LUT6_1387 (
   .O(gates[981]),
   .I0(gatesReg[576]),
   .I1(gatesReg[761]),
   .I2(gatesReg[222]),
   .I3(gatesReg[1504]),
   .I4(gatesReg[25]),
   .I5(gatesReg[738])
);
LUT6 #(
   .INIT(64'b0011101101101110111000110111001011000101110100000001111001101100)  
) LUT6_1388 (
   .O(gates[726]),
   .I0(gatesReg[1415]),
   .I1(gatesReg[484]),
   .I2(gatesReg[1036]),
   .I3(gatesReg[1078]),
   .I4(gatesReg[1243]),
   .I5(gatesReg[305])
);
LUT6 #(
   .INIT(64'b1001111010110010101100001001001000110111001110001111111110001111)  
) LUT6_1389 (
   .O(gates[857]),
   .I0(gatesReg[1253]),
   .I1(gatesReg[928]),
   .I2(gatesReg[1265]),
   .I3(gatesReg[544]),
   .I4(gatesReg[623]),
   .I5(gatesReg[1512])
);
LUT6 #(
   .INIT(64'b0111101110000001110010101010011110000011011010001110110001000111)  
) LUT6_1390 (
   .O(gates[106]),
   .I0(gatesReg[1526]),
   .I1(gatesReg[1196]),
   .I2(gatesReg[1114]),
   .I3(gatesReg[217]),
   .I4(gatesReg[328]),
   .I5(gatesReg[239])
);
LUT6 #(
   .INIT(64'b1111100110010000010000001000101010110101010010010011001010010101)  
) LUT6_1391 (
   .O(gates[1010]),
   .I0(gatesReg[122]),
   .I1(gatesReg[1223]),
   .I2(gatesReg[878]),
   .I3(gatesReg[281]),
   .I4(gatesReg[269]),
   .I5(gatesReg[628])
);
LUT6 #(
   .INIT(64'b0001010011001011100111011001001110011010001001010011011100010011)  
) LUT6_1392 (
   .O(gates[707]),
   .I0(gatesReg[158]),
   .I1(gatesReg[363]),
   .I2(gatesReg[46]),
   .I3(gatesReg[1316]),
   .I4(gatesReg[733]),
   .I5(gatesReg[36])
);
LUT6 #(
   .INIT(64'b1110010001001000111001111111111111011011010110111011111111101001)  
) LUT6_1393 (
   .O(gates[964]),
   .I0(gatesReg[1418]),
   .I1(gatesReg[997]),
   .I2(gatesReg[630]),
   .I3(gatesReg[1368]),
   .I4(gatesReg[472]),
   .I5(gatesReg[748])
);
LUT6 #(
   .INIT(64'b0000110110100011111101010110110011101100000000111000011000011100)  
) LUT6_1394 (
   .O(gates[157]),
   .I0(gatesReg[1449]),
   .I1(gatesReg[317]),
   .I2(gatesReg[608]),
   .I3(gatesReg[711]),
   .I4(gatesReg[132]),
   .I5(gatesReg[1254])
);
LUT6 #(
   .INIT(64'b1110001010010110111011101000101011000101000001010001001010100110)  
) LUT6_1395 (
   .O(gates[65]),
   .I0(gatesReg[1234]),
   .I1(gatesReg[892]),
   .I2(gatesReg[1314]),
   .I3(gatesReg[546]),
   .I4(gatesReg[1428]),
   .I5(gatesReg[537])
);
LUT6 #(
   .INIT(64'b0101111101110110000110100001000011010101110011111101101111001100)  
) LUT6_1396 (
   .O(gates[935]),
   .I0(gatesReg[1474]),
   .I1(gatesReg[125]),
   .I2(gatesReg[522]),
   .I3(gatesReg[1423]),
   .I4(gatesReg[44]),
   .I5(gatesReg[1018])
);
LUT6 #(
   .INIT(64'b0011101000010011100011110111101001011110010110011001001110000110)  
) LUT6_1397 (
   .O(gates[203]),
   .I0(gatesReg[1125]),
   .I1(gatesReg[667]),
   .I2(gatesReg[1007]),
   .I3(gatesReg[1443]),
   .I4(gatesReg[741]),
   .I5(gatesReg[1188])
);
LUT6 #(
   .INIT(64'b1000100001000011000010110100111111100110101001010110000110010100)  
) LUT6_1398 (
   .O(gates[261]),
   .I0(gatesReg[1186]),
   .I1(gatesReg[998]),
   .I2(gatesReg[714]),
   .I3(gatesReg[1280]),
   .I4(gatesReg[313]),
   .I5(gatesReg[529])
);
LUT6 #(
   .INIT(64'b1010001100100000111111101010101111100010101111011100101100010001)  
) LUT6_1399 (
   .O(gates[1213]),
   .I0(gatesReg[1545]),
   .I1(gatesReg[1058]),
   .I2(gatesReg[987]),
   .I3(gatesReg[1324]),
   .I4(gatesReg[397]),
   .I5(gatesReg[1150])
);
LUT6 #(
   .INIT(64'b0010110001011110011111010000011101001001011010000101110011010111)  
) LUT6_1400 (
   .O(gates[1093]),
   .I0(gatesReg[1096]),
   .I1(gatesReg[1535]),
   .I2(gatesReg[1335]),
   .I3(gatesReg[908]),
   .I4(gatesReg[1191]),
   .I5(gatesReg[459])
);
LUT6 #(
   .INIT(64'b1001000100101110101001000101110000010101100011111110110001110011)  
) LUT6_1401 (
   .O(gates[1023]),
   .I0(gatesReg[284]),
   .I1(gatesReg[823]),
   .I2(gatesReg[903]),
   .I3(gatesReg[247]),
   .I4(gatesReg[1340]),
   .I5(gatesReg[165])
);
LUT6 #(
   .INIT(64'b0001011000111110000001111110010110111010001000110110011101110000)  
) LUT6_1402 (
   .O(gates[81]),
   .I0(gatesReg[289]),
   .I1(gatesReg[1495]),
   .I2(gatesReg[729]),
   .I3(gatesReg[2]),
   .I4(gatesReg[771]),
   .I5(gatesReg[808])
);
LUT6 #(
   .INIT(64'b1011101000010010000100011010111000011011011011110101110100111101)  
) LUT6_1403 (
   .O(gates[321]),
   .I0(gatesReg[401]),
   .I1(gatesReg[845]),
   .I2(gatesReg[186]),
   .I3(gatesReg[1231]),
   .I4(gatesReg[1119]),
   .I5(gatesReg[147])
);
LUT6 #(
   .INIT(64'b1101001110001000000011011000110100001011101001101101010101101000)  
) LUT6_1404 (
   .O(gates[1199]),
   .I0(gatesReg[1249]),
   .I1(gatesReg[973]),
   .I2(gatesReg[1046]),
   .I3(gatesReg[1142]),
   .I4(gatesReg[1291]),
   .I5(gatesReg[319])
);
LUT6 #(
   .INIT(64'b1110010010011011111010000100101101101001000000000000001100001101)  
) LUT6_1405 (
   .O(gates[624]),
   .I0(gatesReg[915]),
   .I1(gatesReg[1179]),
   .I2(gatesReg[1456]),
   .I3(gatesReg[1052]),
   .I4(gatesReg[404]),
   .I5(gatesReg[735])
);
LUT6 #(
   .INIT(64'b0011000001100001001011111100100011110000111100110011110010001111)  
) LUT6_1406 (
   .O(gates[1300]),
   .I0(gatesReg[516]),
   .I1(gatesReg[1493]),
   .I2(gatesReg[974]),
   .I3(gatesReg[1551]),
   .I4(gatesReg[702]),
   .I5(gatesReg[1271])
);
LUT6 #(
   .INIT(64'b0100011101110110011011111000100011001011110101011011001000000101)  
) LUT6_1407 (
   .O(gates[792]),
   .I0(gatesReg[344]),
   .I1(gatesReg[636]),
   .I2(gatesReg[1104]),
   .I3(gatesReg[1406]),
   .I4(gatesReg[561]),
   .I5(gatesReg[1133])
);
LUT6 #(
   .INIT(64'b0011000111000000101101000001011000010110101100101011010010111110)  
) LUT6_1408 (
   .O(gates[86]),
   .I0(gatesReg[209]),
   .I1(gatesReg[1118]),
   .I2(gatesReg[357]),
   .I3(gatesReg[117]),
   .I4(gatesReg[1307]),
   .I5(gatesReg[455])
);
LUT6 #(
   .INIT(64'b0000110100001010001110000011011101000001101110000011100001111100)  
) LUT6_1409 (
   .O(gates[1158]),
   .I0(gatesReg[80]),
   .I1(gatesReg[600]),
   .I2(gatesReg[336]),
   .I3(gatesReg[457]),
   .I4(gatesReg[1301]),
   .I5(gatesReg[821])
);
LUT6 #(
   .INIT(64'b0010111001000100101100001110001001010110010110010111011100011110)  
) LUT6_1410 (
   .O(gates[371]),
   .I0(gatesReg[383]),
   .I1(gatesReg[696]),
   .I2(gatesReg[297]),
   .I3(gatesReg[963]),
   .I4(gatesReg[1431]),
   .I5(gatesReg[92])
);
LUT6 #(
   .INIT(64'b0110101010000111110110101001000110010010100100110111000101000111)  
) LUT6_1411 (
   .O(gates[656]),
   .I0(gatesReg[1489]),
   .I1(gatesReg[1212]),
   .I2(gatesReg[10]),
   .I3(gatesReg[980]),
   .I4(gatesReg[550]),
   .I5(gatesReg[1477])
);
LUT6 #(
   .INIT(64'b1000110010111010000000100111110011111010101000101111111010010001)  
) LUT6_1412 (
   .O(gates[1079]),
   .I0(gatesReg[1164]),
   .I1(gatesReg[1081]),
   .I2(gatesReg[505]),
   .I3(gatesReg[670]),
   .I4(gatesReg[1094]),
   .I5(gatesReg[958])
);
LUT6 #(
   .INIT(64'b0110111100100011011101101100100011010001100001011111001000110100)  
) LUT6_1413 (
   .O(gates[204]),
   .I0(gatesReg[419]),
   .I1(gatesReg[995]),
   .I2(gatesReg[1225]),
   .I3(gatesReg[837]),
   .I4(gatesReg[290]),
   .I5(gatesReg[592])
);
LUT6 #(
   .INIT(64'b0100001100110100001110011111011010010000100110011001101100010100)  
) LUT6_1414 (
   .O(gates[1248]),
   .I0(gatesReg[149]),
   .I1(gatesReg[625]),
   .I2(gatesReg[712]),
   .I3(gatesReg[210]),
   .I4(gatesReg[406]),
   .I5(gatesReg[173])
);
LUT6 #(
   .INIT(64'b0010001110101100000101011110101010111001111110001110110001001110)  
) LUT6_1415 (
   .O(gates[1041]),
   .I0(gatesReg[530]),
   .I1(gatesReg[66]),
   .I2(gatesReg[19]),
   .I3(gatesReg[1030]),
   .I4(gatesReg[365]),
   .I5(gatesReg[763])
);
LUT6 #(
   .INIT(64'b0101101000011000110011111101111010110011100001111010011011111100)  
) LUT6_1416 (
   .O(gates[435]),
   .I0(gatesReg[470]),
   .I1(gatesReg[1524]),
   .I2(gatesReg[793]),
   .I3(gatesReg[1205]),
   .I4(gatesReg[1287]),
   .I5(gatesReg[654])
);
LUT6 #(
   .INIT(64'b0110111011111011110001101000000001000011001001010001000101001010)  
) LUT6_1417 (
   .O(gates[814]),
   .I0(gatesReg[570]),
   .I1(gatesReg[252]),
   .I2(gatesReg[1159]),
   .I3(gatesReg[883]),
   .I4(gatesReg[283]),
   .I5(gatesReg[156])
);
LUT6 #(
   .INIT(64'b1001111011101101000000000001001001010101000000101000001111111100)  
) LUT6_1418 (
   .O(gates[1516]),
   .I0(gatesReg[655]),
   .I1(gatesReg[421]),
   .I2(gatesReg[59]),
   .I3(gatesReg[1367]),
   .I4(gatesReg[271]),
   .I5(gatesReg[1226])
);
LUT6 #(
   .INIT(64'b0111001101101010110010110110111000011100101001101000011100101111)  
) LUT6_1419 (
   .O(gates[1482]),
   .I0(gatesReg[1256]),
   .I1(gatesReg[1070]),
   .I2(gatesReg[1024]),
   .I3(gatesReg[491]),
   .I4(gatesReg[864]),
   .I5(gatesReg[219])
);
LUT6 #(
   .INIT(64'b1010111110001101110111001111010110011100100111111001110101000111)  
) LUT6_1420 (
   .O(gates[924]),
   .I0(gatesReg[1016]),
   .I1(gatesReg[13]),
   .I2(gatesReg[799]),
   .I3(gatesReg[1170]),
   .I4(gatesReg[105]),
   .I5(gatesReg[1514])
);
LUT6 #(
   .INIT(64'b0101010110111011100101001100011101001100111111000110100010010101)  
) LUT6_1421 (
   .O(gates[885]),
   .I0(gatesReg[925]),
   .I1(gatesReg[840]),
   .I2(gatesReg[597]),
   .I3(gatesReg[390]),
   .I4(gatesReg[111]),
   .I5(gatesReg[1042])
);
LUT6 #(
   .INIT(64'b0110000000011010101100010101000011101011001100100111011000100011)  
) LUT6_1422 (
   .O(gates[884]),
   .I0(gatesReg[1515]),
   .I1(gatesReg[38]),
   .I2(gatesReg[408]),
   .I3(gatesReg[1411]),
   .I4(gatesReg[1480]),
   .I5(gatesReg[196])
);
LUT6 #(
   .INIT(64'b1011011100110000111100111011101110011010001011011111010110000011)  
) LUT6_1423 (
   .O(gates[1412]),
   .I0(gatesReg[945]),
   .I1(gatesReg[242]),
   .I2(gatesReg[1169]),
   .I3(gatesReg[559]),
   .I4(gatesReg[32]),
   .I5(gatesReg[118])
);
LUT6 #(
   .INIT(64'b0101100110011100001001100000100010011110000010101010001110111111)  
) LUT6_1424 (
   .O(gates[339]),
   .I0(gatesReg[443]),
   .I1(gatesReg[206]),
   .I2(gatesReg[959]),
   .I3(gatesReg[358]),
   .I4(gatesReg[331]),
   .I5(gatesReg[1065])
);
LUT6 #(
   .INIT(64'b0000000101101011010110111001111000001111100100100000001110111001)  
) LUT6_1425 (
   .O(gates[760]),
   .I0(gatesReg[737]),
   .I1(gatesReg[580]),
   .I2(gatesReg[767]),
   .I3(gatesReg[84]),
   .I4(gatesReg[805]),
   .I5(gatesReg[1020])
);
LUT6 #(
   .INIT(64'b0011101000000100010100101011100000110110000010110110000100110100)  
) LUT6_1426 (
   .O(gates[228]),
   .I0(gatesReg[437]),
   .I1(gatesReg[194]),
   .I2(gatesReg[220]),
   .I3(gatesReg[1312]),
   .I4(gatesReg[1257]),
   .I5(gatesReg[846])
);
LUT6 #(
   .INIT(64'b1100110101000111001010101100011101011110010001111001000011000011)  
) LUT6_1427 (
   .O(gates[863]),
   .I0(gatesReg[1021]),
   .I1(gatesReg[31]),
   .I2(gatesReg[1263]),
   .I3(gatesReg[934]),
   .I4(gatesReg[1296]),
   .I5(gatesReg[1553])
);
LUT6 #(
   .INIT(64'b1001001011110000011010111110111100011101100101010110101011010111)  
) LUT6_1428 (
   .O(gates[749]),
   .I0(gatesReg[948]),
   .I1(gatesReg[1303]),
   .I2(gatesReg[572]),
   .I3(gatesReg[968]),
   .I4(gatesReg[675]),
   .I5(gatesReg[1398])
);
LUT6 #(
   .INIT(64'b0111011010100100000000001100100110100100001111011010111100000100)  
) LUT6_1429 (
   .O(gates[531]),
   .I0(gatesReg[226]),
   .I1(gatesReg[15]),
   .I2(gatesReg[527]),
   .I3(gatesReg[431]),
   .I4(gatesReg[1430]),
   .I5(gatesReg[1145])
);
LUT6 #(
   .INIT(64'b1010101110101110011101000000111100111101001010011110100000011101)  
) LUT6_1430 (
   .O(gates[268]),
   .I0(gatesReg[382]),
   .I1(gatesReg[1448]),
   .I2(gatesReg[1506]),
   .I3(gatesReg[62]),
   .I4(gatesReg[833]),
   .I5(gatesReg[139])
);
LUT6 #(
   .INIT(64'b0101110100101000100101110100101100010000000110100110100001011001)  
) LUT6_1431 (
   .O(gates[829]),
   .I0(gatesReg[129]),
   .I1(gatesReg[1472]),
   .I2(gatesReg[548]),
   .I3(gatesReg[926]),
   .I4(gatesReg[859]),
   .I5(gatesReg[1246])
);
LUT6 #(
   .INIT(64'b0011110101101110110000000100011101001110001111011101101010000101)  
) LUT6_1432 (
   .O(gates[345]),
   .I0(gatesReg[1083]),
   .I1(gatesReg[739]),
   .I2(gatesReg[1110]),
   .I3(gatesReg[1293]),
   .I4(gatesReg[876]),
   .I5(gatesReg[662])
);
LUT6 #(
   .INIT(64'b0100111101111111001010110100101001111010111011010010101111100011)  
) LUT6_1433 (
   .O(gates[172]),
   .I0(gatesReg[418]),
   .I1(gatesReg[783]),
   .I2(gatesReg[933]),
   .I3(gatesReg[168]),
   .I4(gatesReg[1357]),
   .I5(gatesReg[135])
);
LUT6 #(
   .INIT(64'b1000000101010100101011110111101100010100111101011001001110100010)  
) LUT6_1434 (
   .O(gates[596]),
   .I0(gatesReg[348]),
   .I1(gatesReg[1518]),
   .I2(gatesReg[1152]),
   .I3(gatesReg[145]),
   .I4(gatesReg[789]),
   .I5(gatesReg[49])
);
LUT6 #(
   .INIT(64'b1110011111001001011001011100111001011111001111100011011111111001)  
) LUT6_1435 (
   .O(gates[1297]),
   .I0(gatesReg[178]),
   .I1(gatesReg[1131]),
   .I2(gatesReg[124]),
   .I3(gatesReg[772]),
   .I4(gatesReg[993]),
   .I5(gatesReg[1090])
);
LUT6 #(
   .INIT(64'b1100011000010101101110110011000010011011010000100110000111010100)  
) LUT6_1436 (
   .O(gates[1521]),
   .I0(gatesReg[627]),
   .I1(gatesReg[1308]),
   .I2(gatesReg[1429]),
   .I3(gatesReg[715]),
   .I4(gatesReg[1374]),
   .I5(gatesReg[23])
);
LUT6 #(
   .INIT(64'b0000010100100101001001111000101101101001101011001010000111010011)  
) LUT6_1437 (
   .O(gates[1366]),
   .I0(gatesReg[388]),
   .I1(gatesReg[364]),
   .I2(gatesReg[1528]),
   .I3(gatesReg[653]),
   .I4(gatesReg[1425]),
   .I5(gatesReg[950])
);
LUT6 #(
   .INIT(64'b1000000011010001101111010001001001001010001000100000011110101110)  
) LUT6_1438 (
   .O(gates[223]),
   .I0(gatesReg[1445]),
   .I1(gatesReg[1025]),
   .I2(gatesReg[509]),
   .I3(gatesReg[1015]),
   .I4(gatesReg[976]),
   .I5(gatesReg[367])
);
LUT6 #(
   .INIT(64'b0100101100011001101101010001001110010101010100000000000100111010)  
) LUT6_1439 (
   .O(gates[613]),
   .I0(gatesReg[716]),
   .I1(gatesReg[940]),
   .I2(gatesReg[1466]),
   .I3(gatesReg[485]),
   .I4(gatesReg[743]),
   .I5(gatesReg[778])
);
LUT6 #(
   .INIT(64'b1110000101111101100000011111101101001011111110000000001001100110)  
) LUT6_1440 (
   .O(gates[721]),
   .I0(gatesReg[685]),
   .I1(gatesReg[21]),
   .I2(gatesReg[523]),
   .I3(gatesReg[720]),
   .I4(gatesReg[1270]),
   .I5(gatesReg[460])
);
LUT6 #(
   .INIT(64'b0001000111110101000011110101000010110010100000100111001101111001)  
) LUT6_1441 (
   .O(gates[1043]),
   .I0(gatesReg[723]),
   .I1(gatesReg[324]),
   .I2(gatesReg[453]),
   .I3(gatesReg[1389]),
   .I4(gatesReg[1460]),
   .I5(gatesReg[244])
);
LUT6 #(
   .INIT(64'b1110101000101111101111001001111110100111100011001110000101010111)  
) LUT6_1442 (
   .O(gates[1255]),
   .I0(gatesReg[1202]),
   .I1(gatesReg[637]),
   .I2(gatesReg[351]),
   .I3(gatesReg[1040]),
   .I4(gatesReg[595]),
   .I5(gatesReg[1138])
);
LUT6 #(
   .INIT(64'b1100011110101101110100010000011111011011111101011001111001000111)  
) LUT6_1443 (
   .O(gates[669]),
   .I0(gatesReg[488]),
   .I1(gatesReg[752]),
   .I2(gatesReg[1012]),
   .I3(gatesReg[1232]),
   .I4(gatesReg[1498]),
   .I5(gatesReg[835])
);
LUT6 #(
   .INIT(64'b0010100001100000101001101001100001101010000100010101101011001111)  
) LUT6_1444 (
   .O(gates[282]),
   .I0(gatesReg[1267]),
   .I1(gatesReg[379]),
   .I2(gatesReg[1032]),
   .I3(gatesReg[1386]),
   .I4(gatesReg[113]),
   .I5(gatesReg[1536])
);
LUT6 #(
   .INIT(64'b1010100000100110101000001111000111101001000000001111101111000010)  
) LUT6_1445 (
   .O(gates[1082]),
   .I0(gatesReg[901]),
   .I1(gatesReg[1035]),
   .I2(gatesReg[152]),
   .I3(gatesReg[342]),
   .I4(gatesReg[452]),
   .I5(gatesReg[862])
);
LUT6 #(
   .INIT(64'b1110001001101001111001010000010101011101001101111010001111111100)  
) LUT6_1446 (
   .O(gates[420]),
   .I0(gatesReg[1419]),
   .I1(gatesReg[579]),
   .I2(gatesReg[295]),
   .I3(gatesReg[341]),
   .I4(gatesReg[1056]),
   .I5(gatesReg[535])
);
LUT6 #(
   .INIT(64'b1001000101111001101001110001010000010000010110001111111100110011)  
) LUT6_1447 (
   .O(gates[121]),
   .I0(gatesReg[77]),
   .I1(gatesReg[683]),
   .I2(gatesReg[541]),
   .I3(gatesReg[1215]),
   .I4(gatesReg[64]),
   .I5(gatesReg[1473])
);
LUT6 #(
   .INIT(64'b0111111110101101100101101011001110001011100101000001101000001100)  
) LUT6_1448 (
   .O(gates[1066]),
   .I0(gatesReg[765]),
   .I1(gatesReg[881]),
   .I2(gatesReg[312]),
   .I3(gatesReg[897]),
   .I4(gatesReg[45]),
   .I5(gatesReg[405])
);
LUT6 #(
   .INIT(64'b1011100101111100010011101010110011110101101111111111011010110010)  
) LUT6_1449 (
   .O(gates[952]),
   .I0(gatesReg[507]),
   .I1(gatesReg[237]),
   .I2(gatesReg[1002]),
   .I3(gatesReg[1173]),
   .I4(gatesReg[370]),
   .I5(gatesReg[309])
);
LUT6 #(
   .INIT(64'b1101000010011101111001001111000110101110110000100010001001001001)  
) LUT6_1450 (
   .O(gates[639]),
   .I0(gatesReg[567]),
   .I1(gatesReg[416]),
   .I2(gatesReg[380]),
   .I3(gatesReg[100]),
   .I4(gatesReg[914]),
   .I5(gatesReg[300])
);
LUT6 #(
   .INIT(64'b1011100011111011111010001000110110111101101100100001000011111111)  
) LUT6_1451 (
   .O(gates[989]),
   .I0(gatesReg[1279]),
   .I1(gatesReg[965]),
   .I2(gatesReg[1258]),
   .I3(gatesReg[1439]),
   .I4(gatesReg[824]),
   .I5(gatesReg[286])
);
LUT6 #(
   .INIT(64'b0001101010001010110011101100101111011000110110110000010100000110)  
) LUT6_1452 (
   .O(gates[494]),
   .I0(gatesReg[1395]),
   .I1(gatesReg[120]),
   .I2(gatesReg[1075]),
   .I3(gatesReg[800]),
   .I4(gatesReg[1148]),
   .I5(gatesReg[392])
);
LUT6 #(
   .INIT(64'b1111011111100101010011101101101111111011110000011011110010111100)  
) LUT6_1453 (
   .O(gates[1505]),
   .I0(gatesReg[254]),
   .I1(gatesReg[1321]),
   .I2(gatesReg[1365]),
   .I3(gatesReg[1407]),
   .I4(gatesReg[496]),
   .I5(gatesReg[605])
);
LUT6 #(
   .INIT(64'b0111111110110100011010010111010011010100000000010001100100101100)  
) LUT6_1454 (
   .O(gates[487]),
   .I0(gatesReg[607]),
   .I1(gatesReg[813]),
   .I2(gatesReg[42]),
   .I3(gatesReg[759]),
   .I4(gatesReg[644]),
   .I5(gatesReg[851])
);
LUT6 #(
   .INIT(64'b1000100010000011111110110011010011111000100011010111001111000011)  
) LUT6_1455 (
   .O(gates[1071]),
   .I0(gatesReg[399]),
   .I1(gatesReg[1228]),
   .I2(gatesReg[235]),
   .I3(gatesReg[1073]),
   .I4(gatesReg[694]),
   .I5(gatesReg[436])
);
LUT6 #(
   .INIT(64'b1010101000000110001011101110001000010110011100110010100111110000)  
) LUT6_1456 (
   .O(gates[1348]),
   .I0(gatesReg[1342]),
   .I1(gatesReg[94]),
   .I2(gatesReg[213]),
   .I3(gatesReg[816]),
   .I4(gatesReg[1103]),
   .I5(gatesReg[1450])
);
LUT6 #(
   .INIT(64'b1111001111001011111000101100001010110010001010100001100010000101)  
) LUT6_1457 (
   .O(gates[238]),
   .I0(gatesReg[568]),
   .I1(gatesReg[296]),
   .I2(gatesReg[265]),
   .I3(gatesReg[1062]),
   .I4(gatesReg[1129]),
   .I5(gatesReg[791])
);
LUT6 #(
   .INIT(64'b1101000001100110011100010001010110111010001011000100011111001000)  
) LUT6_1458 (
   .O(gates[873]),
   .I0(gatesReg[171]),
   .I1(gatesReg[1143]),
   .I2(gatesReg[1355]),
   .I3(gatesReg[386]),
   .I4(gatesReg[916]),
   .I5(gatesReg[1457])
);
LUT6 #(
   .INIT(64'b0101111010101001100010101100011100000010001010101010101100100101)  
) LUT6_1459 (
   .O(gates[577]),
   .I0(gatesReg[445]),
   .I1(gatesReg[200]),
   .I2(gatesReg[1339]),
   .I3(gatesReg[1261]),
   .I4(gatesReg[1352]),
   .I5(gatesReg[329])
);
LUT6 #(
   .INIT(64'b1000100001101111101101010111000100101001010101111111100001001100)  
) LUT6_1460 (
   .O(gates[1137]),
   .I0(gatesReg[525]),
   .I1(gatesReg[27]),
   .I2(gatesReg[787]),
   .I3(gatesReg[161]),
   .I4(gatesReg[582]),
   .I5(gatesReg[109])
);
LUT6 #(
   .INIT(64'b0111101111101111001101111001001010001010111011011001011011011001)  
) LUT6_1461 (
   .O(gates[253]),
   .I0(gatesReg[1310]),
   .I1(gatesReg[557]),
   .I2(gatesReg[718]),
   .I3(gatesReg[1507]),
   .I4(gatesReg[1239]),
   .I5(gatesReg[441])
);
LUT6 #(
   .INIT(64'b0001100000010101011100011010000010101110110001010011111011011100)  
) LUT6_1462 (
   .O(gates[448]),
   .I0(gatesReg[868]),
   .I1(gatesReg[672]),
   .I2(gatesReg[769]),
   .I3(gatesReg[1140]),
   .I4(gatesReg[1181]),
   .I5(gatesReg[275])
);
LUT6 #(
   .INIT(64'b0100110000101111001011101011101101011000100111100001001001001010)  
) LUT6_1463 (
   .O(gates[1227]),
   .I0(gatesReg[983]),
   .I1(gatesReg[803]),
   .I2(gatesReg[197]),
   .I3(gatesReg[853]),
   .I4(gatesReg[751]),
   .I5(gatesReg[60])
);
LUT6 #(
   .INIT(64'b0001101001000100000010011010111010110110100111110110001100000100)  
) LUT6_1464 (
   .O(gates[1417]),
   .I0(gatesReg[1500]),
   .I1(gatesReg[1245]),
   .I2(gatesReg[1400]),
   .I3(gatesReg[691]),
   .I4(gatesReg[1067]),
   .I5(gatesReg[1388])
);
LUT6 #(
   .INIT(64'b1011111111000011010010101110001011111001001101111111110101101000)  
) LUT6_1465 (
   .O(gates[216]),
   .I0(gatesReg[346]),
   .I1(gatesReg[911]),
   .I2(gatesReg[1295]),
   .I3(gatesReg[427]),
   .I4(gatesReg[1111]),
   .I5(gatesReg[677])
);
LUT6 #(
   .INIT(64'b0101011111110000010111000001001000100110000111011000001101010111)  
) LUT6_1466 (
   .O(gates[852]),
   .I0(gatesReg[907]),
   .I1(gatesReg[82]),
   .I2(gatesReg[650]),
   .I3(gatesReg[1154]),
   .I4(gatesReg[590]),
   .I5(gatesReg[1210])
);
LUT6 #(
   .INIT(64'b0011110111010011111100101010101111101110011110100000000011000110)  
) LUT6_1467 (
   .O(gates[643]),
   .I0(gatesReg[895]),
   .I1(gatesReg[69]),
   .I2(gatesReg[1157]),
   .I3(gatesReg[664]),
   .I4(gatesReg[1470]),
   .I5(gatesReg[224])
);
LUT6 #(
   .INIT(64'b0101110110101101001101101010100010101010000001111010101001111100)  
) LUT6_1468 (
   .O(gates[63]),
   .I0(gatesReg[617]),
   .I1(gatesReg[79]),
   .I2(gatesReg[1420]),
   .I3(gatesReg[352]),
   .I4(gatesReg[1006]),
   .I5(gatesReg[126])
);
LUT6 #(
   .INIT(64'b0010111101110001001100101011000010001010010110001100010000101011)  
) LUT6_1469 (
   .O(gates[1120]),
   .I0(gatesReg[251]),
   .I1(gatesReg[1034]),
   .I2(gatesReg[426]),
   .I3(gatesReg[369]),
   .I4(gatesReg[996]),
   .I5(gatesReg[1533])
);
LUT6 #(
   .INIT(64'b1001101110110001111110101100010101101110011110101111011010100110)  
) LUT6_1470 (
   .O(gates[179]),
   .I0(gatesReg[1548]),
   .I1(gatesReg[1435]),
   .I2(gatesReg[651]),
   .I3(gatesReg[279]),
   .I4(gatesReg[176]),
   .I5(gatesReg[956])
);
LUT6 #(
   .INIT(64'b1001010010100100111101010001101010110110110101000011101111101100)  
) LUT6_1471 (
   .O(gates[1532]),
   .I0(gatesReg[498]),
   .I1(gatesReg[483]),
   .I2(gatesReg[629]),
   .I3(gatesReg[947]),
   .I4(gatesReg[256]),
   .I5(gatesReg[372])
);
LUT6 #(
   .INIT(64'b1011001001010000000000011011100111100111001101001111110110100000)  
) LUT6_1472 (
   .O(gates[1475]),
   .I0(gatesReg[1487]),
   .I1(gatesReg[1540]),
   .I2(gatesReg[920]),
   .I3(gatesReg[1330]),
   .I4(gatesReg[1284]),
   .I5(gatesReg[428])
);
LUT6 #(
   .INIT(64'b0010000111101011010111111001111010011110011000000100110111000010)  
) LUT6_1473 (
   .O(gates[1105]),
   .I0(gatesReg[887]),
   .I1(gatesReg[99]),
   .I2(gatesReg[1160]),
   .I3(gatesReg[72]),
   .I4(gatesReg[869]),
   .I5(gatesReg[500])
);
LUT6 #(
   .INIT(64'b1000010011110101010001000110111011111011110010111111111001111100)  
) LUT6_1474 (
   .O(gates[1187]),
   .I0(gatesReg[1496]),
   .I1(gatesReg[1221]),
   .I2(gatesReg[1200]),
   .I3(gatesReg[790]),
   .I4(gatesReg[533]),
   .I5(gatesReg[918])
);
LUT6 #(
   .INIT(64'b0000111110001101110110000110101110010000111111101001010010001100)  
) LUT6_1475 (
   .O(gates[713]),
   .I0(gatesReg[1413]),
   .I1(gatesReg[1122]),
   .I2(gatesReg[1275]),
   .I3(gatesReg[1108]),
   .I4(gatesReg[1053]),
   .I5(gatesReg[414])
);
LUT6 #(
   .INIT(64'b0111101001100001111101011001111000101101111110111001010000111100)  
) LUT6_1476 (
   .O(gates[676]),
   .I0(gatesReg[462]),
   .I1(gatesReg[1014]),
   .I2(gatesReg[843]),
   .I3(gatesReg[1491]),
   .I4(gatesReg[1362]),
   .I5(gatesReg[1209])
);
LUT6 #(
   .INIT(64'b1001011100111010110001001111110110101101111101000111101011010111)  
) LUT6_1477 (
   .O(gates[1334]),
   .I0(gatesReg[632]),
   .I1(gatesReg[263]),
   .I2(gatesReg[1371]),
   .I3(gatesReg[991]),
   .I4(gatesReg[394]),
   .I5(gatesReg[514])
);
LUT6 #(
   .INIT(64'b0111001001111000001000110111110110111010101110110100000110000011)  
) LUT6_1478 (
   .O(gates[1251]),
   .I0(gatesReg[610]),
   .I1(gatesReg[725]),
   .I2(gatesReg[931]),
   .I3(gatesReg[513]),
   .I4(gatesReg[615]),
   .I5(gatesReg[50])
);
LUT6 #(
   .INIT(64'b1000001001100000010111001110001100001011111111000110000110010001)  
) LUT6_1479 (
   .O(gates[277]),
   .I0(gatesReg[476]),
   .I1(gatesReg[1198]),
   .I2(gatesReg[1519]),
   .I3(gatesReg[1409]),
   .I4(gatesReg[797]),
   .I5(gatesReg[1077])
);
LUT6 #(
   .INIT(64'b1111011100110011100101011100101110110111000100111101111111101001)  
) LUT6_1480 (
   .O(gates[1192]),
   .I0(gatesReg[1136]),
   .I1(gatesReg[1175]),
   .I2(gatesReg[293]),
   .I3(gatesReg[1272]),
   .I4(gatesReg[1299]),
   .I5(gatesReg[1236])
);
LUT6 #(
   .INIT(64'b0100101011011010011101001000100100010010010110100101011010001101)  
) LUT6_1481 (
   .O(gates[879]),
   .I0(gatesReg[967]),
   .I1(gatesReg[322]),
   .I2(gatesReg[645]),
   .I3(gatesReg[1326]),
   .I4(gatesReg[469]),
   .I5(gatesReg[635])
);
LUT6 #(
   .INIT(64'b0011011011000011110110100001101010101001011111110010111011100101)  
) LUT6_1482 (
   .O(gates[938]),
   .I0(gatesReg[575]),
   .I1(gatesReg[1088]),
   .I2(gatesReg[1382]),
   .I3(gatesReg[1176]),
   .I4(gatesReg[1452]),
   .I5(gatesReg[1039])
);
LUT6 #(
   .INIT(64'b1111010011111110001001000010011011110111101100100001011001101000)  
) LUT6_1483 (
   .O(gates[1095]),
   .I0(gatesReg[979]),
   .I1(gatesReg[709]),
   .I2(gatesReg[1005]),
   .I3(gatesReg[28]),
   .I4(gatesReg[40]),
   .I5(gatesReg[310])
);
LUT6 #(
   .INIT(64'b0101001110101011110000000100100010001100111111001111100001101101)  
) LUT6_1484 (
   .O(gates[1183]),
   .I0(gatesReg[192]),
   .I1(gatesReg[589]),
   .I2(gatesReg[1337]),
   .I3(gatesReg[699]),
   .I4(gatesReg[215]),
   .I5(gatesReg[687])
);
LUT6 #(
   .INIT(64'b0111010010100111100101010000001111010001000001011001010100001000)  
) LUT6_1485 (
   .O(gates[1262]),
   .I0(gatesReg[1115]),
   .I1(gatesReg[960]),
   .I2(gatesReg[818]),
   .I3(gatesReg[150]),
   .I4(gatesReg[1038]),
   .I5(gatesReg[245])
);
LUT6 #(
   .INIT(64'b0111100011101001111010001000001111100011100100001100000011010101)  
) LUT6_1486 (
   .O(gates[1444]),
   .I0(gatesReg[543]),
   .I1(gatesReg[267]),
   .I2(gatesReg[826]),
   .I3(gatesReg[354]),
   .I4(gatesReg[1437]),
   .I5(gatesReg[1344])
);
LUT6 #(
   .INIT(64'b1111110110000011101100001011001011001111110000010000000010110110)  
) LUT6_1487 (
   .O(gates[1290]),
   .I0(gatesReg[1064]),
   .I1(gatesReg[757]),
   .I2(gatesReg[332]),
   .I3(gatesReg[9]),
   .I4(gatesReg[1099]),
   .I5(gatesReg[1217])
);
LUT6 #(
   .INIT(64'b0011100111100101001011010001101111001111101111101110111011011110)  
) LUT6_1488 (
   .O(gates[1527]),
   .I0(gatesReg[745]),
   .I1(gatesReg[34]),
   .I2(gatesReg[603]),
   .I3(gatesReg[90]),
   .I4(gatesReg[620]),
   .I5(gatesReg[565])
);
LUT6 #(
   .INIT(64'b1111100110010011011110110000010100101011111101010111001001011011)  
) LUT6_1489 (
   .O(gates[1132]),
   .I0(gatesReg[1410]),
   .I1(gatesReg[1346]),
   .I2(gatesReg[1434]),
   .I3(gatesReg[850]),
   .I4(gatesReg[1547]),
   .I5(gatesReg[891])
);
LUT6 #(
   .INIT(64'b0011101011010010110000110100001010110001011111100101100001011010)  
) LUT6_1490 (
   .O(gates[929]),
   .I0(gatesReg[1045]),
   .I1(gatesReg[937]),
   .I2(gatesReg[1004]),
   .I3(gatesReg[730]),
   .I4(gatesReg[16]),
   .I5(gatesReg[921])
);
LUT6 #(
   .INIT(64'b0010010101011110010111000110000111010101000011010111000110010111)  
) LUT6_1491 (
   .O(gates[133]),
   .I0(gatesReg[1360]),
   .I1(gatesReg[1013]),
   .I2(gatesReg[1069]),
   .I3(gatesReg[233]),
   .I4(gatesReg[1224]),
   .I5(gatesReg[1490])
);
LUT6 #(
   .INIT(64'b0101100101001000101001001111111000011101101011100010001011111100)  
) LUT6_1492 (
   .O(gates[123]),
   .I0(gatesReg[368]),
   .I1(gatesReg[316]),
   .I2(gatesReg[994]),
   .I3(gatesReg[611]),
   .I4(gatesReg[1370]),
   .I5(gatesReg[849])
);
LUT6 #(
   .INIT(64'b1110110001011000110010100010011101101000001000110011011111111000)  
) LUT6_1493 (
   .O(gates[304]),
   .I0(gatesReg[11]),
   .I1(gatesReg[492]),
   .I2(gatesReg[208]),
   .I3(gatesReg[842]),
   .I4(gatesReg[511]),
   .I5(gatesReg[1523])
);
LUT6 #(
   .INIT(64'b0010100110010001001110000111111101111101111010111110001011000100)  
) LUT6_1494 (
   .O(gates[547]),
   .I0(gatesReg[93]),
   .I1(gatesReg[899]),
   .I2(gatesReg[292]),
   .I3(gatesReg[291]),
   .I4(gatesReg[374]),
   .I5(gatesReg[114])
);
LUT6 #(
   .INIT(64'b0101001101000111000110101101100001010001011111000000100000010000)  
) LUT6_1495 (
   .O(gates[631]),
   .I0(gatesReg[199]),
   .I1(gatesReg[429]),
   .I2(gatesReg[1306]),
   .I3(gatesReg[1328]),
   .I4(gatesReg[1091]),
   .I5(gatesReg[73])
);
LUT6 #(
   .INIT(64'b0110001011001010010000111100011000110011110000010111101100010100)  
) LUT6_1496 (
   .O(gates[1538]),
   .I0(gatesReg[409]),
   .I1(gatesReg[67]),
   .I2(gatesReg[812]),
   .I3(gatesReg[241]),
   .I4(gatesReg[795]),
   .I5(gatesReg[489])
);
LUT6 #(
   .INIT(64'b1001001110111000000111111000010100000011110010110101101111111011)  
) LUT6_1497 (
   .O(gates[1544]),
   .I0(gatesReg[585]),
   .I1(gatesReg[794]),
   .I2(gatesReg[327]),
   .I3(gatesReg[1392]),
   .I4(gatesReg[1080]),
   .I5(gatesReg[944])
);
LUT6 #(
   .INIT(64'b0100100000101000101011011100100101010111111000011011101010000010)  
) LUT6_1498 (
   .O(gates[396]),
   .I0(gatesReg[1281]),
   .I1(gatesReg[1113]),
   .I2(gatesReg[732]),
   .I3(gatesReg[674]),
   .I4(gatesReg[1317]),
   .I5(gatesReg[280])
);
LUT6 #(
   .INIT(64'b0010001000011110110110111010101011110011010110110011100010100000)  
) LUT6_1499 (
   .O(gates[258]),
   .I0(gatesReg[957]),
   .I1(gatesReg[273]),
   .I2(gatesReg[471]),
   .I3(gatesReg[622]),
   .I4(gatesReg[1503]),
   .I5(gatesReg[970])
);
LUT6 #(
   .INIT(64'b0011010100010110101110011011001111101100111010010100001100100010)  
) LUT6_1500 (
   .O(gates[1422]),
   .I0(gatesReg[1509]),
   .I1(gatesReg[1416]),
   .I2(gatesReg[24]),
   .I3(gatesReg[104]),
   .I4(gatesReg[1325]),
   .I5(gatesReg[131])
);
LUT6 #(
   .INIT(64'b0001001010110001011000101110101010110011100110110100100111111110)  
) LUT6_1501 (
   .O(gates[482]),
   .I0(gatesReg[502]),
   .I1(gatesReg[314]),
   .I2(gatesReg[1286]),
   .I3(gatesReg[1237]),
   .I4(gatesReg[1513]),
   .I5(gatesReg[1502])
);
LUT6 #(
   .INIT(64'b1011001000110010111101001111110001101101100010010111100110000100)  
) LUT6_1502 (
   .O(gates[949]),
   .I0(gatesReg[1264]),
   .I1(gatesReg[355]),
   .I2(gatesReg[553]),
   .I3(gatesReg[159]),
   .I4(gatesReg[747]),
   .I5(gatesReg[1252])
);
LUT6 #(
   .INIT(64'b0011010001101100011000110101000010011010000111111011100001010111)  
) LUT6_1503 (
   .O(gates[499]),
   .I0(gatesReg[555]),
   .I1(gatesReg[47]),
   .I2(gatesReg[1037]),
   .I3(gatesReg[1427]),
   .I4(gatesReg[1484]),
   .I5(gatesReg[37])
);
LUT6 #(
   .INIT(64'b0100100101110111110010011111001011101010100011011000011000011010)  
) LUT6_1504 (
   .O(gates[56]),
   .I0(gatesReg[1017]),
   .I1(gatesReg[855]),
   .I2(gatesReg[270]),
   .I3(gatesReg[195]),
   .I4(gatesReg[1057]),
   .I5(gatesReg[538])
);
LUT6 #(
   .INIT(64'b0100000011101000101100010111010100001101100111000111001101001101)  
) LUT6_1505 (
   .O(gates[1369]),
   .I0(gatesReg[679]),
   .I1(gatesReg[680]),
   .I2(gatesReg[831]),
   .I3(gatesReg[521]),
   .I4(gatesReg[1147]),
   .I5(gatesReg[1332])
);
LUT6 #(
   .INIT(64'b0100011010101100011100111111100110100000011100001101110010000101)  
) LUT6_1506 (
   .O(gates[54]),
   .I0(gatesReg[162]),
   .I1(gatesReg[1241]),
   .I2(gatesReg[433]),
   .I3(gatesReg[880]),
   .I4(gatesReg[1441]),
   .I5(gatesReg[647])
);
LUT6 #(
   .INIT(64'b1101111011010100111100110101111100000010010110111010010010011100)  
) LUT6_1507 (
   .O(gates[1151]),
   .I0(gatesReg[1399]),
   .I1(gatesReg[1206]),
   .I2(gatesReg[334]),
   .I3(gatesReg[986]),
   .I4(gatesReg[786]),
   .I5(gatesReg[1117])
);
LUT6 #(
   .INIT(64'b0100000111111011001011010010101111110100111000100110110011101001)  
) LUT6_1508 (
   .O(gates[306]),
   .I0(gatesReg[740]),
   .I1(gatesReg[1008]),
   .I2(gatesReg[1027]),
   .I3(gatesReg[103]),
   .I4(gatesReg[201]),
   .I5(gatesReg[871])
);
LUT6 #(
   .INIT(64'b1001110000010101011011001110011101111011011110110010101111100011)  
) LUT6_1509 (
   .O(gates[1204]),
   .I0(gatesReg[1401]),
   .I1(gatesReg[423]),
   .I2(gatesReg[719]),
   .I3(gatesReg[1139]),
   .I4(gatesReg[1319]),
   .I5(gatesReg[1529])
);
LUT6 #(
   .INIT(64'b1110011011101111011001011111110100101011100101111111000111101100)  
) LUT6_1510 (
   .O(gates[70]),
   .I0(gatesReg[902]),
   .I1(gatesReg[1222]),
   .I2(gatesReg[827]),
   .I3(gatesReg[266]),
   .I4(gatesReg[1353]),
   .I5(gatesReg[174])
);
LUT6 #(
   .INIT(64'b1000110011110100011001111001101111101110011111110111101111101000)  
) LUT6_1511 (
   .O(gates[1047]),
   .I0(gatesReg[820]),
   .I1(gatesReg[422]),
   .I2(gatesReg[905]),
   .I3(gatesReg[1219]),
   .I4(gatesReg[1194]),
   .I5(gatesReg[1552])
);
LUT6 #(
   .INIT(64'b1000101111110001010011100010110100110111011000010011111110011000)  
) LUT6_1512 (
   .O(gates[839]),
   .I0(gatesReg[97]),
   .I1(gatesReg[41]),
   .I2(gatesReg[668]),
   .I3(gatesReg[52]),
   .I4(gatesReg[688]),
   .I5(gatesReg[750])
);
LUT6 #(
   .INIT(64'b1110001111111111101010110010111101111101110000101100110011010000)  
) LUT6_1513 (
   .O(gates[1055]),
   .I0(gatesReg[302]),
   .I1(gatesReg[1451]),
   .I2(gatesReg[1126]),
   .I3(gatesReg[774]),
   .I4(gatesReg[1453]),
   .I5(gatesReg[866])
);
LUT6 #(
   .INIT(64'b0010010111010110011001000001111110000010000000110111001111110001)  
) LUT6_1514 (
   .O(gates[1276]),
   .I0(gatesReg[910]),
   .I1(gatesReg[1341]),
   .I2(gatesReg[693]),
   .I3(gatesReg[770]),
   .I4(gatesReg[593]),
   .I5(gatesReg[188])
);
LUT6 #(
   .INIT(64'b0100111101011101001110100110011111111010010101000001100000111101)  
) LUT6_1515 (
   .O(gates[166]),
   .I0(gatesReg[402]),
   .I1(gatesReg[1534]),
   .I2(gatesReg[641]),
   .I3(gatesReg[1097]),
   .I4(gatesReg[893]),
   .I5(gatesReg[838])
);
LUT6 #(
   .INIT(64'b0111011010101110100111101111011100010111101110110110011000111110)  
) LUT6_1516 (
   .O(gates[88]),
   .I0(gatesReg[616]),
   .I1(gatesReg[640]),
   .I2(gatesReg[1121]),
   .I3(gatesReg[870]),
   .I4(gatesReg[804]),
   .I5(gatesReg[83])
);
LUT6 #(
   .INIT(64'b0110001101101000010001000110101110011000100000111000100010100001)  
) LUT6_1517 (
   .O(gates[1009]),
   .I0(gatesReg[1384]),
   .I1(gatesReg[896]),
   .I2(gatesReg[1468]),
   .I3(gatesReg[1385]),
   .I4(gatesReg[1464]),
   .I5(gatesReg[1494])
);
LUT6 #(
   .INIT(64'b0111001010111000001010000100000111111100000000101111101110011000)  
) LUT6_1518 (
   .O(gates[141]),
   .I0(gatesReg[962]),
   .I1(gatesReg[1085]),
   .I2(gatesReg[755]),
   .I3(gatesReg[777]),
   .I4(gatesReg[143]),
   .I5(gatesReg[464])
);
LUT6 #(
   .INIT(64'b1101110110010101111110001001000111010110000000110101000011010000)  
) LUT6_1519 (
   .O(gates[30]),
   .I0(gatesReg[1403]),
   .I1(gatesReg[6]),
   .I2(gatesReg[1051]),
   .I3(gatesReg[562]),
   .I4(gatesReg[1497]),
   .I5(gatesReg[1304])
);
LUT6 #(
   .INIT(64'b1101001101010100011110101111010110001101010011110111110110010010)  
) LUT6_1520 (
   .O(gates[909]),
   .I0(gatesReg[183]),
   .I1(gatesReg[497]),
   .I2(gatesReg[1102]),
   .I3(gatesReg[518]),
   .I4(gatesReg[1478]),
   .I5(gatesReg[439])
);
LUT6 #(
   .INIT(64'b0001101100110110110110001101101111101010010101000111010000100111)  
) LUT6_1521 (
   .O(gates[403]),
   .I0(gatesReg[1211]),
   .I1(gatesReg[362]),
   .I2(gatesReg[1379]),
   .I3(gatesReg[169]),
   .I4(gatesReg[411]),
   .I5(gatesReg[1542])
);
LUT6 #(
   .INIT(64'b1000011110110101101011101010010100000100101111100010011010100111)  
) LUT6_1522 (
   .O(gates[466]),
   .I0(gatesReg[705]),
   .I1(gatesReg[478]),
   .I2(gatesReg[398]),
   .I3(gatesReg[384]),
   .I4(gatesReg[836]),
   .I5(gatesReg[942])
);
LUT6 #(
   .INIT(64'b0110110011001001101100010100010110010011110011110101011111001010)  
) LUT6_1523 (
   .O(gates[1124]),
   .I0(gatesReg[955]),
   .I1(gatesReg[1376]),
   .I2(gatesReg[407]),
   .I3(gatesReg[18]),
   .I4(gatesReg[376]),
   .I5(gatesReg[912])
);
LUT6 #(
   .INIT(64'b0000101001011100111000100001101110110000100101101011011111010100)  
) LUT6_1524 (
   .O(gates[1230]),
   .I0(gatesReg[785]),
   .I1(gatesReg[1432]),
   .I2(gatesReg[599]),
   .I3(gatesReg[1167]),
   .I4(gatesReg[587]),
   .I5(gatesReg[1393])
);
LUT6 #(
   .INIT(64'b1011111000101001101000011011111000010110000001010101011000000101)  
) LUT6_1525 (
   .O(gates[134]),
   .I0(gatesReg[609]),
   .I1(gatesReg[1235]),
   .I2(gatesReg[190]),
   .I3(gatesReg[95]),
   .I4(gatesReg[298]),
   .I5(gatesReg[923])
);
LUT6 #(
   .INIT(64'b1111110000011001101110100011001010110011101111110110100001111100)  
) LUT6_1526 (
   .O(gates[75]),
   .I0(gatesReg[601]),
   .I1(gatesReg[822]),
   .I2(gatesReg[231]),
   .I3(gatesReg[243]),
   .I4(gatesReg[779]),
   .I5(gatesReg[551])
);
LUT6 #(
   .INIT(64'b1011111011001100011111101110001011100101010111111000010100001000)  
) LUT6_1527 (
   .O(gates[618]),
   .I0(gatesReg[148]),
   .I1(gatesReg[343]),
   .I2(gatesReg[504]),
   .I3(gatesReg[753]),
   .I4(gatesReg[1343]),
   .I5(gatesReg[697])
);
LUT6 #(
   .INIT(64'b1001010000110100010101110000100011110001110000101010111000011011)  
) LUT6_1528 (
   .O(gates[848]),
   .I0(gatesReg[981]),
   .I1(gatesReg[726]),
   .I2(gatesReg[857]),
   .I3(gatesReg[106]),
   .I4(gatesReg[1010]),
   .I5(gatesReg[707])
);
LUT6 #(
   .INIT(64'b1001101100010011101000011000111100001110011010101001010110010111)  
) LUT6_1529 (
   .O(gates[1163]),
   .I0(gatesReg[964]),
   .I1(gatesReg[157]),
   .I2(gatesReg[65]),
   .I3(gatesReg[935]),
   .I4(gatesReg[203]),
   .I5(gatesReg[261])
);
LUT6 #(
   .INIT(64'b0010100011101010000111000000001010101001101011111101101100110101)  
) LUT6_1530 (
   .O(gates[450]),
   .I0(gatesReg[1213]),
   .I1(gatesReg[1093]),
   .I2(gatesReg[1023]),
   .I3(gatesReg[81]),
   .I4(gatesReg[321]),
   .I5(gatesReg[1199])
);
LUT6 #(
   .INIT(64'b0000000100100010000110101111111100010010101111010101011010011000)  
) LUT6_1531 (
   .O(gates[1323]),
   .I0(gatesReg[624]),
   .I1(gatesReg[1300]),
   .I2(gatesReg[792]),
   .I3(gatesReg[86]),
   .I4(gatesReg[1158]),
   .I5(gatesReg[371])
);
LUT6 #(
   .INIT(64'b0100101001001001111001010000111010100110100011110101010100101001)  
) LUT6_1532 (
   .O(gates[1455]),
   .I0(gatesReg[656]),
   .I1(gatesReg[1079]),
   .I2(gatesReg[204]),
   .I3(gatesReg[1248]),
   .I4(gatesReg[1041]),
   .I5(gatesReg[435])
);
LUT6 #(
   .INIT(64'b0100010011100001001010000001001100100101010101010101000000000000)  
) LUT6_1533 (
   .O(gates[1405]),
   .I0(gatesReg[814]),
   .I1(gatesReg[1516]),
   .I2(gatesReg[1482]),
   .I3(gatesReg[924]),
   .I4(gatesReg[885]),
   .I5(gatesReg[884])
);
LUT6 #(
   .INIT(64'b1110010011000010110110110011101110110010000110101111000010111011)  
) LUT6_1534 (
   .O(gates[1060]),
   .I0(gatesReg[1412]),
   .I1(gatesReg[339]),
   .I2(gatesReg[760]),
   .I3(gatesReg[228]),
   .I4(gatesReg[863]),
   .I5(gatesReg[749])
);
LUT6 #(
   .INIT(64'b0111101011010000101010110111101011110111000111001000111010100001)  
) LUT6_1535 (
   .O(gates[1492]),
   .I0(gatesReg[531]),
   .I1(gatesReg[268]),
   .I2(gatesReg[829]),
   .I3(gatesReg[345]),
   .I4(gatesReg[172]),
   .I5(gatesReg[596])
);
LUT6 #(
   .INIT(64'b0000001001011001100110110000001011101001010010110001000011111011)  
) LUT6_1536 (
   .O(gates[703]),
   .I0(gatesReg[1297]),
   .I1(gatesReg[1521]),
   .I2(gatesReg[1366]),
   .I3(gatesReg[223]),
   .I4(gatesReg[613]),
   .I5(gatesReg[721])
);
LUT6 #(
   .INIT(64'b0000110011010101101111110010100111111101110011100001010100010100)  
) LUT6_1537 (
   .O(gates[900]),
   .I0(gatesReg[1043]),
   .I1(gatesReg[1255]),
   .I2(gatesReg[669]),
   .I3(gatesReg[282]),
   .I4(gatesReg[1082]),
   .I5(gatesReg[420])
);
LUT6 #(
   .INIT(64'b0101001100100001101101101000100010101011010100001100111011000101)  
) LUT6_1538 (
   .O(gates[1134]),
   .I0(gatesReg[121]),
   .I1(gatesReg[1066]),
   .I2(gatesReg[952]),
   .I3(gatesReg[639]),
   .I4(gatesReg[989]),
   .I5(gatesReg[494])
);
LUT6 #(
   .INIT(64'b1011100001011110010101011111110101011101001110000011001010110101)  
) LUT6_1539 (
   .O(gates[318]),
   .I0(gatesReg[1505]),
   .I1(gatesReg[487]),
   .I2(gatesReg[1071]),
   .I3(gatesReg[1348]),
   .I4(gatesReg[238]),
   .I5(gatesReg[873])
);
LUT6 #(
   .INIT(64'b1101011101110101101100100110001001101010010110110110111011001110)  
) LUT6_1540 (
   .O(gates[972]),
   .I0(gatesReg[577]),
   .I1(gatesReg[1137]),
   .I2(gatesReg[253]),
   .I3(gatesReg[448]),
   .I4(gatesReg[1227]),
   .I5(gatesReg[1417])
);
LUT6 #(
   .INIT(64'b0101110000111011001111010010110000100000111110001011101010100000)  
) LUT6_1541 (
   .O(gates[1100]),
   .I0(gatesReg[216]),
   .I1(gatesReg[852]),
   .I2(gatesReg[643]),
   .I3(gatesReg[63]),
   .I4(gatesReg[1120]),
   .I5(gatesReg[179])
);
LUT6 #(
   .INIT(64'b1011010001011000110011000011110010110000010100110000011101111111)  
) LUT6_1542 (
   .O(gates[473]),
   .I0(gatesReg[1532]),
   .I1(gatesReg[1475]),
   .I2(gatesReg[1105]),
   .I3(gatesReg[1187]),
   .I4(gatesReg[713]),
   .I5(gatesReg[676])
);
LUT6 #(
   .INIT(64'b0110100111100011010010000000110010101111011100001111010111110000)  
) LUT6_1543 (
   .O(gates[1377]),
   .I0(gatesReg[1334]),
   .I1(gatesReg[1251]),
   .I2(gatesReg[277]),
   .I3(gatesReg[1192]),
   .I4(gatesReg[879]),
   .I5(gatesReg[938])
);
LUT6 #(
   .INIT(64'b1111001111100000100101000111101111010110001011010000011101000011)  
) LUT6_1544 (
   .O(gates[1461]),
   .I0(gatesReg[1095]),
   .I1(gatesReg[1183]),
   .I2(gatesReg[1262]),
   .I3(gatesReg[1444]),
   .I4(gatesReg[1290]),
   .I5(gatesReg[1527])
);
LUT6 #(
   .INIT(64'b1000110100111011010110000111110000100100001110100011001010101101)  
) LUT6_1545 (
   .O(gates[185]),
   .I0(gatesReg[1132]),
   .I1(gatesReg[929]),
   .I2(gatesReg[133]),
   .I3(gatesReg[123]),
   .I4(gatesReg[304]),
   .I5(gatesReg[547])
);
LUT6 #(
   .INIT(64'b0110111110101001000000001100011010011001101001011010101001101011)  
) LUT6_1546 (
   .O(gates[3]),
   .I0(gatesReg[631]),
   .I1(gatesReg[1538]),
   .I2(gatesReg[1544]),
   .I3(gatesReg[396]),
   .I4(gatesReg[258]),
   .I5(gatesReg[1422])
);
LUT6 #(
   .INIT(64'b0101101111011011100110001011100111001110100111111110000001100010)  
) LUT6_1547 (
   .O(gates[248]),
   .I0(gatesReg[482]),
   .I1(gatesReg[949]),
   .I2(gatesReg[499]),
   .I3(gatesReg[56]),
   .I4(gatesReg[1369]),
   .I5(gatesReg[54])
);
LUT6 #(
   .INIT(64'b1100011100101001010001111111001000101111000111010101000100000100)  
) LUT6_1548 (
   .O(gates[146]),
   .I0(gatesReg[1151]),
   .I1(gatesReg[306]),
   .I2(gatesReg[1204]),
   .I3(gatesReg[70]),
   .I4(gatesReg[1047]),
   .I5(gatesReg[839])
);
LUT6 #(
   .INIT(64'b1010010111100110111101111011100001011011111110100011110001011111)  
) LUT6_1549 (
   .O(gates[1351]),
   .I0(gatesReg[1055]),
   .I1(gatesReg[1276]),
   .I2(gatesReg[166]),
   .I3(gatesReg[88]),
   .I4(gatesReg[1009]),
   .I5(gatesReg[141])
);
LUT6 #(
   .INIT(64'b0010110010010111100110000001010010110001100110010100111111100010)  
) LUT6_1550 (
   .O(gates[356]),
   .I0(gatesReg[30]),
   .I1(gatesReg[909]),
   .I2(gatesReg[403]),
   .I3(gatesReg[466]),
   .I4(gatesReg[1124]),
   .I5(gatesReg[1230])
);
LUT6 #(
   .INIT(64'b1111110001110100110110110110001010111000010000001010011010100011)  
) LUT6_1551 (
   .O(gates[802]),
   .I0(gatesReg[134]),
   .I1(gatesReg[75]),
   .I2(gatesReg[618]),
   .I3(gatesReg[848]),
   .I4(gatesReg[1163]),
   .I5(gatesReg[450])
);
LUT6 #(
   .INIT(64'b0011011111100111011001110110111001100000111001000101111010011011)  
) LUT6_1552 (
   .O(gates[4]),
   .I0(gatesReg[1323]),
   .I1(gatesReg[1455]),
   .I2(gatesReg[1405]),
   .I3(gatesReg[1060]),
   .I4(gatesReg[1492]),
   .I5(gatesReg[703])
);
LUT6 #(
   .INIT(64'b0000111101001100100011010111111100000011101010101110011000100010)  
) LUT6_1553 (
   .O(gates[528]),
   .I0(gatesReg[900]),
   .I1(gatesReg[1134]),
   .I2(gatesReg[318]),
   .I3(gatesReg[972]),
   .I4(gatesReg[1100]),
   .I5(gatesReg[473])
);
LUT6 #(
   .INIT(64'b0001111010000101100001000110011101011110110000011010010010100111)  
) LUT6_1554 (
   .O(gates[164]),
   .I0(gatesReg[1377]),
   .I1(gatesReg[1461]),
   .I2(gatesReg[185]),
   .I3(gatesReg[3]),
   .I4(gatesReg[248]),
   .I5(gatesReg[146])
);
LUT6 #(
   .INIT(64'b0000111010110101100010000110110011001001001011001110001100010110)  
) LUT6_1555 (
   .O(gates[807]),
   .I0(gatesReg[1351]),
   .I1(gatesReg[356]),
   .I2(gatesReg[802]),
   .I3(gatesReg[4]),
   .I4(gatesReg[528]),
   .I5(gatesReg[164])
);



endmodule