// 2014-8-29, 19:58:54

module mux_to7776_tree12(
                    input      [1727:0]data_in,
                    input                rx_fifo_clock,
                    input                rx_fifo_resetn,
                    input                valid,
                    output     [7775:0]data_out
                    );

     assign  data_out[0] = data_in[288];
     assign  data_out[1] = data_in[643];
     assign  data_out[2] = data_in[273];
     assign  data_out[3] = data_in[1407];
     assign  data_out[4] = data_in[1112];
     assign  data_out[5] = data_in[1284];
     assign  data_out[6] = data_in[406];
     assign  data_out[7] = data_in[390];
     assign  data_out[8] = data_in[1452];
     assign  data_out[9] = data_in[1340];
     assign  data_out[10] = data_in[908];
     assign  data_out[11] = data_in[753];
     assign  data_out[12] = data_in[406];
     assign  data_out[13] = data_in[1238];
     assign  data_out[14] = data_in[1272];
     assign  data_out[15] = data_in[830];
     assign  data_out[16] = data_in[1292];
     assign  data_out[17] = data_in[374];
     assign  data_out[18] = data_in[316];
     assign  data_out[19] = data_in[182];
     assign  data_out[20] = data_in[955];
     assign  data_out[21] = data_in[28];
     assign  data_out[22] = data_in[616];
     assign  data_out[23] = data_in[349];
     assign  data_out[24] = data_in[691];
     assign  data_out[25] = data_in[184];
     assign  data_out[26] = data_in[122];
     assign  data_out[27] = data_in[820];
     assign  data_out[28] = data_in[394];
     assign  data_out[29] = data_in[16];
     assign  data_out[30] = data_in[409];
     assign  data_out[31] = data_in[441];
     assign  data_out[32] = data_in[606];
     assign  data_out[33] = data_in[603];
     assign  data_out[34] = data_in[1348];
     assign  data_out[35] = data_in[1496];
     assign  data_out[36] = data_in[1724];
     assign  data_out[37] = data_in[620];
     assign  data_out[38] = data_in[1293];
     assign  data_out[39] = data_in[751];
     assign  data_out[40] = data_in[837];
     assign  data_out[41] = data_in[834];
     assign  data_out[42] = data_in[209];
     assign  data_out[43] = data_in[993];
     assign  data_out[44] = data_in[1395];
     assign  data_out[45] = data_in[1267];
     assign  data_out[46] = data_in[645];
     assign  data_out[47] = data_in[1435];
     assign  data_out[48] = data_in[1599];
     assign  data_out[49] = data_in[1645];
     assign  data_out[50] = data_in[536];
     assign  data_out[51] = data_in[511];
     assign  data_out[52] = data_in[917];
     assign  data_out[53] = data_in[1105];
     assign  data_out[54] = data_in[358];
     assign  data_out[55] = data_in[546];
     assign  data_out[56] = data_in[988];
     assign  data_out[57] = data_in[867];
     assign  data_out[58] = data_in[1368];
     assign  data_out[59] = data_in[1162];
     assign  data_out[60] = data_in[553];
     assign  data_out[61] = data_in[651];
     assign  data_out[62] = data_in[153];
     assign  data_out[63] = data_in[279];
     assign  data_out[64] = data_in[448];
     assign  data_out[65] = data_in[1200];
     assign  data_out[66] = data_in[1165];
     assign  data_out[67] = data_in[1682];
     assign  data_out[68] = data_in[995];
     assign  data_out[69] = data_in[210];
     assign  data_out[70] = data_in[608];
     assign  data_out[71] = data_in[1335];
     assign  data_out[72] = data_in[934];
     assign  data_out[73] = data_in[965];
     assign  data_out[74] = data_in[1383];
     assign  data_out[75] = data_in[1543];
     assign  data_out[76] = data_in[945];
     assign  data_out[77] = data_in[230];
     assign  data_out[78] = data_in[360];
     assign  data_out[79] = data_in[952];
     assign  data_out[80] = data_in[177];
     assign  data_out[81] = data_in[614];
     assign  data_out[82] = data_in[757];
     assign  data_out[83] = data_in[826];
     assign  data_out[84] = data_in[951];
     assign  data_out[85] = data_in[148];
     assign  data_out[86] = data_in[1292];
     assign  data_out[87] = data_in[1534];
     assign  data_out[88] = data_in[1373];
     assign  data_out[89] = data_in[819];
     assign  data_out[90] = data_in[1029];
     assign  data_out[91] = data_in[306];
     assign  data_out[92] = data_in[1421];
     assign  data_out[93] = data_in[908];
     assign  data_out[94] = data_in[983];
     assign  data_out[95] = data_in[469];
     assign  data_out[96] = data_in[508];
     assign  data_out[97] = data_in[779];
     assign  data_out[98] = data_in[1662];
     assign  data_out[99] = data_in[29];
     assign  data_out[100] = data_in[1709];
     assign  data_out[101] = data_in[784];
     assign  data_out[102] = data_in[56];
     assign  data_out[103] = data_in[915];
     assign  data_out[104] = data_in[670];
     assign  data_out[105] = data_in[199];
     assign  data_out[106] = data_in[823];
     assign  data_out[107] = data_in[1562];
     assign  data_out[108] = data_in[285];
     assign  data_out[109] = data_in[56];
     assign  data_out[110] = data_in[244];
     assign  data_out[111] = data_in[329];
     assign  data_out[112] = data_in[1529];
     assign  data_out[113] = data_in[1483];
     assign  data_out[114] = data_in[896];
     assign  data_out[115] = data_in[83];
     assign  data_out[116] = data_in[1164];
     assign  data_out[117] = data_in[719];
     assign  data_out[118] = data_in[72];
     assign  data_out[119] = data_in[1681];
     assign  data_out[120] = data_in[259];
     assign  data_out[121] = data_in[45];
     assign  data_out[122] = data_in[1249];
     assign  data_out[123] = data_in[893];
     assign  data_out[124] = data_in[689];
     assign  data_out[125] = data_in[1230];
     assign  data_out[126] = data_in[270];
     assign  data_out[127] = data_in[688];
     assign  data_out[128] = data_in[457];
     assign  data_out[129] = data_in[763];
     assign  data_out[130] = data_in[732];
     assign  data_out[131] = data_in[1569];
     assign  data_out[132] = data_in[1301];
     assign  data_out[133] = data_in[98];
     assign  data_out[134] = data_in[1612];
     assign  data_out[135] = data_in[911];
     assign  data_out[136] = data_in[1402];
     assign  data_out[137] = data_in[81];
     assign  data_out[138] = data_in[1240];
     assign  data_out[139] = data_in[260];
     assign  data_out[140] = data_in[482];
     assign  data_out[141] = data_in[1431];
     assign  data_out[142] = data_in[396];
     assign  data_out[143] = data_in[1431];
     assign  data_out[144] = data_in[492];
     assign  data_out[145] = data_in[1167];
     assign  data_out[146] = data_in[274];
     assign  data_out[147] = data_in[749];
     assign  data_out[148] = data_in[1504];
     assign  data_out[149] = data_in[1685];
     assign  data_out[150] = data_in[537];
     assign  data_out[151] = data_in[275];
     assign  data_out[152] = data_in[219];
     assign  data_out[153] = data_in[1630];
     assign  data_out[154] = data_in[123];
     assign  data_out[155] = data_in[436];
     assign  data_out[156] = data_in[1070];
     assign  data_out[157] = data_in[820];
     assign  data_out[158] = data_in[839];
     assign  data_out[159] = data_in[1532];
     assign  data_out[160] = data_in[666];
     assign  data_out[161] = data_in[469];
     assign  data_out[162] = data_in[856];
     assign  data_out[163] = data_in[1017];
     assign  data_out[164] = data_in[499];
     assign  data_out[165] = data_in[1580];
     assign  data_out[166] = data_in[609];
     assign  data_out[167] = data_in[206];
     assign  data_out[168] = data_in[4];
     assign  data_out[169] = data_in[49];
     assign  data_out[170] = data_in[1294];
     assign  data_out[171] = data_in[362];
     assign  data_out[172] = data_in[713];
     assign  data_out[173] = data_in[345];
     assign  data_out[174] = data_in[1184];
     assign  data_out[175] = data_in[128];
     assign  data_out[176] = data_in[1244];
     assign  data_out[177] = data_in[1386];
     assign  data_out[178] = data_in[1075];
     assign  data_out[179] = data_in[158];
     assign  data_out[180] = data_in[27];
     assign  data_out[181] = data_in[666];
     assign  data_out[182] = data_in[1611];
     assign  data_out[183] = data_in[976];
     assign  data_out[184] = data_in[1070];
     assign  data_out[185] = data_in[1366];
     assign  data_out[186] = data_in[333];
     assign  data_out[187] = data_in[1683];
     assign  data_out[188] = data_in[1661];
     assign  data_out[189] = data_in[1094];
     assign  data_out[190] = data_in[601];
     assign  data_out[191] = data_in[1059];
     assign  data_out[192] = data_in[482];
     assign  data_out[193] = data_in[564];
     assign  data_out[194] = data_in[464];
     assign  data_out[195] = data_in[58];
     assign  data_out[196] = data_in[1600];
     assign  data_out[197] = data_in[504];
     assign  data_out[198] = data_in[1289];
     assign  data_out[199] = data_in[325];
     assign  data_out[200] = data_in[967];
     assign  data_out[201] = data_in[892];
     assign  data_out[202] = data_in[779];
     assign  data_out[203] = data_in[1186];
     assign  data_out[204] = data_in[1721];
     assign  data_out[205] = data_in[186];
     assign  data_out[206] = data_in[1518];
     assign  data_out[207] = data_in[122];
     assign  data_out[208] = data_in[27];
     assign  data_out[209] = data_in[25];
     assign  data_out[210] = data_in[1433];
     assign  data_out[211] = data_in[884];
     assign  data_out[212] = data_in[1539];
     assign  data_out[213] = data_in[957];
     assign  data_out[214] = data_in[758];
     assign  data_out[215] = data_in[1450];
     assign  data_out[216] = data_in[1606];
     assign  data_out[217] = data_in[1582];
     assign  data_out[218] = data_in[514];
     assign  data_out[219] = data_in[525];
     assign  data_out[220] = data_in[1395];
     assign  data_out[221] = data_in[498];
     assign  data_out[222] = data_in[1195];
     assign  data_out[223] = data_in[1702];
     assign  data_out[224] = data_in[1679];
     assign  data_out[225] = data_in[1336];
     assign  data_out[226] = data_in[850];
     assign  data_out[227] = data_in[428];
     assign  data_out[228] = data_in[1552];
     assign  data_out[229] = data_in[1270];
     assign  data_out[230] = data_in[1254];
     assign  data_out[231] = data_in[260];
     assign  data_out[232] = data_in[840];
     assign  data_out[233] = data_in[1291];
     assign  data_out[234] = data_in[624];
     assign  data_out[235] = data_in[381];
     assign  data_out[236] = data_in[631];
     assign  data_out[237] = data_in[1370];
     assign  data_out[238] = data_in[579];
     assign  data_out[239] = data_in[848];
     assign  data_out[240] = data_in[694];
     assign  data_out[241] = data_in[1505];
     assign  data_out[242] = data_in[617];
     assign  data_out[243] = data_in[373];
     assign  data_out[244] = data_in[316];
     assign  data_out[245] = data_in[1152];
     assign  data_out[246] = data_in[899];
     assign  data_out[247] = data_in[282];
     assign  data_out[248] = data_in[1319];
     assign  data_out[249] = data_in[770];
     assign  data_out[250] = data_in[432];
     assign  data_out[251] = data_in[1548];
     assign  data_out[252] = data_in[773];
     assign  data_out[253] = data_in[1420];
     assign  data_out[254] = data_in[1070];
     assign  data_out[255] = data_in[1627];
     assign  data_out[256] = data_in[1551];
     assign  data_out[257] = data_in[970];
     assign  data_out[258] = data_in[984];
     assign  data_out[259] = data_in[461];
     assign  data_out[260] = data_in[600];
     assign  data_out[261] = data_in[124];
     assign  data_out[262] = data_in[102];
     assign  data_out[263] = data_in[1645];
     assign  data_out[264] = data_in[334];
     assign  data_out[265] = data_in[1281];
     assign  data_out[266] = data_in[1164];
     assign  data_out[267] = data_in[829];
     assign  data_out[268] = data_in[1317];
     assign  data_out[269] = data_in[1346];
     assign  data_out[270] = data_in[1273];
     assign  data_out[271] = data_in[931];
     assign  data_out[272] = data_in[890];
     assign  data_out[273] = data_in[1227];
     assign  data_out[274] = data_in[757];
     assign  data_out[275] = data_in[1304];
     assign  data_out[276] = data_in[842];
     assign  data_out[277] = data_in[331];
     assign  data_out[278] = data_in[40];
     assign  data_out[279] = data_in[431];
     assign  data_out[280] = data_in[407];
     assign  data_out[281] = data_in[502];
     assign  data_out[282] = data_in[989];
     assign  data_out[283] = data_in[752];
     assign  data_out[284] = data_in[132];
     assign  data_out[285] = data_in[1551];
     assign  data_out[286] = data_in[676];
     assign  data_out[287] = data_in[1646];
     assign  data_out[288] = data_in[1550];
     assign  data_out[289] = data_in[725];
     assign  data_out[290] = data_in[972];
     assign  data_out[291] = data_in[275];
     assign  data_out[292] = data_in[552];
     assign  data_out[293] = data_in[708];
     assign  data_out[294] = data_in[1157];
     assign  data_out[295] = data_in[123];
     assign  data_out[296] = data_in[860];
     assign  data_out[297] = data_in[514];
     assign  data_out[298] = data_in[411];
     assign  data_out[299] = data_in[285];
     assign  data_out[300] = data_in[582];
     assign  data_out[301] = data_in[1501];
     assign  data_out[302] = data_in[1592];
     assign  data_out[303] = data_in[1642];
     assign  data_out[304] = data_in[691];
     assign  data_out[305] = data_in[1128];
     assign  data_out[306] = data_in[1660];
     assign  data_out[307] = data_in[1231];
     assign  data_out[308] = data_in[524];
     assign  data_out[309] = data_in[1517];
     assign  data_out[310] = data_in[1641];
     assign  data_out[311] = data_in[590];
     assign  data_out[312] = data_in[1495];
     assign  data_out[313] = data_in[243];
     assign  data_out[314] = data_in[765];
     assign  data_out[315] = data_in[1101];
     assign  data_out[316] = data_in[1377];
     assign  data_out[317] = data_in[796];
     assign  data_out[318] = data_in[734];
     assign  data_out[319] = data_in[32];
     assign  data_out[320] = data_in[374];
     assign  data_out[321] = data_in[1486];
     assign  data_out[322] = data_in[326];
     assign  data_out[323] = data_in[41];
     assign  data_out[324] = data_in[1328];
     assign  data_out[325] = data_in[241];
     assign  data_out[326] = data_in[1103];
     assign  data_out[327] = data_in[893];
     assign  data_out[328] = data_in[1075];
     assign  data_out[329] = data_in[1724];
     assign  data_out[330] = data_in[968];
     assign  data_out[331] = data_in[14];
     assign  data_out[332] = data_in[246];
     assign  data_out[333] = data_in[255];
     assign  data_out[334] = data_in[1527];
     assign  data_out[335] = data_in[1714];
     assign  data_out[336] = data_in[872];
     assign  data_out[337] = data_in[1038];
     assign  data_out[338] = data_in[812];
     assign  data_out[339] = data_in[1216];
     assign  data_out[340] = data_in[65];
     assign  data_out[341] = data_in[1307];
     assign  data_out[342] = data_in[791];
     assign  data_out[343] = data_in[368];
     assign  data_out[344] = data_in[1000];
     assign  data_out[345] = data_in[810];
     assign  data_out[346] = data_in[1201];
     assign  data_out[347] = data_in[431];
     assign  data_out[348] = data_in[1064];
     assign  data_out[349] = data_in[1271];
     assign  data_out[350] = data_in[503];
     assign  data_out[351] = data_in[1163];
     assign  data_out[352] = data_in[879];
     assign  data_out[353] = data_in[300];
     assign  data_out[354] = data_in[1417];
     assign  data_out[355] = data_in[1711];
     assign  data_out[356] = data_in[957];
     assign  data_out[357] = data_in[1611];
     assign  data_out[358] = data_in[349];
     assign  data_out[359] = data_in[1432];
     assign  data_out[360] = data_in[337];
     assign  data_out[361] = data_in[353];
     assign  data_out[362] = data_in[1388];
     assign  data_out[363] = data_in[1334];
     assign  data_out[364] = data_in[244];
     assign  data_out[365] = data_in[1698];
     assign  data_out[366] = data_in[1338];
     assign  data_out[367] = data_in[798];
     assign  data_out[368] = data_in[1185];
     assign  data_out[369] = data_in[408];
     assign  data_out[370] = data_in[290];
     assign  data_out[371] = data_in[645];
     assign  data_out[372] = data_in[6];
     assign  data_out[373] = data_in[240];
     assign  data_out[374] = data_in[1490];
     assign  data_out[375] = data_in[294];
     assign  data_out[376] = data_in[1223];
     assign  data_out[377] = data_in[911];
     assign  data_out[378] = data_in[1417];
     assign  data_out[379] = data_in[88];
     assign  data_out[380] = data_in[775];
     assign  data_out[381] = data_in[397];
     assign  data_out[382] = data_in[1244];
     assign  data_out[383] = data_in[1692];
     assign  data_out[384] = data_in[1437];
     assign  data_out[385] = data_in[751];
     assign  data_out[386] = data_in[840];
     assign  data_out[387] = data_in[380];
     assign  data_out[388] = data_in[764];
     assign  data_out[389] = data_in[1280];
     assign  data_out[390] = data_in[1301];
     assign  data_out[391] = data_in[136];
     assign  data_out[392] = data_in[437];
     assign  data_out[393] = data_in[105];
     assign  data_out[394] = data_in[1356];
     assign  data_out[395] = data_in[433];
     assign  data_out[396] = data_in[347];
     assign  data_out[397] = data_in[37];
     assign  data_out[398] = data_in[1554];
     assign  data_out[399] = data_in[1192];
     assign  data_out[400] = data_in[354];
     assign  data_out[401] = data_in[41];
     assign  data_out[402] = data_in[1576];
     assign  data_out[403] = data_in[689];
     assign  data_out[404] = data_in[724];
     assign  data_out[405] = data_in[1069];
     assign  data_out[406] = data_in[1096];
     assign  data_out[407] = data_in[88];
     assign  data_out[408] = data_in[1714];
     assign  data_out[409] = data_in[606];
     assign  data_out[410] = data_in[1666];
     assign  data_out[411] = data_in[1470];
     assign  data_out[412] = data_in[200];
     assign  data_out[413] = data_in[1265];
     assign  data_out[414] = data_in[1029];
     assign  data_out[415] = data_in[918];
     assign  data_out[416] = data_in[1125];
     assign  data_out[417] = data_in[860];
     assign  data_out[418] = data_in[1510];
     assign  data_out[419] = data_in[1565];
     assign  data_out[420] = data_in[180];
     assign  data_out[421] = data_in[1378];
     assign  data_out[422] = data_in[1452];
     assign  data_out[423] = data_in[1503];
     assign  data_out[424] = data_in[409];
     assign  data_out[425] = data_in[851];
     assign  data_out[426] = data_in[1693];
     assign  data_out[427] = data_in[466];
     assign  data_out[428] = data_in[162];
     assign  data_out[429] = data_in[333];
     assign  data_out[430] = data_in[1250];
     assign  data_out[431] = data_in[927];
     assign  data_out[432] = data_in[1261];
     assign  data_out[433] = data_in[361];
     assign  data_out[434] = data_in[374];
     assign  data_out[435] = data_in[843];
     assign  data_out[436] = data_in[709];
     assign  data_out[437] = data_in[120];
     assign  data_out[438] = data_in[693];
     assign  data_out[439] = data_in[386];
     assign  data_out[440] = data_in[993];
     assign  data_out[441] = data_in[1305];
     assign  data_out[442] = data_in[1608];
     assign  data_out[443] = data_in[848];
     assign  data_out[444] = data_in[593];
     assign  data_out[445] = data_in[540];
     assign  data_out[446] = data_in[1658];
     assign  data_out[447] = data_in[790];
     assign  data_out[448] = data_in[1448];
     assign  data_out[449] = data_in[1725];
     assign  data_out[450] = data_in[561];
     assign  data_out[451] = data_in[469];
     assign  data_out[452] = data_in[206];
     assign  data_out[453] = data_in[1069];
     assign  data_out[454] = data_in[292];
     assign  data_out[455] = data_in[580];
     assign  data_out[456] = data_in[1718];
     assign  data_out[457] = data_in[356];
     assign  data_out[458] = data_in[899];
     assign  data_out[459] = data_in[1185];
     assign  data_out[460] = data_in[866];
     assign  data_out[461] = data_in[1221];
     assign  data_out[462] = data_in[1494];
     assign  data_out[463] = data_in[679];
     assign  data_out[464] = data_in[580];
     assign  data_out[465] = data_in[1413];
     assign  data_out[466] = data_in[433];
     assign  data_out[467] = data_in[659];
     assign  data_out[468] = data_in[14];
     assign  data_out[469] = data_in[1118];
     assign  data_out[470] = data_in[1634];
     assign  data_out[471] = data_in[1014];
     assign  data_out[472] = data_in[14];
     assign  data_out[473] = data_in[583];
     assign  data_out[474] = data_in[309];
     assign  data_out[475] = data_in[1456];
     assign  data_out[476] = data_in[1321];
     assign  data_out[477] = data_in[554];
     assign  data_out[478] = data_in[16];
     assign  data_out[479] = data_in[713];
     assign  data_out[480] = data_in[1159];
     assign  data_out[481] = data_in[612];
     assign  data_out[482] = data_in[1446];
     assign  data_out[483] = data_in[988];
     assign  data_out[484] = data_in[1680];
     assign  data_out[485] = data_in[1727];
     assign  data_out[486] = data_in[1040];
     assign  data_out[487] = data_in[245];
     assign  data_out[488] = data_in[1348];
     assign  data_out[489] = data_in[1190];
     assign  data_out[490] = data_in[332];
     assign  data_out[491] = data_in[669];
     assign  data_out[492] = data_in[15];
     assign  data_out[493] = data_in[94];
     assign  data_out[494] = data_in[171];
     assign  data_out[495] = data_in[315];
     assign  data_out[496] = data_in[870];
     assign  data_out[497] = data_in[1137];
     assign  data_out[498] = data_in[1454];
     assign  data_out[499] = data_in[1467];
     assign  data_out[500] = data_in[260];
     assign  data_out[501] = data_in[1361];
     assign  data_out[502] = data_in[359];
     assign  data_out[503] = data_in[989];
     assign  data_out[504] = data_in[431];
     assign  data_out[505] = data_in[821];
     assign  data_out[506] = data_in[1424];
     assign  data_out[507] = data_in[1400];
     assign  data_out[508] = data_in[1588];
     assign  data_out[509] = data_in[672];
     assign  data_out[510] = data_in[170];
     assign  data_out[511] = data_in[1016];
     assign  data_out[512] = data_in[1438];
     assign  data_out[513] = data_in[1321];
     assign  data_out[514] = data_in[112];
     assign  data_out[515] = data_in[163];
     assign  data_out[516] = data_in[91];
     assign  data_out[517] = data_in[30];
     assign  data_out[518] = data_in[269];
     assign  data_out[519] = data_in[837];
     assign  data_out[520] = data_in[440];
     assign  data_out[521] = data_in[361];
     assign  data_out[522] = data_in[761];
     assign  data_out[523] = data_in[505];
     assign  data_out[524] = data_in[189];
     assign  data_out[525] = data_in[16];
     assign  data_out[526] = data_in[619];
     assign  data_out[527] = data_in[622];
     assign  data_out[528] = data_in[206];
     assign  data_out[529] = data_in[552];
     assign  data_out[530] = data_in[815];
     assign  data_out[531] = data_in[1197];
     assign  data_out[532] = data_in[1178];
     assign  data_out[533] = data_in[363];
     assign  data_out[534] = data_in[491];
     assign  data_out[535] = data_in[245];
     assign  data_out[536] = data_in[1143];
     assign  data_out[537] = data_in[567];
     assign  data_out[538] = data_in[1102];
     assign  data_out[539] = data_in[567];
     assign  data_out[540] = data_in[435];
     assign  data_out[541] = data_in[745];
     assign  data_out[542] = data_in[1274];
     assign  data_out[543] = data_in[1212];
     assign  data_out[544] = data_in[714];
     assign  data_out[545] = data_in[358];
     assign  data_out[546] = data_in[552];
     assign  data_out[547] = data_in[268];
     assign  data_out[548] = data_in[1139];
     assign  data_out[549] = data_in[54];
     assign  data_out[550] = data_in[8];
     assign  data_out[551] = data_in[159];
     assign  data_out[552] = data_in[837];
     assign  data_out[553] = data_in[1412];
     assign  data_out[554] = data_in[630];
     assign  data_out[555] = data_in[608];
     assign  data_out[556] = data_in[347];
     assign  data_out[557] = data_in[1080];
     assign  data_out[558] = data_in[1263];
     assign  data_out[559] = data_in[1574];
     assign  data_out[560] = data_in[823];
     assign  data_out[561] = data_in[298];
     assign  data_out[562] = data_in[484];
     assign  data_out[563] = data_in[1289];
     assign  data_out[564] = data_in[608];
     assign  data_out[565] = data_in[1578];
     assign  data_out[566] = data_in[736];
     assign  data_out[567] = data_in[1364];
     assign  data_out[568] = data_in[25];
     assign  data_out[569] = data_in[1446];
     assign  data_out[570] = data_in[84];
     assign  data_out[571] = data_in[627];
     assign  data_out[572] = data_in[200];
     assign  data_out[573] = data_in[1109];
     assign  data_out[574] = data_in[1024];
     assign  data_out[575] = data_in[10];
     assign  data_out[576] = data_in[1571];
     assign  data_out[577] = data_in[769];
     assign  data_out[578] = data_in[981];
     assign  data_out[579] = data_in[180];
     assign  data_out[580] = data_in[1718];
     assign  data_out[581] = data_in[1177];
     assign  data_out[582] = data_in[828];
     assign  data_out[583] = data_in[385];
     assign  data_out[584] = data_in[1628];
     assign  data_out[585] = data_in[596];
     assign  data_out[586] = data_in[1245];
     assign  data_out[587] = data_in[947];
     assign  data_out[588] = data_in[1017];
     assign  data_out[589] = data_in[409];
     assign  data_out[590] = data_in[797];
     assign  data_out[591] = data_in[607];
     assign  data_out[592] = data_in[475];
     assign  data_out[593] = data_in[636];
     assign  data_out[594] = data_in[107];
     assign  data_out[595] = data_in[1509];
     assign  data_out[596] = data_in[1412];
     assign  data_out[597] = data_in[307];
     assign  data_out[598] = data_in[73];
     assign  data_out[599] = data_in[932];
     assign  data_out[600] = data_in[837];
     assign  data_out[601] = data_in[1250];
     assign  data_out[602] = data_in[242];
     assign  data_out[603] = data_in[1574];
     assign  data_out[604] = data_in[1327];
     assign  data_out[605] = data_in[857];
     assign  data_out[606] = data_in[839];
     assign  data_out[607] = data_in[489];
     assign  data_out[608] = data_in[386];
     assign  data_out[609] = data_in[33];
     assign  data_out[610] = data_in[749];
     assign  data_out[611] = data_in[556];
     assign  data_out[612] = data_in[290];
     assign  data_out[613] = data_in[1535];
     assign  data_out[614] = data_in[114];
     assign  data_out[615] = data_in[1154];
     assign  data_out[616] = data_in[876];
     assign  data_out[617] = data_in[698];
     assign  data_out[618] = data_in[1590];
     assign  data_out[619] = data_in[1544];
     assign  data_out[620] = data_in[836];
     assign  data_out[621] = data_in[797];
     assign  data_out[622] = data_in[1641];
     assign  data_out[623] = data_in[1262];
     assign  data_out[624] = data_in[1071];
     assign  data_out[625] = data_in[1450];
     assign  data_out[626] = data_in[464];
     assign  data_out[627] = data_in[1677];
     assign  data_out[628] = data_in[1107];
     assign  data_out[629] = data_in[977];
     assign  data_out[630] = data_in[1206];
     assign  data_out[631] = data_in[1636];
     assign  data_out[632] = data_in[1129];
     assign  data_out[633] = data_in[849];
     assign  data_out[634] = data_in[1128];
     assign  data_out[635] = data_in[3];
     assign  data_out[636] = data_in[644];
     assign  data_out[637] = data_in[1300];
     assign  data_out[638] = data_in[685];
     assign  data_out[639] = data_in[1462];
     assign  data_out[640] = data_in[1149];
     assign  data_out[641] = data_in[438];
     assign  data_out[642] = data_in[337];
     assign  data_out[643] = data_in[377];
     assign  data_out[644] = data_in[339];
     assign  data_out[645] = data_in[1477];
     assign  data_out[646] = data_in[705];
     assign  data_out[647] = data_in[1293];
     assign  data_out[648] = data_in[803];
     assign  data_out[649] = data_in[672];
     assign  data_out[650] = data_in[56];
     assign  data_out[651] = data_in[747];
     assign  data_out[652] = data_in[6];
     assign  data_out[653] = data_in[338];
     assign  data_out[654] = data_in[1302];
     assign  data_out[655] = data_in[1084];
     assign  data_out[656] = data_in[41];
     assign  data_out[657] = data_in[519];
     assign  data_out[658] = data_in[13];
     assign  data_out[659] = data_in[1667];
     assign  data_out[660] = data_in[502];
     assign  data_out[661] = data_in[1588];
     assign  data_out[662] = data_in[196];
     assign  data_out[663] = data_in[173];
     assign  data_out[664] = data_in[881];
     assign  data_out[665] = data_in[734];
     assign  data_out[666] = data_in[1700];
     assign  data_out[667] = data_in[1201];
     assign  data_out[668] = data_in[2];
     assign  data_out[669] = data_in[773];
     assign  data_out[670] = data_in[793];
     assign  data_out[671] = data_in[935];
     assign  data_out[672] = data_in[1639];
     assign  data_out[673] = data_in[437];
     assign  data_out[674] = data_in[1364];
     assign  data_out[675] = data_in[409];
     assign  data_out[676] = data_in[0];
     assign  data_out[677] = data_in[110];
     assign  data_out[678] = data_in[525];
     assign  data_out[679] = data_in[547];
     assign  data_out[680] = data_in[876];
     assign  data_out[681] = data_in[820];
     assign  data_out[682] = data_in[1353];
     assign  data_out[683] = data_in[414];
     assign  data_out[684] = data_in[298];
     assign  data_out[685] = data_in[1070];
     assign  data_out[686] = data_in[1011];
     assign  data_out[687] = data_in[262];
     assign  data_out[688] = data_in[699];
     assign  data_out[689] = data_in[426];
     assign  data_out[690] = data_in[74];
     assign  data_out[691] = data_in[1406];
     assign  data_out[692] = data_in[248];
     assign  data_out[693] = data_in[627];
     assign  data_out[694] = data_in[287];
     assign  data_out[695] = data_in[1067];
     assign  data_out[696] = data_in[776];
     assign  data_out[697] = data_in[1018];
     assign  data_out[698] = data_in[321];
     assign  data_out[699] = data_in[140];
     assign  data_out[700] = data_in[1088];
     assign  data_out[701] = data_in[1558];
     assign  data_out[702] = data_in[1667];
     assign  data_out[703] = data_in[1285];
     assign  data_out[704] = data_in[337];
     assign  data_out[705] = data_in[1560];
     assign  data_out[706] = data_in[1397];
     assign  data_out[707] = data_in[1471];
     assign  data_out[708] = data_in[707];
     assign  data_out[709] = data_in[486];
     assign  data_out[710] = data_in[1225];
     assign  data_out[711] = data_in[1308];
     assign  data_out[712] = data_in[1263];
     assign  data_out[713] = data_in[1066];
     assign  data_out[714] = data_in[953];
     assign  data_out[715] = data_in[731];
     assign  data_out[716] = data_in[1588];
     assign  data_out[717] = data_in[332];
     assign  data_out[718] = data_in[544];
     assign  data_out[719] = data_in[1635];
     assign  data_out[720] = data_in[150];
     assign  data_out[721] = data_in[1650];
     assign  data_out[722] = data_in[1373];
     assign  data_out[723] = data_in[877];
     assign  data_out[724] = data_in[830];
     assign  data_out[725] = data_in[523];
     assign  data_out[726] = data_in[1537];
     assign  data_out[727] = data_in[1120];
     assign  data_out[728] = data_in[470];
     assign  data_out[729] = data_in[1437];
     assign  data_out[730] = data_in[1673];
     assign  data_out[731] = data_in[489];
     assign  data_out[732] = data_in[245];
     assign  data_out[733] = data_in[1237];
     assign  data_out[734] = data_in[625];
     assign  data_out[735] = data_in[624];
     assign  data_out[736] = data_in[1612];
     assign  data_out[737] = data_in[1505];
     assign  data_out[738] = data_in[864];
     assign  data_out[739] = data_in[980];
     assign  data_out[740] = data_in[273];
     assign  data_out[741] = data_in[955];
     assign  data_out[742] = data_in[1271];
     assign  data_out[743] = data_in[1703];
     assign  data_out[744] = data_in[1108];
     assign  data_out[745] = data_in[957];
     assign  data_out[746] = data_in[651];
     assign  data_out[747] = data_in[206];
     assign  data_out[748] = data_in[140];
     assign  data_out[749] = data_in[1133];
     assign  data_out[750] = data_in[1672];
     assign  data_out[751] = data_in[318];
     assign  data_out[752] = data_in[1384];
     assign  data_out[753] = data_in[834];
     assign  data_out[754] = data_in[586];
     assign  data_out[755] = data_in[115];
     assign  data_out[756] = data_in[844];
     assign  data_out[757] = data_in[734];
     assign  data_out[758] = data_in[817];
     assign  data_out[759] = data_in[1508];
     assign  data_out[760] = data_in[320];
     assign  data_out[761] = data_in[1348];
     assign  data_out[762] = data_in[1204];
     assign  data_out[763] = data_in[785];
     assign  data_out[764] = data_in[564];
     assign  data_out[765] = data_in[1335];
     assign  data_out[766] = data_in[438];
     assign  data_out[767] = data_in[1438];
     assign  data_out[768] = data_in[165];
     assign  data_out[769] = data_in[1047];
     assign  data_out[770] = data_in[1328];
     assign  data_out[771] = data_in[1590];
     assign  data_out[772] = data_in[1532];
     assign  data_out[773] = data_in[355];
     assign  data_out[774] = data_in[1124];
     assign  data_out[775] = data_in[773];
     assign  data_out[776] = data_in[257];
     assign  data_out[777] = data_in[1389];
     assign  data_out[778] = data_in[1644];
     assign  data_out[779] = data_in[862];
     assign  data_out[780] = data_in[691];
     assign  data_out[781] = data_in[57];
     assign  data_out[782] = data_in[1253];
     assign  data_out[783] = data_in[984];
     assign  data_out[784] = data_in[1183];
     assign  data_out[785] = data_in[1157];
     assign  data_out[786] = data_in[708];
     assign  data_out[787] = data_in[939];
     assign  data_out[788] = data_in[452];
     assign  data_out[789] = data_in[1206];
     assign  data_out[790] = data_in[454];
     assign  data_out[791] = data_in[871];
     assign  data_out[792] = data_in[1387];
     assign  data_out[793] = data_in[1459];
     assign  data_out[794] = data_in[678];
     assign  data_out[795] = data_in[1346];
     assign  data_out[796] = data_in[1519];
     assign  data_out[797] = data_in[405];
     assign  data_out[798] = data_in[690];
     assign  data_out[799] = data_in[221];
     assign  data_out[800] = data_in[40];
     assign  data_out[801] = data_in[582];
     assign  data_out[802] = data_in[303];
     assign  data_out[803] = data_in[827];
     assign  data_out[804] = data_in[246];
     assign  data_out[805] = data_in[1466];
     assign  data_out[806] = data_in[1518];
     assign  data_out[807] = data_in[210];
     assign  data_out[808] = data_in[984];
     assign  data_out[809] = data_in[1153];
     assign  data_out[810] = data_in[1081];
     assign  data_out[811] = data_in[1315];
     assign  data_out[812] = data_in[906];
     assign  data_out[813] = data_in[1085];
     assign  data_out[814] = data_in[1601];
     assign  data_out[815] = data_in[583];
     assign  data_out[816] = data_in[484];
     assign  data_out[817] = data_in[233];
     assign  data_out[818] = data_in[682];
     assign  data_out[819] = data_in[35];
     assign  data_out[820] = data_in[1384];
     assign  data_out[821] = data_in[641];
     assign  data_out[822] = data_in[1315];
     assign  data_out[823] = data_in[493];
     assign  data_out[824] = data_in[250];
     assign  data_out[825] = data_in[371];
     assign  data_out[826] = data_in[1268];
     assign  data_out[827] = data_in[820];
     assign  data_out[828] = data_in[694];
     assign  data_out[829] = data_in[943];
     assign  data_out[830] = data_in[1239];
     assign  data_out[831] = data_in[1292];
     assign  data_out[832] = data_in[798];
     assign  data_out[833] = data_in[130];
     assign  data_out[834] = data_in[1619];
     assign  data_out[835] = data_in[1452];
     assign  data_out[836] = data_in[656];
     assign  data_out[837] = data_in[642];
     assign  data_out[838] = data_in[1727];
     assign  data_out[839] = data_in[892];
     assign  data_out[840] = data_in[1082];
     assign  data_out[841] = data_in[390];
     assign  data_out[842] = data_in[700];
     assign  data_out[843] = data_in[239];
     assign  data_out[844] = data_in[17];
     assign  data_out[845] = data_in[43];
     assign  data_out[846] = data_in[113];
     assign  data_out[847] = data_in[441];
     assign  data_out[848] = data_in[929];
     assign  data_out[849] = data_in[487];
     assign  data_out[850] = data_in[586];
     assign  data_out[851] = data_in[1059];
     assign  data_out[852] = data_in[22];
     assign  data_out[853] = data_in[1683];
     assign  data_out[854] = data_in[1083];
     assign  data_out[855] = data_in[849];
     assign  data_out[856] = data_in[1100];
     assign  data_out[857] = data_in[1492];
     assign  data_out[858] = data_in[95];
     assign  data_out[859] = data_in[1359];
     assign  data_out[860] = data_in[695];
     assign  data_out[861] = data_in[748];
     assign  data_out[862] = data_in[480];
     assign  data_out[863] = data_in[1254];
     assign  data_out[864] = data_in[975];
     assign  data_out[865] = data_in[1060];
     assign  data_out[866] = data_in[1602];
     assign  data_out[867] = data_in[1100];
     assign  data_out[868] = data_in[1653];
     assign  data_out[869] = data_in[1634];
     assign  data_out[870] = data_in[1296];
     assign  data_out[871] = data_in[1162];
     assign  data_out[872] = data_in[775];
     assign  data_out[873] = data_in[589];
     assign  data_out[874] = data_in[1647];
     assign  data_out[875] = data_in[1543];
     assign  data_out[876] = data_in[547];
     assign  data_out[877] = data_in[158];
     assign  data_out[878] = data_in[1370];
     assign  data_out[879] = data_in[1073];
     assign  data_out[880] = data_in[1404];
     assign  data_out[881] = data_in[504];
     assign  data_out[882] = data_in[1632];
     assign  data_out[883] = data_in[805];
     assign  data_out[884] = data_in[1226];
     assign  data_out[885] = data_in[552];
     assign  data_out[886] = data_in[1164];
     assign  data_out[887] = data_in[1603];
     assign  data_out[888] = data_in[191];
     assign  data_out[889] = data_in[939];
     assign  data_out[890] = data_in[599];
     assign  data_out[891] = data_in[1719];
     assign  data_out[892] = data_in[510];
     assign  data_out[893] = data_in[1561];
     assign  data_out[894] = data_in[536];
     assign  data_out[895] = data_in[1079];
     assign  data_out[896] = data_in[1537];
     assign  data_out[897] = data_in[906];
     assign  data_out[898] = data_in[1167];
     assign  data_out[899] = data_in[913];
     assign  data_out[900] = data_in[242];
     assign  data_out[901] = data_in[40];
     assign  data_out[902] = data_in[41];
     assign  data_out[903] = data_in[278];
     assign  data_out[904] = data_in[988];
     assign  data_out[905] = data_in[1135];
     assign  data_out[906] = data_in[1015];
     assign  data_out[907] = data_in[553];
     assign  data_out[908] = data_in[1405];
     assign  data_out[909] = data_in[1685];
     assign  data_out[910] = data_in[1581];
     assign  data_out[911] = data_in[457];
     assign  data_out[912] = data_in[1498];
     assign  data_out[913] = data_in[224];
     assign  data_out[914] = data_in[983];
     assign  data_out[915] = data_in[1307];
     assign  data_out[916] = data_in[1055];
     assign  data_out[917] = data_in[865];
     assign  data_out[918] = data_in[1509];
     assign  data_out[919] = data_in[1610];
     assign  data_out[920] = data_in[1393];
     assign  data_out[921] = data_in[1364];
     assign  data_out[922] = data_in[440];
     assign  data_out[923] = data_in[707];
     assign  data_out[924] = data_in[693];
     assign  data_out[925] = data_in[422];
     assign  data_out[926] = data_in[347];
     assign  data_out[927] = data_in[933];
     assign  data_out[928] = data_in[696];
     assign  data_out[929] = data_in[282];
     assign  data_out[930] = data_in[634];
     assign  data_out[931] = data_in[360];
     assign  data_out[932] = data_in[176];
     assign  data_out[933] = data_in[584];
     assign  data_out[934] = data_in[1501];
     assign  data_out[935] = data_in[147];
     assign  data_out[936] = data_in[1620];
     assign  data_out[937] = data_in[1035];
     assign  data_out[938] = data_in[489];
     assign  data_out[939] = data_in[1286];
     assign  data_out[940] = data_in[1335];
     assign  data_out[941] = data_in[180];
     assign  data_out[942] = data_in[684];
     assign  data_out[943] = data_in[943];
     assign  data_out[944] = data_in[1501];
     assign  data_out[945] = data_in[934];
     assign  data_out[946] = data_in[391];
     assign  data_out[947] = data_in[1198];
     assign  data_out[948] = data_in[588];
     assign  data_out[949] = data_in[1539];
     assign  data_out[950] = data_in[609];
     assign  data_out[951] = data_in[643];
     assign  data_out[952] = data_in[634];
     assign  data_out[953] = data_in[1585];
     assign  data_out[954] = data_in[144];
     assign  data_out[955] = data_in[639];
     assign  data_out[956] = data_in[1636];
     assign  data_out[957] = data_in[46];
     assign  data_out[958] = data_in[846];
     assign  data_out[959] = data_in[168];
     assign  data_out[960] = data_in[820];
     assign  data_out[961] = data_in[1150];
     assign  data_out[962] = data_in[1459];
     assign  data_out[963] = data_in[691];
     assign  data_out[964] = data_in[1591];
     assign  data_out[965] = data_in[1564];
     assign  data_out[966] = data_in[848];
     assign  data_out[967] = data_in[135];
     assign  data_out[968] = data_in[1544];
     assign  data_out[969] = data_in[646];
     assign  data_out[970] = data_in[1160];
     assign  data_out[971] = data_in[902];
     assign  data_out[972] = data_in[648];
     assign  data_out[973] = data_in[327];
     assign  data_out[974] = data_in[612];
     assign  data_out[975] = data_in[616];
     assign  data_out[976] = data_in[679];
     assign  data_out[977] = data_in[89];
     assign  data_out[978] = data_in[1013];
     assign  data_out[979] = data_in[892];
     assign  data_out[980] = data_in[745];
     assign  data_out[981] = data_in[252];
     assign  data_out[982] = data_in[683];
     assign  data_out[983] = data_in[1119];
     assign  data_out[984] = data_in[1459];
     assign  data_out[985] = data_in[40];
     assign  data_out[986] = data_in[1366];
     assign  data_out[987] = data_in[432];
     assign  data_out[988] = data_in[112];
     assign  data_out[989] = data_in[173];
     assign  data_out[990] = data_in[1510];
     assign  data_out[991] = data_in[786];
     assign  data_out[992] = data_in[1527];
     assign  data_out[993] = data_in[1639];
     assign  data_out[994] = data_in[1047];
     assign  data_out[995] = data_in[1483];
     assign  data_out[996] = data_in[1003];
     assign  data_out[997] = data_in[35];
     assign  data_out[998] = data_in[434];
     assign  data_out[999] = data_in[530];
     assign  data_out[1000] = data_in[336];
     assign  data_out[1001] = data_in[1673];
     assign  data_out[1002] = data_in[68];
     assign  data_out[1003] = data_in[73];
     assign  data_out[1004] = data_in[1221];
     assign  data_out[1005] = data_in[384];
     assign  data_out[1006] = data_in[114];
     assign  data_out[1007] = data_in[208];
     assign  data_out[1008] = data_in[725];
     assign  data_out[1009] = data_in[1675];
     assign  data_out[1010] = data_in[1685];
     assign  data_out[1011] = data_in[855];
     assign  data_out[1012] = data_in[554];
     assign  data_out[1013] = data_in[350];
     assign  data_out[1014] = data_in[762];
     assign  data_out[1015] = data_in[1193];
     assign  data_out[1016] = data_in[1202];
     assign  data_out[1017] = data_in[1703];
     assign  data_out[1018] = data_in[1715];
     assign  data_out[1019] = data_in[782];
     assign  data_out[1020] = data_in[1374];
     assign  data_out[1021] = data_in[1032];
     assign  data_out[1022] = data_in[360];
     assign  data_out[1023] = data_in[520];
     assign  data_out[1024] = data_in[1404];
     assign  data_out[1025] = data_in[1230];
     assign  data_out[1026] = data_in[1393];
     assign  data_out[1027] = data_in[640];
     assign  data_out[1028] = data_in[1680];
     assign  data_out[1029] = data_in[451];
     assign  data_out[1030] = data_in[1155];
     assign  data_out[1031] = data_in[806];
     assign  data_out[1032] = data_in[0];
     assign  data_out[1033] = data_in[261];
     assign  data_out[1034] = data_in[572];
     assign  data_out[1035] = data_in[1251];
     assign  data_out[1036] = data_in[1312];
     assign  data_out[1037] = data_in[820];
     assign  data_out[1038] = data_in[1664];
     assign  data_out[1039] = data_in[1367];
     assign  data_out[1040] = data_in[581];
     assign  data_out[1041] = data_in[664];
     assign  data_out[1042] = data_in[650];
     assign  data_out[1043] = data_in[1611];
     assign  data_out[1044] = data_in[608];
     assign  data_out[1045] = data_in[483];
     assign  data_out[1046] = data_in[147];
     assign  data_out[1047] = data_in[1661];
     assign  data_out[1048] = data_in[1356];
     assign  data_out[1049] = data_in[802];
     assign  data_out[1050] = data_in[1661];
     assign  data_out[1051] = data_in[713];
     assign  data_out[1052] = data_in[144];
     assign  data_out[1053] = data_in[1610];
     assign  data_out[1054] = data_in[869];
     assign  data_out[1055] = data_in[1478];
     assign  data_out[1056] = data_in[1473];
     assign  data_out[1057] = data_in[749];
     assign  data_out[1058] = data_in[441];
     assign  data_out[1059] = data_in[1303];
     assign  data_out[1060] = data_in[1545];
     assign  data_out[1061] = data_in[840];
     assign  data_out[1062] = data_in[718];
     assign  data_out[1063] = data_in[1356];
     assign  data_out[1064] = data_in[1516];
     assign  data_out[1065] = data_in[817];
     assign  data_out[1066] = data_in[252];
     assign  data_out[1067] = data_in[29];
     assign  data_out[1068] = data_in[748];
     assign  data_out[1069] = data_in[867];
     assign  data_out[1070] = data_in[1095];
     assign  data_out[1071] = data_in[1477];
     assign  data_out[1072] = data_in[1618];
     assign  data_out[1073] = data_in[287];
     assign  data_out[1074] = data_in[740];
     assign  data_out[1075] = data_in[279];
     assign  data_out[1076] = data_in[1342];
     assign  data_out[1077] = data_in[1512];
     assign  data_out[1078] = data_in[139];
     assign  data_out[1079] = data_in[786];
     assign  data_out[1080] = data_in[658];
     assign  data_out[1081] = data_in[1554];
     assign  data_out[1082] = data_in[1078];
     assign  data_out[1083] = data_in[1031];
     assign  data_out[1084] = data_in[1349];
     assign  data_out[1085] = data_in[1378];
     assign  data_out[1086] = data_in[1595];
     assign  data_out[1087] = data_in[1503];
     assign  data_out[1088] = data_in[1727];
     assign  data_out[1089] = data_in[650];
     assign  data_out[1090] = data_in[728];
     assign  data_out[1091] = data_in[1481];
     assign  data_out[1092] = data_in[83];
     assign  data_out[1093] = data_in[1443];
     assign  data_out[1094] = data_in[559];
     assign  data_out[1095] = data_in[37];
     assign  data_out[1096] = data_in[1381];
     assign  data_out[1097] = data_in[457];
     assign  data_out[1098] = data_in[1279];
     assign  data_out[1099] = data_in[696];
     assign  data_out[1100] = data_in[918];
     assign  data_out[1101] = data_in[238];
     assign  data_out[1102] = data_in[1420];
     assign  data_out[1103] = data_in[567];
     assign  data_out[1104] = data_in[723];
     assign  data_out[1105] = data_in[1671];
     assign  data_out[1106] = data_in[736];
     assign  data_out[1107] = data_in[944];
     assign  data_out[1108] = data_in[1297];
     assign  data_out[1109] = data_in[1332];
     assign  data_out[1110] = data_in[580];
     assign  data_out[1111] = data_in[1201];
     assign  data_out[1112] = data_in[277];
     assign  data_out[1113] = data_in[887];
     assign  data_out[1114] = data_in[977];
     assign  data_out[1115] = data_in[866];
     assign  data_out[1116] = data_in[1115];
     assign  data_out[1117] = data_in[295];
     assign  data_out[1118] = data_in[1368];
     assign  data_out[1119] = data_in[1083];
     assign  data_out[1120] = data_in[1133];
     assign  data_out[1121] = data_in[1003];
     assign  data_out[1122] = data_in[737];
     assign  data_out[1123] = data_in[968];
     assign  data_out[1124] = data_in[77];
     assign  data_out[1125] = data_in[1261];
     assign  data_out[1126] = data_in[655];
     assign  data_out[1127] = data_in[807];
     assign  data_out[1128] = data_in[250];
     assign  data_out[1129] = data_in[1104];
     assign  data_out[1130] = data_in[45];
     assign  data_out[1131] = data_in[684];
     assign  data_out[1132] = data_in[1323];
     assign  data_out[1133] = data_in[864];
     assign  data_out[1134] = data_in[740];
     assign  data_out[1135] = data_in[1312];
     assign  data_out[1136] = data_in[671];
     assign  data_out[1137] = data_in[378];
     assign  data_out[1138] = data_in[556];
     assign  data_out[1139] = data_in[835];
     assign  data_out[1140] = data_in[581];
     assign  data_out[1141] = data_in[47];
     assign  data_out[1142] = data_in[1581];
     assign  data_out[1143] = data_in[1275];
     assign  data_out[1144] = data_in[355];
     assign  data_out[1145] = data_in[534];
     assign  data_out[1146] = data_in[45];
     assign  data_out[1147] = data_in[1132];
     assign  data_out[1148] = data_in[590];
     assign  data_out[1149] = data_in[533];
     assign  data_out[1150] = data_in[1016];
     assign  data_out[1151] = data_in[1623];
     assign  data_out[1152] = data_in[1090];
     assign  data_out[1153] = data_in[1505];
     assign  data_out[1154] = data_in[89];
     assign  data_out[1155] = data_in[1340];
     assign  data_out[1156] = data_in[690];
     assign  data_out[1157] = data_in[1506];
     assign  data_out[1158] = data_in[1253];
     assign  data_out[1159] = data_in[1628];
     assign  data_out[1160] = data_in[1208];
     assign  data_out[1161] = data_in[846];
     assign  data_out[1162] = data_in[990];
     assign  data_out[1163] = data_in[931];
     assign  data_out[1164] = data_in[1303];
     assign  data_out[1165] = data_in[1702];
     assign  data_out[1166] = data_in[882];
     assign  data_out[1167] = data_in[393];
     assign  data_out[1168] = data_in[1484];
     assign  data_out[1169] = data_in[236];
     assign  data_out[1170] = data_in[1248];
     assign  data_out[1171] = data_in[689];
     assign  data_out[1172] = data_in[869];
     assign  data_out[1173] = data_in[1708];
     assign  data_out[1174] = data_in[68];
     assign  data_out[1175] = data_in[295];
     assign  data_out[1176] = data_in[9];
     assign  data_out[1177] = data_in[122];
     assign  data_out[1178] = data_in[1559];
     assign  data_out[1179] = data_in[1069];
     assign  data_out[1180] = data_in[761];
     assign  data_out[1181] = data_in[1294];
     assign  data_out[1182] = data_in[1635];
     assign  data_out[1183] = data_in[265];
     assign  data_out[1184] = data_in[240];
     assign  data_out[1185] = data_in[1473];
     assign  data_out[1186] = data_in[1263];
     assign  data_out[1187] = data_in[767];
     assign  data_out[1188] = data_in[923];
     assign  data_out[1189] = data_in[424];
     assign  data_out[1190] = data_in[1140];
     assign  data_out[1191] = data_in[1382];
     assign  data_out[1192] = data_in[1130];
     assign  data_out[1193] = data_in[849];
     assign  data_out[1194] = data_in[1045];
     assign  data_out[1195] = data_in[704];
     assign  data_out[1196] = data_in[35];
     assign  data_out[1197] = data_in[472];
     assign  data_out[1198] = data_in[485];
     assign  data_out[1199] = data_in[593];
     assign  data_out[1200] = data_in[428];
     assign  data_out[1201] = data_in[1236];
     assign  data_out[1202] = data_in[1541];
     assign  data_out[1203] = data_in[1299];
     assign  data_out[1204] = data_in[217];
     assign  data_out[1205] = data_in[480];
     assign  data_out[1206] = data_in[148];
     assign  data_out[1207] = data_in[193];
     assign  data_out[1208] = data_in[783];
     assign  data_out[1209] = data_in[630];
     assign  data_out[1210] = data_in[1292];
     assign  data_out[1211] = data_in[1697];
     assign  data_out[1212] = data_in[723];
     assign  data_out[1213] = data_in[538];
     assign  data_out[1214] = data_in[1137];
     assign  data_out[1215] = data_in[249];
     assign  data_out[1216] = data_in[1385];
     assign  data_out[1217] = data_in[1573];
     assign  data_out[1218] = data_in[964];
     assign  data_out[1219] = data_in[935];
     assign  data_out[1220] = data_in[1344];
     assign  data_out[1221] = data_in[198];
     assign  data_out[1222] = data_in[1104];
     assign  data_out[1223] = data_in[1597];
     assign  data_out[1224] = data_in[1051];
     assign  data_out[1225] = data_in[175];
     assign  data_out[1226] = data_in[5];
     assign  data_out[1227] = data_in[1052];
     assign  data_out[1228] = data_in[1716];
     assign  data_out[1229] = data_in[559];
     assign  data_out[1230] = data_in[188];
     assign  data_out[1231] = data_in[429];
     assign  data_out[1232] = data_in[655];
     assign  data_out[1233] = data_in[1264];
     assign  data_out[1234] = data_in[1296];
     assign  data_out[1235] = data_in[54];
     assign  data_out[1236] = data_in[1704];
     assign  data_out[1237] = data_in[1385];
     assign  data_out[1238] = data_in[1017];
     assign  data_out[1239] = data_in[365];
     assign  data_out[1240] = data_in[1471];
     assign  data_out[1241] = data_in[928];
     assign  data_out[1242] = data_in[1332];
     assign  data_out[1243] = data_in[637];
     assign  data_out[1244] = data_in[1138];
     assign  data_out[1245] = data_in[169];
     assign  data_out[1246] = data_in[1160];
     assign  data_out[1247] = data_in[552];
     assign  data_out[1248] = data_in[1118];
     assign  data_out[1249] = data_in[366];
     assign  data_out[1250] = data_in[484];
     assign  data_out[1251] = data_in[122];
     assign  data_out[1252] = data_in[631];
     assign  data_out[1253] = data_in[46];
     assign  data_out[1254] = data_in[475];
     assign  data_out[1255] = data_in[1263];
     assign  data_out[1256] = data_in[976];
     assign  data_out[1257] = data_in[961];
     assign  data_out[1258] = data_in[527];
     assign  data_out[1259] = data_in[1349];
     assign  data_out[1260] = data_in[18];
     assign  data_out[1261] = data_in[653];
     assign  data_out[1262] = data_in[899];
     assign  data_out[1263] = data_in[1065];
     assign  data_out[1264] = data_in[837];
     assign  data_out[1265] = data_in[1285];
     assign  data_out[1266] = data_in[1511];
     assign  data_out[1267] = data_in[1310];
     assign  data_out[1268] = data_in[1335];
     assign  data_out[1269] = data_in[1290];
     assign  data_out[1270] = data_in[408];
     assign  data_out[1271] = data_in[1122];
     assign  data_out[1272] = data_in[1566];
     assign  data_out[1273] = data_in[1238];
     assign  data_out[1274] = data_in[1447];
     assign  data_out[1275] = data_in[745];
     assign  data_out[1276] = data_in[778];
     assign  data_out[1277] = data_in[845];
     assign  data_out[1278] = data_in[154];
     assign  data_out[1279] = data_in[1068];
     assign  data_out[1280] = data_in[188];
     assign  data_out[1281] = data_in[1220];
     assign  data_out[1282] = data_in[522];
     assign  data_out[1283] = data_in[121];
     assign  data_out[1284] = data_in[754];
     assign  data_out[1285] = data_in[1397];
     assign  data_out[1286] = data_in[577];
     assign  data_out[1287] = data_in[286];
     assign  data_out[1288] = data_in[1614];
     assign  data_out[1289] = data_in[1512];
     assign  data_out[1290] = data_in[1216];
     assign  data_out[1291] = data_in[1024];
     assign  data_out[1292] = data_in[541];
     assign  data_out[1293] = data_in[1658];
     assign  data_out[1294] = data_in[340];
     assign  data_out[1295] = data_in[1125];
     assign  data_out[1296] = data_in[346];
     assign  data_out[1297] = data_in[155];
     assign  data_out[1298] = data_in[859];
     assign  data_out[1299] = data_in[837];
     assign  data_out[1300] = data_in[135];
     assign  data_out[1301] = data_in[1002];
     assign  data_out[1302] = data_in[1513];
     assign  data_out[1303] = data_in[239];
     assign  data_out[1304] = data_in[1265];
     assign  data_out[1305] = data_in[1404];
     assign  data_out[1306] = data_in[811];
     assign  data_out[1307] = data_in[1476];
     assign  data_out[1308] = data_in[1709];
     assign  data_out[1309] = data_in[257];
     assign  data_out[1310] = data_in[297];
     assign  data_out[1311] = data_in[882];
     assign  data_out[1312] = data_in[46];
     assign  data_out[1313] = data_in[211];
     assign  data_out[1314] = data_in[1183];
     assign  data_out[1315] = data_in[1048];
     assign  data_out[1316] = data_in[67];
     assign  data_out[1317] = data_in[983];
     assign  data_out[1318] = data_in[1282];
     assign  data_out[1319] = data_in[1222];
     assign  data_out[1320] = data_in[922];
     assign  data_out[1321] = data_in[1483];
     assign  data_out[1322] = data_in[87];
     assign  data_out[1323] = data_in[1286];
     assign  data_out[1324] = data_in[87];
     assign  data_out[1325] = data_in[1506];
     assign  data_out[1326] = data_in[1688];
     assign  data_out[1327] = data_in[153];
     assign  data_out[1328] = data_in[984];
     assign  data_out[1329] = data_in[1540];
     assign  data_out[1330] = data_in[875];
     assign  data_out[1331] = data_in[1371];
     assign  data_out[1332] = data_in[697];
     assign  data_out[1333] = data_in[89];
     assign  data_out[1334] = data_in[879];
     assign  data_out[1335] = data_in[1593];
     assign  data_out[1336] = data_in[1466];
     assign  data_out[1337] = data_in[891];
     assign  data_out[1338] = data_in[1459];
     assign  data_out[1339] = data_in[613];
     assign  data_out[1340] = data_in[651];
     assign  data_out[1341] = data_in[38];
     assign  data_out[1342] = data_in[580];
     assign  data_out[1343] = data_in[1723];
     assign  data_out[1344] = data_in[1118];
     assign  data_out[1345] = data_in[1678];
     assign  data_out[1346] = data_in[251];
     assign  data_out[1347] = data_in[1346];
     assign  data_out[1348] = data_in[217];
     assign  data_out[1349] = data_in[1205];
     assign  data_out[1350] = data_in[998];
     assign  data_out[1351] = data_in[629];
     assign  data_out[1352] = data_in[1013];
     assign  data_out[1353] = data_in[150];
     assign  data_out[1354] = data_in[1469];
     assign  data_out[1355] = data_in[1672];
     assign  data_out[1356] = data_in[480];
     assign  data_out[1357] = data_in[345];
     assign  data_out[1358] = data_in[1478];
     assign  data_out[1359] = data_in[337];
     assign  data_out[1360] = data_in[72];
     assign  data_out[1361] = data_in[84];
     assign  data_out[1362] = data_in[775];
     assign  data_out[1363] = data_in[518];
     assign  data_out[1364] = data_in[267];
     assign  data_out[1365] = data_in[332];
     assign  data_out[1366] = data_in[508];
     assign  data_out[1367] = data_in[1338];
     assign  data_out[1368] = data_in[313];
     assign  data_out[1369] = data_in[514];
     assign  data_out[1370] = data_in[1376];
     assign  data_out[1371] = data_in[1175];
     assign  data_out[1372] = data_in[1073];
     assign  data_out[1373] = data_in[578];
     assign  data_out[1374] = data_in[265];
     assign  data_out[1375] = data_in[1056];
     assign  data_out[1376] = data_in[1076];
     assign  data_out[1377] = data_in[943];
     assign  data_out[1378] = data_in[98];
     assign  data_out[1379] = data_in[1240];
     assign  data_out[1380] = data_in[963];
     assign  data_out[1381] = data_in[1495];
     assign  data_out[1382] = data_in[135];
     assign  data_out[1383] = data_in[1169];
     assign  data_out[1384] = data_in[1244];
     assign  data_out[1385] = data_in[1595];
     assign  data_out[1386] = data_in[458];
     assign  data_out[1387] = data_in[45];
     assign  data_out[1388] = data_in[1651];
     assign  data_out[1389] = data_in[536];
     assign  data_out[1390] = data_in[1696];
     assign  data_out[1391] = data_in[1329];
     assign  data_out[1392] = data_in[817];
     assign  data_out[1393] = data_in[425];
     assign  data_out[1394] = data_in[906];
     assign  data_out[1395] = data_in[1120];
     assign  data_out[1396] = data_in[1114];
     assign  data_out[1397] = data_in[541];
     assign  data_out[1398] = data_in[944];
     assign  data_out[1399] = data_in[4];
     assign  data_out[1400] = data_in[109];
     assign  data_out[1401] = data_in[712];
     assign  data_out[1402] = data_in[1411];
     assign  data_out[1403] = data_in[1050];
     assign  data_out[1404] = data_in[1100];
     assign  data_out[1405] = data_in[1024];
     assign  data_out[1406] = data_in[610];
     assign  data_out[1407] = data_in[718];
     assign  data_out[1408] = data_in[22];
     assign  data_out[1409] = data_in[1588];
     assign  data_out[1410] = data_in[775];
     assign  data_out[1411] = data_in[1009];
     assign  data_out[1412] = data_in[170];
     assign  data_out[1413] = data_in[43];
     assign  data_out[1414] = data_in[1100];
     assign  data_out[1415] = data_in[1238];
     assign  data_out[1416] = data_in[1679];
     assign  data_out[1417] = data_in[884];
     assign  data_out[1418] = data_in[198];
     assign  data_out[1419] = data_in[1233];
     assign  data_out[1420] = data_in[1644];
     assign  data_out[1421] = data_in[1470];
     assign  data_out[1422] = data_in[1147];
     assign  data_out[1423] = data_in[243];
     assign  data_out[1424] = data_in[216];
     assign  data_out[1425] = data_in[1636];
     assign  data_out[1426] = data_in[1022];
     assign  data_out[1427] = data_in[894];
     assign  data_out[1428] = data_in[161];
     assign  data_out[1429] = data_in[13];
     assign  data_out[1430] = data_in[1272];
     assign  data_out[1431] = data_in[764];
     assign  data_out[1432] = data_in[401];
     assign  data_out[1433] = data_in[1543];
     assign  data_out[1434] = data_in[89];
     assign  data_out[1435] = data_in[1639];
     assign  data_out[1436] = data_in[422];
     assign  data_out[1437] = data_in[1011];
     assign  data_out[1438] = data_in[1417];
     assign  data_out[1439] = data_in[10];
     assign  data_out[1440] = data_in[487];
     assign  data_out[1441] = data_in[1635];
     assign  data_out[1442] = data_in[12];
     assign  data_out[1443] = data_in[985];
     assign  data_out[1444] = data_in[730];
     assign  data_out[1445] = data_in[709];
     assign  data_out[1446] = data_in[1386];
     assign  data_out[1447] = data_in[148];
     assign  data_out[1448] = data_in[1351];
     assign  data_out[1449] = data_in[1342];
     assign  data_out[1450] = data_in[1509];
     assign  data_out[1451] = data_in[1478];
     assign  data_out[1452] = data_in[68];
     assign  data_out[1453] = data_in[1297];
     assign  data_out[1454] = data_in[629];
     assign  data_out[1455] = data_in[292];
     assign  data_out[1456] = data_in[1151];
     assign  data_out[1457] = data_in[685];
     assign  data_out[1458] = data_in[283];
     assign  data_out[1459] = data_in[1061];
     assign  data_out[1460] = data_in[1079];
     assign  data_out[1461] = data_in[259];
     assign  data_out[1462] = data_in[848];
     assign  data_out[1463] = data_in[799];
     assign  data_out[1464] = data_in[1439];
     assign  data_out[1465] = data_in[961];
     assign  data_out[1466] = data_in[526];
     assign  data_out[1467] = data_in[938];
     assign  data_out[1468] = data_in[294];
     assign  data_out[1469] = data_in[660];
     assign  data_out[1470] = data_in[1030];
     assign  data_out[1471] = data_in[878];
     assign  data_out[1472] = data_in[520];
     assign  data_out[1473] = data_in[454];
     assign  data_out[1474] = data_in[127];
     assign  data_out[1475] = data_in[1555];
     assign  data_out[1476] = data_in[184];
     assign  data_out[1477] = data_in[926];
     assign  data_out[1478] = data_in[483];
     assign  data_out[1479] = data_in[1589];
     assign  data_out[1480] = data_in[1726];
     assign  data_out[1481] = data_in[733];
     assign  data_out[1482] = data_in[1162];
     assign  data_out[1483] = data_in[532];
     assign  data_out[1484] = data_in[1554];
     assign  data_out[1485] = data_in[379];
     assign  data_out[1486] = data_in[1213];
     assign  data_out[1487] = data_in[426];
     assign  data_out[1488] = data_in[295];
     assign  data_out[1489] = data_in[1074];
     assign  data_out[1490] = data_in[712];
     assign  data_out[1491] = data_in[1173];
     assign  data_out[1492] = data_in[468];
     assign  data_out[1493] = data_in[1547];
     assign  data_out[1494] = data_in[1026];
     assign  data_out[1495] = data_in[1664];
     assign  data_out[1496] = data_in[721];
     assign  data_out[1497] = data_in[1725];
     assign  data_out[1498] = data_in[58];
     assign  data_out[1499] = data_in[455];
     assign  data_out[1500] = data_in[83];
     assign  data_out[1501] = data_in[576];
     assign  data_out[1502] = data_in[1517];
     assign  data_out[1503] = data_in[1001];
     assign  data_out[1504] = data_in[603];
     assign  data_out[1505] = data_in[494];
     assign  data_out[1506] = data_in[1118];
     assign  data_out[1507] = data_in[1433];
     assign  data_out[1508] = data_in[1100];
     assign  data_out[1509] = data_in[342];
     assign  data_out[1510] = data_in[1608];
     assign  data_out[1511] = data_in[1525];
     assign  data_out[1512] = data_in[1515];
     assign  data_out[1513] = data_in[1630];
     assign  data_out[1514] = data_in[516];
     assign  data_out[1515] = data_in[1659];
     assign  data_out[1516] = data_in[203];
     assign  data_out[1517] = data_in[1295];
     assign  data_out[1518] = data_in[785];
     assign  data_out[1519] = data_in[513];
     assign  data_out[1520] = data_in[207];
     assign  data_out[1521] = data_in[743];
     assign  data_out[1522] = data_in[280];
     assign  data_out[1523] = data_in[832];
     assign  data_out[1524] = data_in[1675];
     assign  data_out[1525] = data_in[1176];
     assign  data_out[1526] = data_in[1702];
     assign  data_out[1527] = data_in[648];
     assign  data_out[1528] = data_in[1627];
     assign  data_out[1529] = data_in[1034];
     assign  data_out[1530] = data_in[614];
     assign  data_out[1531] = data_in[24];
     assign  data_out[1532] = data_in[720];
     assign  data_out[1533] = data_in[125];
     assign  data_out[1534] = data_in[35];
     assign  data_out[1535] = data_in[707];
     assign  data_out[1536] = data_in[187];
     assign  data_out[1537] = data_in[370];
     assign  data_out[1538] = data_in[659];
     assign  data_out[1539] = data_in[1113];
     assign  data_out[1540] = data_in[695];
     assign  data_out[1541] = data_in[819];
     assign  data_out[1542] = data_in[1336];
     assign  data_out[1543] = data_in[296];
     assign  data_out[1544] = data_in[131];
     assign  data_out[1545] = data_in[1039];
     assign  data_out[1546] = data_in[339];
     assign  data_out[1547] = data_in[1261];
     assign  data_out[1548] = data_in[321];
     assign  data_out[1549] = data_in[194];
     assign  data_out[1550] = data_in[952];
     assign  data_out[1551] = data_in[1337];
     assign  data_out[1552] = data_in[691];
     assign  data_out[1553] = data_in[710];
     assign  data_out[1554] = data_in[1549];
     assign  data_out[1555] = data_in[1426];
     assign  data_out[1556] = data_in[975];
     assign  data_out[1557] = data_in[387];
     assign  data_out[1558] = data_in[1313];
     assign  data_out[1559] = data_in[1141];
     assign  data_out[1560] = data_in[1330];
     assign  data_out[1561] = data_in[889];
     assign  data_out[1562] = data_in[71];
     assign  data_out[1563] = data_in[1259];
     assign  data_out[1564] = data_in[1247];
     assign  data_out[1565] = data_in[883];
     assign  data_out[1566] = data_in[919];
     assign  data_out[1567] = data_in[1239];
     assign  data_out[1568] = data_in[1157];
     assign  data_out[1569] = data_in[47];
     assign  data_out[1570] = data_in[1016];
     assign  data_out[1571] = data_in[1143];
     assign  data_out[1572] = data_in[1212];
     assign  data_out[1573] = data_in[1248];
     assign  data_out[1574] = data_in[1696];
     assign  data_out[1575] = data_in[887];
     assign  data_out[1576] = data_in[1146];
     assign  data_out[1577] = data_in[776];
     assign  data_out[1578] = data_in[803];
     assign  data_out[1579] = data_in[983];
     assign  data_out[1580] = data_in[869];
     assign  data_out[1581] = data_in[627];
     assign  data_out[1582] = data_in[141];
     assign  data_out[1583] = data_in[1145];
     assign  data_out[1584] = data_in[526];
     assign  data_out[1585] = data_in[1614];
     assign  data_out[1586] = data_in[1304];
     assign  data_out[1587] = data_in[937];
     assign  data_out[1588] = data_in[1392];
     assign  data_out[1589] = data_in[907];
     assign  data_out[1590] = data_in[296];
     assign  data_out[1591] = data_in[539];
     assign  data_out[1592] = data_in[1161];
     assign  data_out[1593] = data_in[1190];
     assign  data_out[1594] = data_in[896];
     assign  data_out[1595] = data_in[646];
     assign  data_out[1596] = data_in[544];
     assign  data_out[1597] = data_in[1459];
     assign  data_out[1598] = data_in[138];
     assign  data_out[1599] = data_in[1303];
     assign  data_out[1600] = data_in[915];
     assign  data_out[1601] = data_in[841];
     assign  data_out[1602] = data_in[404];
     assign  data_out[1603] = data_in[400];
     assign  data_out[1604] = data_in[1274];
     assign  data_out[1605] = data_in[1008];
     assign  data_out[1606] = data_in[1530];
     assign  data_out[1607] = data_in[291];
     assign  data_out[1608] = data_in[193];
     assign  data_out[1609] = data_in[548];
     assign  data_out[1610] = data_in[1486];
     assign  data_out[1611] = data_in[791];
     assign  data_out[1612] = data_in[647];
     assign  data_out[1613] = data_in[1445];
     assign  data_out[1614] = data_in[502];
     assign  data_out[1615] = data_in[831];
     assign  data_out[1616] = data_in[921];
     assign  data_out[1617] = data_in[263];
     assign  data_out[1618] = data_in[918];
     assign  data_out[1619] = data_in[859];
     assign  data_out[1620] = data_in[605];
     assign  data_out[1621] = data_in[1493];
     assign  data_out[1622] = data_in[1084];
     assign  data_out[1623] = data_in[614];
     assign  data_out[1624] = data_in[1423];
     assign  data_out[1625] = data_in[1455];
     assign  data_out[1626] = data_in[1508];
     assign  data_out[1627] = data_in[1637];
     assign  data_out[1628] = data_in[786];
     assign  data_out[1629] = data_in[948];
     assign  data_out[1630] = data_in[841];
     assign  data_out[1631] = data_in[524];
     assign  data_out[1632] = data_in[1020];
     assign  data_out[1633] = data_in[232];
     assign  data_out[1634] = data_in[1628];
     assign  data_out[1635] = data_in[1267];
     assign  data_out[1636] = data_in[1069];
     assign  data_out[1637] = data_in[1689];
     assign  data_out[1638] = data_in[1680];
     assign  data_out[1639] = data_in[1601];
     assign  data_out[1640] = data_in[518];
     assign  data_out[1641] = data_in[1415];
     assign  data_out[1642] = data_in[1374];
     assign  data_out[1643] = data_in[708];
     assign  data_out[1644] = data_in[19];
     assign  data_out[1645] = data_in[256];
     assign  data_out[1646] = data_in[998];
     assign  data_out[1647] = data_in[478];
     assign  data_out[1648] = data_in[330];
     assign  data_out[1649] = data_in[1724];
     assign  data_out[1650] = data_in[1171];
     assign  data_out[1651] = data_in[1013];
     assign  data_out[1652] = data_in[1315];
     assign  data_out[1653] = data_in[1386];
     assign  data_out[1654] = data_in[1197];
     assign  data_out[1655] = data_in[597];
     assign  data_out[1656] = data_in[1395];
     assign  data_out[1657] = data_in[826];
     assign  data_out[1658] = data_in[1457];
     assign  data_out[1659] = data_in[824];
     assign  data_out[1660] = data_in[527];
     assign  data_out[1661] = data_in[658];
     assign  data_out[1662] = data_in[1263];
     assign  data_out[1663] = data_in[1171];
     assign  data_out[1664] = data_in[278];
     assign  data_out[1665] = data_in[507];
     assign  data_out[1666] = data_in[1714];
     assign  data_out[1667] = data_in[1000];
     assign  data_out[1668] = data_in[627];
     assign  data_out[1669] = data_in[187];
     assign  data_out[1670] = data_in[1528];
     assign  data_out[1671] = data_in[188];
     assign  data_out[1672] = data_in[888];
     assign  data_out[1673] = data_in[601];
     assign  data_out[1674] = data_in[584];
     assign  data_out[1675] = data_in[812];
     assign  data_out[1676] = data_in[917];
     assign  data_out[1677] = data_in[341];
     assign  data_out[1678] = data_in[864];
     assign  data_out[1679] = data_in[1087];
     assign  data_out[1680] = data_in[1366];
     assign  data_out[1681] = data_in[319];
     assign  data_out[1682] = data_in[523];
     assign  data_out[1683] = data_in[1272];
     assign  data_out[1684] = data_in[875];
     assign  data_out[1685] = data_in[316];
     assign  data_out[1686] = data_in[153];
     assign  data_out[1687] = data_in[640];
     assign  data_out[1688] = data_in[1057];
     assign  data_out[1689] = data_in[1523];
     assign  data_out[1690] = data_in[1430];
     assign  data_out[1691] = data_in[40];
     assign  data_out[1692] = data_in[1619];
     assign  data_out[1693] = data_in[655];
     assign  data_out[1694] = data_in[1638];
     assign  data_out[1695] = data_in[1249];
     assign  data_out[1696] = data_in[1653];
     assign  data_out[1697] = data_in[120];
     assign  data_out[1698] = data_in[552];
     assign  data_out[1699] = data_in[363];
     assign  data_out[1700] = data_in[1540];
     assign  data_out[1701] = data_in[792];
     assign  data_out[1702] = data_in[726];
     assign  data_out[1703] = data_in[982];
     assign  data_out[1704] = data_in[769];
     assign  data_out[1705] = data_in[137];
     assign  data_out[1706] = data_in[370];
     assign  data_out[1707] = data_in[1231];
     assign  data_out[1708] = data_in[1652];
     assign  data_out[1709] = data_in[280];
     assign  data_out[1710] = data_in[1333];
     assign  data_out[1711] = data_in[1120];
     assign  data_out[1712] = data_in[431];
     assign  data_out[1713] = data_in[360];
     assign  data_out[1714] = data_in[291];
     assign  data_out[1715] = data_in[1564];
     assign  data_out[1716] = data_in[1662];
     assign  data_out[1717] = data_in[226];
     assign  data_out[1718] = data_in[1195];
     assign  data_out[1719] = data_in[84];
     assign  data_out[1720] = data_in[1091];
     assign  data_out[1721] = data_in[202];
     assign  data_out[1722] = data_in[1517];
     assign  data_out[1723] = data_in[1169];
     assign  data_out[1724] = data_in[565];
     assign  data_out[1725] = data_in[1491];
     assign  data_out[1726] = data_in[740];
     assign  data_out[1727] = data_in[1407];
     assign  data_out[1728] = data_in[169];
     assign  data_out[1729] = data_in[600];
     assign  data_out[1730] = data_in[893];
     assign  data_out[1731] = data_in[176];
     assign  data_out[1732] = data_in[55];
     assign  data_out[1733] = data_in[1370];
     assign  data_out[1734] = data_in[927];
     assign  data_out[1735] = data_in[1191];
     assign  data_out[1736] = data_in[329];
     assign  data_out[1737] = data_in[1674];
     assign  data_out[1738] = data_in[1389];
     assign  data_out[1739] = data_in[423];
     assign  data_out[1740] = data_in[377];
     assign  data_out[1741] = data_in[868];
     assign  data_out[1742] = data_in[450];
     assign  data_out[1743] = data_in[1687];
     assign  data_out[1744] = data_in[1543];
     assign  data_out[1745] = data_in[596];
     assign  data_out[1746] = data_in[1204];
     assign  data_out[1747] = data_in[143];
     assign  data_out[1748] = data_in[707];
     assign  data_out[1749] = data_in[89];
     assign  data_out[1750] = data_in[926];
     assign  data_out[1751] = data_in[913];
     assign  data_out[1752] = data_in[1153];
     assign  data_out[1753] = data_in[56];
     assign  data_out[1754] = data_in[1217];
     assign  data_out[1755] = data_in[967];
     assign  data_out[1756] = data_in[618];
     assign  data_out[1757] = data_in[748];
     assign  data_out[1758] = data_in[1071];
     assign  data_out[1759] = data_in[1487];
     assign  data_out[1760] = data_in[196];
     assign  data_out[1761] = data_in[1374];
     assign  data_out[1762] = data_in[1438];
     assign  data_out[1763] = data_in[1311];
     assign  data_out[1764] = data_in[898];
     assign  data_out[1765] = data_in[273];
     assign  data_out[1766] = data_in[594];
     assign  data_out[1767] = data_in[668];
     assign  data_out[1768] = data_in[442];
     assign  data_out[1769] = data_in[1303];
     assign  data_out[1770] = data_in[251];
     assign  data_out[1771] = data_in[353];
     assign  data_out[1772] = data_in[264];
     assign  data_out[1773] = data_in[1660];
     assign  data_out[1774] = data_in[1716];
     assign  data_out[1775] = data_in[1360];
     assign  data_out[1776] = data_in[780];
     assign  data_out[1777] = data_in[1129];
     assign  data_out[1778] = data_in[1664];
     assign  data_out[1779] = data_in[501];
     assign  data_out[1780] = data_in[61];
     assign  data_out[1781] = data_in[1090];
     assign  data_out[1782] = data_in[1401];
     assign  data_out[1783] = data_in[851];
     assign  data_out[1784] = data_in[1601];
     assign  data_out[1785] = data_in[441];
     assign  data_out[1786] = data_in[1161];
     assign  data_out[1787] = data_in[1427];
     assign  data_out[1788] = data_in[1415];
     assign  data_out[1789] = data_in[1679];
     assign  data_out[1790] = data_in[219];
     assign  data_out[1791] = data_in[517];
     assign  data_out[1792] = data_in[1618];
     assign  data_out[1793] = data_in[1488];
     assign  data_out[1794] = data_in[294];
     assign  data_out[1795] = data_in[1238];
     assign  data_out[1796] = data_in[1721];
     assign  data_out[1797] = data_in[1523];
     assign  data_out[1798] = data_in[190];
     assign  data_out[1799] = data_in[185];
     assign  data_out[1800] = data_in[951];
     assign  data_out[1801] = data_in[1649];
     assign  data_out[1802] = data_in[1610];
     assign  data_out[1803] = data_in[1315];
     assign  data_out[1804] = data_in[868];
     assign  data_out[1805] = data_in[965];
     assign  data_out[1806] = data_in[261];
     assign  data_out[1807] = data_in[1355];
     assign  data_out[1808] = data_in[107];
     assign  data_out[1809] = data_in[1679];
     assign  data_out[1810] = data_in[1210];
     assign  data_out[1811] = data_in[1000];
     assign  data_out[1812] = data_in[1616];
     assign  data_out[1813] = data_in[1447];
     assign  data_out[1814] = data_in[1490];
     assign  data_out[1815] = data_in[262];
     assign  data_out[1816] = data_in[40];
     assign  data_out[1817] = data_in[338];
     assign  data_out[1818] = data_in[1386];
     assign  data_out[1819] = data_in[1141];
     assign  data_out[1820] = data_in[701];
     assign  data_out[1821] = data_in[1110];
     assign  data_out[1822] = data_in[1224];
     assign  data_out[1823] = data_in[174];
     assign  data_out[1824] = data_in[1568];
     assign  data_out[1825] = data_in[1339];
     assign  data_out[1826] = data_in[157];
     assign  data_out[1827] = data_in[940];
     assign  data_out[1828] = data_in[13];
     assign  data_out[1829] = data_in[987];
     assign  data_out[1830] = data_in[449];
     assign  data_out[1831] = data_in[1432];
     assign  data_out[1832] = data_in[676];
     assign  data_out[1833] = data_in[1503];
     assign  data_out[1834] = data_in[886];
     assign  data_out[1835] = data_in[198];
     assign  data_out[1836] = data_in[1581];
     assign  data_out[1837] = data_in[1038];
     assign  data_out[1838] = data_in[126];
     assign  data_out[1839] = data_in[351];
     assign  data_out[1840] = data_in[461];
     assign  data_out[1841] = data_in[1591];
     assign  data_out[1842] = data_in[513];
     assign  data_out[1843] = data_in[55];
     assign  data_out[1844] = data_in[188];
     assign  data_out[1845] = data_in[1591];
     assign  data_out[1846] = data_in[333];
     assign  data_out[1847] = data_in[432];
     assign  data_out[1848] = data_in[1688];
     assign  data_out[1849] = data_in[75];
     assign  data_out[1850] = data_in[1336];
     assign  data_out[1851] = data_in[482];
     assign  data_out[1852] = data_in[1246];
     assign  data_out[1853] = data_in[1537];
     assign  data_out[1854] = data_in[486];
     assign  data_out[1855] = data_in[1324];
     assign  data_out[1856] = data_in[1334];
     assign  data_out[1857] = data_in[946];
     assign  data_out[1858] = data_in[1404];
     assign  data_out[1859] = data_in[1450];
     assign  data_out[1860] = data_in[12];
     assign  data_out[1861] = data_in[203];
     assign  data_out[1862] = data_in[644];
     assign  data_out[1863] = data_in[104];
     assign  data_out[1864] = data_in[866];
     assign  data_out[1865] = data_in[1004];
     assign  data_out[1866] = data_in[1547];
     assign  data_out[1867] = data_in[859];
     assign  data_out[1868] = data_in[1636];
     assign  data_out[1869] = data_in[1161];
     assign  data_out[1870] = data_in[437];
     assign  data_out[1871] = data_in[1402];
     assign  data_out[1872] = data_in[29];
     assign  data_out[1873] = data_in[1560];
     assign  data_out[1874] = data_in[1381];
     assign  data_out[1875] = data_in[1321];
     assign  data_out[1876] = data_in[799];
     assign  data_out[1877] = data_in[710];
     assign  data_out[1878] = data_in[795];
     assign  data_out[1879] = data_in[107];
     assign  data_out[1880] = data_in[368];
     assign  data_out[1881] = data_in[1333];
     assign  data_out[1882] = data_in[1589];
     assign  data_out[1883] = data_in[1605];
     assign  data_out[1884] = data_in[469];
     assign  data_out[1885] = data_in[759];
     assign  data_out[1886] = data_in[1586];
     assign  data_out[1887] = data_in[568];
     assign  data_out[1888] = data_in[1181];
     assign  data_out[1889] = data_in[1678];
     assign  data_out[1890] = data_in[359];
     assign  data_out[1891] = data_in[402];
     assign  data_out[1892] = data_in[614];
     assign  data_out[1893] = data_in[1195];
     assign  data_out[1894] = data_in[321];
     assign  data_out[1895] = data_in[1454];
     assign  data_out[1896] = data_in[16];
     assign  data_out[1897] = data_in[1644];
     assign  data_out[1898] = data_in[1279];
     assign  data_out[1899] = data_in[297];
     assign  data_out[1900] = data_in[100];
     assign  data_out[1901] = data_in[1104];
     assign  data_out[1902] = data_in[589];
     assign  data_out[1903] = data_in[1566];
     assign  data_out[1904] = data_in[1153];
     assign  data_out[1905] = data_in[171];
     assign  data_out[1906] = data_in[1568];
     assign  data_out[1907] = data_in[1592];
     assign  data_out[1908] = data_in[1398];
     assign  data_out[1909] = data_in[207];
     assign  data_out[1910] = data_in[829];
     assign  data_out[1911] = data_in[680];
     assign  data_out[1912] = data_in[975];
     assign  data_out[1913] = data_in[229];
     assign  data_out[1914] = data_in[399];
     assign  data_out[1915] = data_in[1536];
     assign  data_out[1916] = data_in[817];
     assign  data_out[1917] = data_in[515];
     assign  data_out[1918] = data_in[1464];
     assign  data_out[1919] = data_in[607];
     assign  data_out[1920] = data_in[347];
     assign  data_out[1921] = data_in[1070];
     assign  data_out[1922] = data_in[1393];
     assign  data_out[1923] = data_in[666];
     assign  data_out[1924] = data_in[548];
     assign  data_out[1925] = data_in[1289];
     assign  data_out[1926] = data_in[1023];
     assign  data_out[1927] = data_in[1287];
     assign  data_out[1928] = data_in[780];
     assign  data_out[1929] = data_in[1078];
     assign  data_out[1930] = data_in[635];
     assign  data_out[1931] = data_in[746];
     assign  data_out[1932] = data_in[1064];
     assign  data_out[1933] = data_in[1122];
     assign  data_out[1934] = data_in[251];
     assign  data_out[1935] = data_in[549];
     assign  data_out[1936] = data_in[1693];
     assign  data_out[1937] = data_in[821];
     assign  data_out[1938] = data_in[1693];
     assign  data_out[1939] = data_in[1176];
     assign  data_out[1940] = data_in[1499];
     assign  data_out[1941] = data_in[242];
     assign  data_out[1942] = data_in[384];
     assign  data_out[1943] = data_in[1005];
     assign  data_out[1944] = data_in[466];
     assign  data_out[1945] = data_in[1142];
     assign  data_out[1946] = data_in[613];
     assign  data_out[1947] = data_in[809];
     assign  data_out[1948] = data_in[1113];
     assign  data_out[1949] = data_in[1304];
     assign  data_out[1950] = data_in[784];
     assign  data_out[1951] = data_in[1606];
     assign  data_out[1952] = data_in[498];
     assign  data_out[1953] = data_in[1464];
     assign  data_out[1954] = data_in[1372];
     assign  data_out[1955] = data_in[1712];
     assign  data_out[1956] = data_in[113];
     assign  data_out[1957] = data_in[24];
     assign  data_out[1958] = data_in[1106];
     assign  data_out[1959] = data_in[1508];
     assign  data_out[1960] = data_in[1328];
     assign  data_out[1961] = data_in[42];
     assign  data_out[1962] = data_in[1299];
     assign  data_out[1963] = data_in[1043];
     assign  data_out[1964] = data_in[1547];
     assign  data_out[1965] = data_in[228];
     assign  data_out[1966] = data_in[1084];
     assign  data_out[1967] = data_in[701];
     assign  data_out[1968] = data_in[212];
     assign  data_out[1969] = data_in[1341];
     assign  data_out[1970] = data_in[52];
     assign  data_out[1971] = data_in[432];
     assign  data_out[1972] = data_in[454];
     assign  data_out[1973] = data_in[1463];
     assign  data_out[1974] = data_in[1407];
     assign  data_out[1975] = data_in[855];
     assign  data_out[1976] = data_in[1682];
     assign  data_out[1977] = data_in[1161];
     assign  data_out[1978] = data_in[1027];
     assign  data_out[1979] = data_in[15];
     assign  data_out[1980] = data_in[23];
     assign  data_out[1981] = data_in[654];
     assign  data_out[1982] = data_in[483];
     assign  data_out[1983] = data_in[1190];
     assign  data_out[1984] = data_in[549];
     assign  data_out[1985] = data_in[1365];
     assign  data_out[1986] = data_in[21];
     assign  data_out[1987] = data_in[1333];
     assign  data_out[1988] = data_in[1172];
     assign  data_out[1989] = data_in[882];
     assign  data_out[1990] = data_in[925];
     assign  data_out[1991] = data_in[1484];
     assign  data_out[1992] = data_in[534];
     assign  data_out[1993] = data_in[620];
     assign  data_out[1994] = data_in[904];
     assign  data_out[1995] = data_in[75];
     assign  data_out[1996] = data_in[129];
     assign  data_out[1997] = data_in[1378];
     assign  data_out[1998] = data_in[1569];
     assign  data_out[1999] = data_in[109];
     assign  data_out[2000] = data_in[1158];
     assign  data_out[2001] = data_in[912];
     assign  data_out[2002] = data_in[1259];
     assign  data_out[2003] = data_in[1502];
     assign  data_out[2004] = data_in[910];
     assign  data_out[2005] = data_in[1547];
     assign  data_out[2006] = data_in[934];
     assign  data_out[2007] = data_in[921];
     assign  data_out[2008] = data_in[1256];
     assign  data_out[2009] = data_in[455];
     assign  data_out[2010] = data_in[1569];
     assign  data_out[2011] = data_in[1525];
     assign  data_out[2012] = data_in[1232];
     assign  data_out[2013] = data_in[36];
     assign  data_out[2014] = data_in[37];
     assign  data_out[2015] = data_in[1359];
     assign  data_out[2016] = data_in[115];
     assign  data_out[2017] = data_in[631];
     assign  data_out[2018] = data_in[1659];
     assign  data_out[2019] = data_in[836];
     assign  data_out[2020] = data_in[243];
     assign  data_out[2021] = data_in[920];
     assign  data_out[2022] = data_in[1105];
     assign  data_out[2023] = data_in[1501];
     assign  data_out[2024] = data_in[1429];
     assign  data_out[2025] = data_in[1061];
     assign  data_out[2026] = data_in[1677];
     assign  data_out[2027] = data_in[241];
     assign  data_out[2028] = data_in[417];
     assign  data_out[2029] = data_in[1100];
     assign  data_out[2030] = data_in[453];
     assign  data_out[2031] = data_in[1230];
     assign  data_out[2032] = data_in[1043];
     assign  data_out[2033] = data_in[67];
     assign  data_out[2034] = data_in[695];
     assign  data_out[2035] = data_in[1397];
     assign  data_out[2036] = data_in[167];
     assign  data_out[2037] = data_in[383];
     assign  data_out[2038] = data_in[1451];
     assign  data_out[2039] = data_in[1083];
     assign  data_out[2040] = data_in[1705];
     assign  data_out[2041] = data_in[540];
     assign  data_out[2042] = data_in[1575];
     assign  data_out[2043] = data_in[852];
     assign  data_out[2044] = data_in[1352];
     assign  data_out[2045] = data_in[1405];
     assign  data_out[2046] = data_in[922];
     assign  data_out[2047] = data_in[1577];
     assign  data_out[2048] = data_in[1242];
     assign  data_out[2049] = data_in[470];
     assign  data_out[2050] = data_in[1368];
     assign  data_out[2051] = data_in[1579];
     assign  data_out[2052] = data_in[592];
     assign  data_out[2053] = data_in[1133];
     assign  data_out[2054] = data_in[813];
     assign  data_out[2055] = data_in[1035];
     assign  data_out[2056] = data_in[834];
     assign  data_out[2057] = data_in[967];
     assign  data_out[2058] = data_in[63];
     assign  data_out[2059] = data_in[537];
     assign  data_out[2060] = data_in[670];
     assign  data_out[2061] = data_in[1594];
     assign  data_out[2062] = data_in[211];
     assign  data_out[2063] = data_in[531];
     assign  data_out[2064] = data_in[535];
     assign  data_out[2065] = data_in[688];
     assign  data_out[2066] = data_in[56];
     assign  data_out[2067] = data_in[640];
     assign  data_out[2068] = data_in[548];
     assign  data_out[2069] = data_in[77];
     assign  data_out[2070] = data_in[532];
     assign  data_out[2071] = data_in[411];
     assign  data_out[2072] = data_in[1066];
     assign  data_out[2073] = data_in[829];
     assign  data_out[2074] = data_in[1516];
     assign  data_out[2075] = data_in[475];
     assign  data_out[2076] = data_in[289];
     assign  data_out[2077] = data_in[291];
     assign  data_out[2078] = data_in[1426];
     assign  data_out[2079] = data_in[494];
     assign  data_out[2080] = data_in[1493];
     assign  data_out[2081] = data_in[1709];
     assign  data_out[2082] = data_in[550];
     assign  data_out[2083] = data_in[1518];
     assign  data_out[2084] = data_in[141];
     assign  data_out[2085] = data_in[1279];
     assign  data_out[2086] = data_in[1213];
     assign  data_out[2087] = data_in[480];
     assign  data_out[2088] = data_in[1456];
     assign  data_out[2089] = data_in[1289];
     assign  data_out[2090] = data_in[554];
     assign  data_out[2091] = data_in[13];
     assign  data_out[2092] = data_in[711];
     assign  data_out[2093] = data_in[362];
     assign  data_out[2094] = data_in[130];
     assign  data_out[2095] = data_in[578];
     assign  data_out[2096] = data_in[1005];
     assign  data_out[2097] = data_in[823];
     assign  data_out[2098] = data_in[448];
     assign  data_out[2099] = data_in[1535];
     assign  data_out[2100] = data_in[758];
     assign  data_out[2101] = data_in[1491];
     assign  data_out[2102] = data_in[1206];
     assign  data_out[2103] = data_in[624];
     assign  data_out[2104] = data_in[1533];
     assign  data_out[2105] = data_in[355];
     assign  data_out[2106] = data_in[1265];
     assign  data_out[2107] = data_in[1200];
     assign  data_out[2108] = data_in[1243];
     assign  data_out[2109] = data_in[1352];
     assign  data_out[2110] = data_in[110];
     assign  data_out[2111] = data_in[1138];
     assign  data_out[2112] = data_in[863];
     assign  data_out[2113] = data_in[1344];
     assign  data_out[2114] = data_in[11];
     assign  data_out[2115] = data_in[393];
     assign  data_out[2116] = data_in[106];
     assign  data_out[2117] = data_in[1599];
     assign  data_out[2118] = data_in[284];
     assign  data_out[2119] = data_in[1147];
     assign  data_out[2120] = data_in[1520];
     assign  data_out[2121] = data_in[870];
     assign  data_out[2122] = data_in[138];
     assign  data_out[2123] = data_in[1230];
     assign  data_out[2124] = data_in[205];
     assign  data_out[2125] = data_in[573];
     assign  data_out[2126] = data_in[1498];
     assign  data_out[2127] = data_in[1400];
     assign  data_out[2128] = data_in[1069];
     assign  data_out[2129] = data_in[1597];
     assign  data_out[2130] = data_in[651];
     assign  data_out[2131] = data_in[1254];
     assign  data_out[2132] = data_in[1065];
     assign  data_out[2133] = data_in[791];
     assign  data_out[2134] = data_in[1586];
     assign  data_out[2135] = data_in[898];
     assign  data_out[2136] = data_in[819];
     assign  data_out[2137] = data_in[1228];
     assign  data_out[2138] = data_in[106];
     assign  data_out[2139] = data_in[431];
     assign  data_out[2140] = data_in[340];
     assign  data_out[2141] = data_in[1089];
     assign  data_out[2142] = data_in[987];
     assign  data_out[2143] = data_in[540];
     assign  data_out[2144] = data_in[47];
     assign  data_out[2145] = data_in[1177];
     assign  data_out[2146] = data_in[1692];
     assign  data_out[2147] = data_in[1452];
     assign  data_out[2148] = data_in[1540];
     assign  data_out[2149] = data_in[1093];
     assign  data_out[2150] = data_in[1460];
     assign  data_out[2151] = data_in[81];
     assign  data_out[2152] = data_in[1682];
     assign  data_out[2153] = data_in[1633];
     assign  data_out[2154] = data_in[391];
     assign  data_out[2155] = data_in[1618];
     assign  data_out[2156] = data_in[380];
     assign  data_out[2157] = data_in[703];
     assign  data_out[2158] = data_in[686];
     assign  data_out[2159] = data_in[489];
     assign  data_out[2160] = data_in[46];
     assign  data_out[2161] = data_in[303];
     assign  data_out[2162] = data_in[583];
     assign  data_out[2163] = data_in[483];
     assign  data_out[2164] = data_in[1580];
     assign  data_out[2165] = data_in[1538];
     assign  data_out[2166] = data_in[55];
     assign  data_out[2167] = data_in[1331];
     assign  data_out[2168] = data_in[793];
     assign  data_out[2169] = data_in[1727];
     assign  data_out[2170] = data_in[181];
     assign  data_out[2171] = data_in[807];
     assign  data_out[2172] = data_in[455];
     assign  data_out[2173] = data_in[1675];
     assign  data_out[2174] = data_in[1427];
     assign  data_out[2175] = data_in[106];
     assign  data_out[2176] = data_in[443];
     assign  data_out[2177] = data_in[901];
     assign  data_out[2178] = data_in[29];
     assign  data_out[2179] = data_in[1087];
     assign  data_out[2180] = data_in[150];
     assign  data_out[2181] = data_in[974];
     assign  data_out[2182] = data_in[1530];
     assign  data_out[2183] = data_in[430];
     assign  data_out[2184] = data_in[1571];
     assign  data_out[2185] = data_in[1667];
     assign  data_out[2186] = data_in[568];
     assign  data_out[2187] = data_in[390];
     assign  data_out[2188] = data_in[575];
     assign  data_out[2189] = data_in[1437];
     assign  data_out[2190] = data_in[1249];
     assign  data_out[2191] = data_in[1437];
     assign  data_out[2192] = data_in[1413];
     assign  data_out[2193] = data_in[767];
     assign  data_out[2194] = data_in[1294];
     assign  data_out[2195] = data_in[1687];
     assign  data_out[2196] = data_in[521];
     assign  data_out[2197] = data_in[870];
     assign  data_out[2198] = data_in[452];
     assign  data_out[2199] = data_in[1209];
     assign  data_out[2200] = data_in[571];
     assign  data_out[2201] = data_in[1480];
     assign  data_out[2202] = data_in[1312];
     assign  data_out[2203] = data_in[1570];
     assign  data_out[2204] = data_in[848];
     assign  data_out[2205] = data_in[583];
     assign  data_out[2206] = data_in[801];
     assign  data_out[2207] = data_in[432];
     assign  data_out[2208] = data_in[694];
     assign  data_out[2209] = data_in[1562];
     assign  data_out[2210] = data_in[959];
     assign  data_out[2211] = data_in[926];
     assign  data_out[2212] = data_in[122];
     assign  data_out[2213] = data_in[1214];
     assign  data_out[2214] = data_in[1013];
     assign  data_out[2215] = data_in[1076];
     assign  data_out[2216] = data_in[1518];
     assign  data_out[2217] = data_in[410];
     assign  data_out[2218] = data_in[1056];
     assign  data_out[2219] = data_in[267];
     assign  data_out[2220] = data_in[1695];
     assign  data_out[2221] = data_in[494];
     assign  data_out[2222] = data_in[99];
     assign  data_out[2223] = data_in[116];
     assign  data_out[2224] = data_in[709];
     assign  data_out[2225] = data_in[1252];
     assign  data_out[2226] = data_in[1510];
     assign  data_out[2227] = data_in[473];
     assign  data_out[2228] = data_in[1127];
     assign  data_out[2229] = data_in[1593];
     assign  data_out[2230] = data_in[1700];
     assign  data_out[2231] = data_in[737];
     assign  data_out[2232] = data_in[1700];
     assign  data_out[2233] = data_in[1462];
     assign  data_out[2234] = data_in[998];
     assign  data_out[2235] = data_in[284];
     assign  data_out[2236] = data_in[613];
     assign  data_out[2237] = data_in[959];
     assign  data_out[2238] = data_in[475];
     assign  data_out[2239] = data_in[1305];
     assign  data_out[2240] = data_in[146];
     assign  data_out[2241] = data_in[371];
     assign  data_out[2242] = data_in[1184];
     assign  data_out[2243] = data_in[923];
     assign  data_out[2244] = data_in[296];
     assign  data_out[2245] = data_in[544];
     assign  data_out[2246] = data_in[693];
     assign  data_out[2247] = data_in[91];
     assign  data_out[2248] = data_in[828];
     assign  data_out[2249] = data_in[379];
     assign  data_out[2250] = data_in[1651];
     assign  data_out[2251] = data_in[570];
     assign  data_out[2252] = data_in[1027];
     assign  data_out[2253] = data_in[1259];
     assign  data_out[2254] = data_in[1331];
     assign  data_out[2255] = data_in[226];
     assign  data_out[2256] = data_in[1085];
     assign  data_out[2257] = data_in[1373];
     assign  data_out[2258] = data_in[1095];
     assign  data_out[2259] = data_in[1145];
     assign  data_out[2260] = data_in[1293];
     assign  data_out[2261] = data_in[89];
     assign  data_out[2262] = data_in[1265];
     assign  data_out[2263] = data_in[1038];
     assign  data_out[2264] = data_in[1244];
     assign  data_out[2265] = data_in[547];
     assign  data_out[2266] = data_in[1330];
     assign  data_out[2267] = data_in[1481];
     assign  data_out[2268] = data_in[412];
     assign  data_out[2269] = data_in[1247];
     assign  data_out[2270] = data_in[359];
     assign  data_out[2271] = data_in[1700];
     assign  data_out[2272] = data_in[574];
     assign  data_out[2273] = data_in[1073];
     assign  data_out[2274] = data_in[270];
     assign  data_out[2275] = data_in[1089];
     assign  data_out[2276] = data_in[1076];
     assign  data_out[2277] = data_in[1634];
     assign  data_out[2278] = data_in[1629];
     assign  data_out[2279] = data_in[1648];
     assign  data_out[2280] = data_in[1236];
     assign  data_out[2281] = data_in[256];
     assign  data_out[2282] = data_in[1553];
     assign  data_out[2283] = data_in[674];
     assign  data_out[2284] = data_in[879];
     assign  data_out[2285] = data_in[696];
     assign  data_out[2286] = data_in[668];
     assign  data_out[2287] = data_in[1204];
     assign  data_out[2288] = data_in[1213];
     assign  data_out[2289] = data_in[366];
     assign  data_out[2290] = data_in[1045];
     assign  data_out[2291] = data_in[1144];
     assign  data_out[2292] = data_in[480];
     assign  data_out[2293] = data_in[135];
     assign  data_out[2294] = data_in[339];
     assign  data_out[2295] = data_in[695];
     assign  data_out[2296] = data_in[426];
     assign  data_out[2297] = data_in[684];
     assign  data_out[2298] = data_in[346];
     assign  data_out[2299] = data_in[1105];
     assign  data_out[2300] = data_in[746];
     assign  data_out[2301] = data_in[381];
     assign  data_out[2302] = data_in[632];
     assign  data_out[2303] = data_in[1512];
     assign  data_out[2304] = data_in[1001];
     assign  data_out[2305] = data_in[123];
     assign  data_out[2306] = data_in[643];
     assign  data_out[2307] = data_in[1485];
     assign  data_out[2308] = data_in[978];
     assign  data_out[2309] = data_in[731];
     assign  data_out[2310] = data_in[1691];
     assign  data_out[2311] = data_in[470];
     assign  data_out[2312] = data_in[1723];
     assign  data_out[2313] = data_in[73];
     assign  data_out[2314] = data_in[1097];
     assign  data_out[2315] = data_in[7];
     assign  data_out[2316] = data_in[1671];
     assign  data_out[2317] = data_in[1434];
     assign  data_out[2318] = data_in[1017];
     assign  data_out[2319] = data_in[1673];
     assign  data_out[2320] = data_in[466];
     assign  data_out[2321] = data_in[545];
     assign  data_out[2322] = data_in[33];
     assign  data_out[2323] = data_in[1427];
     assign  data_out[2324] = data_in[1442];
     assign  data_out[2325] = data_in[813];
     assign  data_out[2326] = data_in[384];
     assign  data_out[2327] = data_in[941];
     assign  data_out[2328] = data_in[1168];
     assign  data_out[2329] = data_in[1716];
     assign  data_out[2330] = data_in[676];
     assign  data_out[2331] = data_in[341];
     assign  data_out[2332] = data_in[225];
     assign  data_out[2333] = data_in[1235];
     assign  data_out[2334] = data_in[15];
     assign  data_out[2335] = data_in[1553];
     assign  data_out[2336] = data_in[1150];
     assign  data_out[2337] = data_in[510];
     assign  data_out[2338] = data_in[682];
     assign  data_out[2339] = data_in[501];
     assign  data_out[2340] = data_in[84];
     assign  data_out[2341] = data_in[1477];
     assign  data_out[2342] = data_in[748];
     assign  data_out[2343] = data_in[839];
     assign  data_out[2344] = data_in[245];
     assign  data_out[2345] = data_in[1213];
     assign  data_out[2346] = data_in[23];
     assign  data_out[2347] = data_in[1507];
     assign  data_out[2348] = data_in[204];
     assign  data_out[2349] = data_in[1407];
     assign  data_out[2350] = data_in[370];
     assign  data_out[2351] = data_in[1178];
     assign  data_out[2352] = data_in[645];
     assign  data_out[2353] = data_in[388];
     assign  data_out[2354] = data_in[1323];
     assign  data_out[2355] = data_in[1271];
     assign  data_out[2356] = data_in[1588];
     assign  data_out[2357] = data_in[1689];
     assign  data_out[2358] = data_in[1404];
     assign  data_out[2359] = data_in[466];
     assign  data_out[2360] = data_in[914];
     assign  data_out[2361] = data_in[1380];
     assign  data_out[2362] = data_in[900];
     assign  data_out[2363] = data_in[426];
     assign  data_out[2364] = data_in[751];
     assign  data_out[2365] = data_in[256];
     assign  data_out[2366] = data_in[956];
     assign  data_out[2367] = data_in[96];
     assign  data_out[2368] = data_in[1447];
     assign  data_out[2369] = data_in[1389];
     assign  data_out[2370] = data_in[1624];
     assign  data_out[2371] = data_in[36];
     assign  data_out[2372] = data_in[41];
     assign  data_out[2373] = data_in[1092];
     assign  data_out[2374] = data_in[666];
     assign  data_out[2375] = data_in[1044];
     assign  data_out[2376] = data_in[643];
     assign  data_out[2377] = data_in[1225];
     assign  data_out[2378] = data_in[933];
     assign  data_out[2379] = data_in[1255];
     assign  data_out[2380] = data_in[28];
     assign  data_out[2381] = data_in[762];
     assign  data_out[2382] = data_in[446];
     assign  data_out[2383] = data_in[179];
     assign  data_out[2384] = data_in[801];
     assign  data_out[2385] = data_in[1456];
     assign  data_out[2386] = data_in[674];
     assign  data_out[2387] = data_in[12];
     assign  data_out[2388] = data_in[1620];
     assign  data_out[2389] = data_in[1088];
     assign  data_out[2390] = data_in[215];
     assign  data_out[2391] = data_in[611];
     assign  data_out[2392] = data_in[1264];
     assign  data_out[2393] = data_in[492];
     assign  data_out[2394] = data_in[732];
     assign  data_out[2395] = data_in[922];
     assign  data_out[2396] = data_in[612];
     assign  data_out[2397] = data_in[1292];
     assign  data_out[2398] = data_in[988];
     assign  data_out[2399] = data_in[1519];
     assign  data_out[2400] = data_in[1291];
     assign  data_out[2401] = data_in[1536];
     assign  data_out[2402] = data_in[659];
     assign  data_out[2403] = data_in[314];
     assign  data_out[2404] = data_in[607];
     assign  data_out[2405] = data_in[734];
     assign  data_out[2406] = data_in[127];
     assign  data_out[2407] = data_in[289];
     assign  data_out[2408] = data_in[548];
     assign  data_out[2409] = data_in[735];
     assign  data_out[2410] = data_in[653];
     assign  data_out[2411] = data_in[569];
     assign  data_out[2412] = data_in[1077];
     assign  data_out[2413] = data_in[133];
     assign  data_out[2414] = data_in[1505];
     assign  data_out[2415] = data_in[55];
     assign  data_out[2416] = data_in[683];
     assign  data_out[2417] = data_in[1471];
     assign  data_out[2418] = data_in[162];
     assign  data_out[2419] = data_in[493];
     assign  data_out[2420] = data_in[349];
     assign  data_out[2421] = data_in[1277];
     assign  data_out[2422] = data_in[819];
     assign  data_out[2423] = data_in[175];
     assign  data_out[2424] = data_in[1063];
     assign  data_out[2425] = data_in[1218];
     assign  data_out[2426] = data_in[1018];
     assign  data_out[2427] = data_in[1448];
     assign  data_out[2428] = data_in[1388];
     assign  data_out[2429] = data_in[34];
     assign  data_out[2430] = data_in[1370];
     assign  data_out[2431] = data_in[747];
     assign  data_out[2432] = data_in[784];
     assign  data_out[2433] = data_in[1080];
     assign  data_out[2434] = data_in[1294];
     assign  data_out[2435] = data_in[1614];
     assign  data_out[2436] = data_in[1376];
     assign  data_out[2437] = data_in[322];
     assign  data_out[2438] = data_in[1538];
     assign  data_out[2439] = data_in[426];
     assign  data_out[2440] = data_in[21];
     assign  data_out[2441] = data_in[1720];
     assign  data_out[2442] = data_in[597];
     assign  data_out[2443] = data_in[821];
     assign  data_out[2444] = data_in[1393];
     assign  data_out[2445] = data_in[639];
     assign  data_out[2446] = data_in[621];
     assign  data_out[2447] = data_in[1375];
     assign  data_out[2448] = data_in[744];
     assign  data_out[2449] = data_in[1236];
     assign  data_out[2450] = data_in[1268];
     assign  data_out[2451] = data_in[427];
     assign  data_out[2452] = data_in[1612];
     assign  data_out[2453] = data_in[1552];
     assign  data_out[2454] = data_in[573];
     assign  data_out[2455] = data_in[605];
     assign  data_out[2456] = data_in[1588];
     assign  data_out[2457] = data_in[161];
     assign  data_out[2458] = data_in[284];
     assign  data_out[2459] = data_in[1675];
     assign  data_out[2460] = data_in[1039];
     assign  data_out[2461] = data_in[1301];
     assign  data_out[2462] = data_in[176];
     assign  data_out[2463] = data_in[536];
     assign  data_out[2464] = data_in[729];
     assign  data_out[2465] = data_in[1496];
     assign  data_out[2466] = data_in[1257];
     assign  data_out[2467] = data_in[813];
     assign  data_out[2468] = data_in[54];
     assign  data_out[2469] = data_in[258];
     assign  data_out[2470] = data_in[662];
     assign  data_out[2471] = data_in[768];
     assign  data_out[2472] = data_in[1553];
     assign  data_out[2473] = data_in[593];
     assign  data_out[2474] = data_in[1585];
     assign  data_out[2475] = data_in[1710];
     assign  data_out[2476] = data_in[585];
     assign  data_out[2477] = data_in[429];
     assign  data_out[2478] = data_in[322];
     assign  data_out[2479] = data_in[444];
     assign  data_out[2480] = data_in[410];
     assign  data_out[2481] = data_in[1174];
     assign  data_out[2482] = data_in[1425];
     assign  data_out[2483] = data_in[1039];
     assign  data_out[2484] = data_in[440];
     assign  data_out[2485] = data_in[1697];
     assign  data_out[2486] = data_in[561];
     assign  data_out[2487] = data_in[810];
     assign  data_out[2488] = data_in[1362];
     assign  data_out[2489] = data_in[458];
     assign  data_out[2490] = data_in[1647];
     assign  data_out[2491] = data_in[1328];
     assign  data_out[2492] = data_in[822];
     assign  data_out[2493] = data_in[28];
     assign  data_out[2494] = data_in[932];
     assign  data_out[2495] = data_in[1104];
     assign  data_out[2496] = data_in[905];
     assign  data_out[2497] = data_in[428];
     assign  data_out[2498] = data_in[1141];
     assign  data_out[2499] = data_in[26];
     assign  data_out[2500] = data_in[1098];
     assign  data_out[2501] = data_in[1434];
     assign  data_out[2502] = data_in[447];
     assign  data_out[2503] = data_in[1548];
     assign  data_out[2504] = data_in[1426];
     assign  data_out[2505] = data_in[304];
     assign  data_out[2506] = data_in[388];
     assign  data_out[2507] = data_in[1260];
     assign  data_out[2508] = data_in[1557];
     assign  data_out[2509] = data_in[1594];
     assign  data_out[2510] = data_in[1679];
     assign  data_out[2511] = data_in[1392];
     assign  data_out[2512] = data_in[1539];
     assign  data_out[2513] = data_in[1332];
     assign  data_out[2514] = data_in[927];
     assign  data_out[2515] = data_in[151];
     assign  data_out[2516] = data_in[344];
     assign  data_out[2517] = data_in[251];
     assign  data_out[2518] = data_in[408];
     assign  data_out[2519] = data_in[617];
     assign  data_out[2520] = data_in[1336];
     assign  data_out[2521] = data_in[1413];
     assign  data_out[2522] = data_in[715];
     assign  data_out[2523] = data_in[186];
     assign  data_out[2524] = data_in[103];
     assign  data_out[2525] = data_in[279];
     assign  data_out[2526] = data_in[525];
     assign  data_out[2527] = data_in[132];
     assign  data_out[2528] = data_in[63];
     assign  data_out[2529] = data_in[324];
     assign  data_out[2530] = data_in[942];
     assign  data_out[2531] = data_in[1421];
     assign  data_out[2532] = data_in[159];
     assign  data_out[2533] = data_in[40];
     assign  data_out[2534] = data_in[654];
     assign  data_out[2535] = data_in[459];
     assign  data_out[2536] = data_in[78];
     assign  data_out[2537] = data_in[1695];
     assign  data_out[2538] = data_in[95];
     assign  data_out[2539] = data_in[1005];
     assign  data_out[2540] = data_in[137];
     assign  data_out[2541] = data_in[1527];
     assign  data_out[2542] = data_in[848];
     assign  data_out[2543] = data_in[633];
     assign  data_out[2544] = data_in[1506];
     assign  data_out[2545] = data_in[1377];
     assign  data_out[2546] = data_in[1201];
     assign  data_out[2547] = data_in[822];
     assign  data_out[2548] = data_in[1216];
     assign  data_out[2549] = data_in[1426];
     assign  data_out[2550] = data_in[10];
     assign  data_out[2551] = data_in[769];
     assign  data_out[2552] = data_in[1436];
     assign  data_out[2553] = data_in[224];
     assign  data_out[2554] = data_in[1144];
     assign  data_out[2555] = data_in[1539];
     assign  data_out[2556] = data_in[1543];
     assign  data_out[2557] = data_in[1417];
     assign  data_out[2558] = data_in[1293];
     assign  data_out[2559] = data_in[1401];
     assign  data_out[2560] = data_in[1113];
     assign  data_out[2561] = data_in[1529];
     assign  data_out[2562] = data_in[63];
     assign  data_out[2563] = data_in[311];
     assign  data_out[2564] = data_in[1370];
     assign  data_out[2565] = data_in[1395];
     assign  data_out[2566] = data_in[1313];
     assign  data_out[2567] = data_in[1297];
     assign  data_out[2568] = data_in[379];
     assign  data_out[2569] = data_in[46];
     assign  data_out[2570] = data_in[1472];
     assign  data_out[2571] = data_in[806];
     assign  data_out[2572] = data_in[632];
     assign  data_out[2573] = data_in[1564];
     assign  data_out[2574] = data_in[1168];
     assign  data_out[2575] = data_in[678];
     assign  data_out[2576] = data_in[114];
     assign  data_out[2577] = data_in[600];
     assign  data_out[2578] = data_in[1355];
     assign  data_out[2579] = data_in[983];
     assign  data_out[2580] = data_in[1058];
     assign  data_out[2581] = data_in[1279];
     assign  data_out[2582] = data_in[1261];
     assign  data_out[2583] = data_in[1202];
     assign  data_out[2584] = data_in[563];
     assign  data_out[2585] = data_in[621];
     assign  data_out[2586] = data_in[811];
     assign  data_out[2587] = data_in[91];
     assign  data_out[2588] = data_in[725];
     assign  data_out[2589] = data_in[1564];
     assign  data_out[2590] = data_in[662];
     assign  data_out[2591] = data_in[972];
     assign  data_out[2592] = data_in[754];
     assign  data_out[2593] = data_in[550];
     assign  data_out[2594] = data_in[769];
     assign  data_out[2595] = data_in[699];
     assign  data_out[2596] = data_in[59];
     assign  data_out[2597] = data_in[933];
     assign  data_out[2598] = data_in[998];
     assign  data_out[2599] = data_in[134];
     assign  data_out[2600] = data_in[716];
     assign  data_out[2601] = data_in[629];
     assign  data_out[2602] = data_in[1235];
     assign  data_out[2603] = data_in[577];
     assign  data_out[2604] = data_in[275];
     assign  data_out[2605] = data_in[70];
     assign  data_out[2606] = data_in[1062];
     assign  data_out[2607] = data_in[1503];
     assign  data_out[2608] = data_in[1326];
     assign  data_out[2609] = data_in[1368];
     assign  data_out[2610] = data_in[1627];
     assign  data_out[2611] = data_in[345];
     assign  data_out[2612] = data_in[1167];
     assign  data_out[2613] = data_in[1536];
     assign  data_out[2614] = data_in[1142];
     assign  data_out[2615] = data_in[1040];
     assign  data_out[2616] = data_in[46];
     assign  data_out[2617] = data_in[775];
     assign  data_out[2618] = data_in[457];
     assign  data_out[2619] = data_in[966];
     assign  data_out[2620] = data_in[1716];
     assign  data_out[2621] = data_in[1057];
     assign  data_out[2622] = data_in[1511];
     assign  data_out[2623] = data_in[1007];
     assign  data_out[2624] = data_in[1572];
     assign  data_out[2625] = data_in[431];
     assign  data_out[2626] = data_in[1275];
     assign  data_out[2627] = data_in[1460];
     assign  data_out[2628] = data_in[35];
     assign  data_out[2629] = data_in[1489];
     assign  data_out[2630] = data_in[278];
     assign  data_out[2631] = data_in[876];
     assign  data_out[2632] = data_in[179];
     assign  data_out[2633] = data_in[1422];
     assign  data_out[2634] = data_in[691];
     assign  data_out[2635] = data_in[286];
     assign  data_out[2636] = data_in[1320];
     assign  data_out[2637] = data_in[1080];
     assign  data_out[2638] = data_in[953];
     assign  data_out[2639] = data_in[546];
     assign  data_out[2640] = data_in[1168];
     assign  data_out[2641] = data_in[488];
     assign  data_out[2642] = data_in[1665];
     assign  data_out[2643] = data_in[401];
     assign  data_out[2644] = data_in[949];
     assign  data_out[2645] = data_in[954];
     assign  data_out[2646] = data_in[357];
     assign  data_out[2647] = data_in[326];
     assign  data_out[2648] = data_in[191];
     assign  data_out[2649] = data_in[205];
     assign  data_out[2650] = data_in[226];
     assign  data_out[2651] = data_in[704];
     assign  data_out[2652] = data_in[1504];
     assign  data_out[2653] = data_in[718];
     assign  data_out[2654] = data_in[77];
     assign  data_out[2655] = data_in[1130];
     assign  data_out[2656] = data_in[1671];
     assign  data_out[2657] = data_in[381];
     assign  data_out[2658] = data_in[931];
     assign  data_out[2659] = data_in[1523];
     assign  data_out[2660] = data_in[1487];
     assign  data_out[2661] = data_in[1199];
     assign  data_out[2662] = data_in[1724];
     assign  data_out[2663] = data_in[1430];
     assign  data_out[2664] = data_in[285];
     assign  data_out[2665] = data_in[30];
     assign  data_out[2666] = data_in[553];
     assign  data_out[2667] = data_in[1685];
     assign  data_out[2668] = data_in[678];
     assign  data_out[2669] = data_in[475];
     assign  data_out[2670] = data_in[1533];
     assign  data_out[2671] = data_in[1344];
     assign  data_out[2672] = data_in[1549];
     assign  data_out[2673] = data_in[1300];
     assign  data_out[2674] = data_in[519];
     assign  data_out[2675] = data_in[973];
     assign  data_out[2676] = data_in[1378];
     assign  data_out[2677] = data_in[503];
     assign  data_out[2678] = data_in[1610];
     assign  data_out[2679] = data_in[20];
     assign  data_out[2680] = data_in[275];
     assign  data_out[2681] = data_in[1509];
     assign  data_out[2682] = data_in[1399];
     assign  data_out[2683] = data_in[1082];
     assign  data_out[2684] = data_in[374];
     assign  data_out[2685] = data_in[128];
     assign  data_out[2686] = data_in[1508];
     assign  data_out[2687] = data_in[155];
     assign  data_out[2688] = data_in[1584];
     assign  data_out[2689] = data_in[958];
     assign  data_out[2690] = data_in[218];
     assign  data_out[2691] = data_in[1599];
     assign  data_out[2692] = data_in[986];
     assign  data_out[2693] = data_in[412];
     assign  data_out[2694] = data_in[1261];
     assign  data_out[2695] = data_in[626];
     assign  data_out[2696] = data_in[1529];
     assign  data_out[2697] = data_in[588];
     assign  data_out[2698] = data_in[940];
     assign  data_out[2699] = data_in[1393];
     assign  data_out[2700] = data_in[278];
     assign  data_out[2701] = data_in[1535];
     assign  data_out[2702] = data_in[309];
     assign  data_out[2703] = data_in[1444];
     assign  data_out[2704] = data_in[1627];
     assign  data_out[2705] = data_in[1580];
     assign  data_out[2706] = data_in[104];
     assign  data_out[2707] = data_in[205];
     assign  data_out[2708] = data_in[1534];
     assign  data_out[2709] = data_in[1641];
     assign  data_out[2710] = data_in[964];
     assign  data_out[2711] = data_in[274];
     assign  data_out[2712] = data_in[278];
     assign  data_out[2713] = data_in[1721];
     assign  data_out[2714] = data_in[1204];
     assign  data_out[2715] = data_in[476];
     assign  data_out[2716] = data_in[175];
     assign  data_out[2717] = data_in[1080];
     assign  data_out[2718] = data_in[853];
     assign  data_out[2719] = data_in[1269];
     assign  data_out[2720] = data_in[819];
     assign  data_out[2721] = data_in[616];
     assign  data_out[2722] = data_in[756];
     assign  data_out[2723] = data_in[726];
     assign  data_out[2724] = data_in[126];
     assign  data_out[2725] = data_in[1692];
     assign  data_out[2726] = data_in[270];
     assign  data_out[2727] = data_in[1664];
     assign  data_out[2728] = data_in[1650];
     assign  data_out[2729] = data_in[1670];
     assign  data_out[2730] = data_in[1375];
     assign  data_out[2731] = data_in[1268];
     assign  data_out[2732] = data_in[162];
     assign  data_out[2733] = data_in[1113];
     assign  data_out[2734] = data_in[241];
     assign  data_out[2735] = data_in[1036];
     assign  data_out[2736] = data_in[1260];
     assign  data_out[2737] = data_in[458];
     assign  data_out[2738] = data_in[13];
     assign  data_out[2739] = data_in[1482];
     assign  data_out[2740] = data_in[339];
     assign  data_out[2741] = data_in[1125];
     assign  data_out[2742] = data_in[1662];
     assign  data_out[2743] = data_in[427];
     assign  data_out[2744] = data_in[883];
     assign  data_out[2745] = data_in[955];
     assign  data_out[2746] = data_in[1462];
     assign  data_out[2747] = data_in[770];
     assign  data_out[2748] = data_in[867];
     assign  data_out[2749] = data_in[670];
     assign  data_out[2750] = data_in[343];
     assign  data_out[2751] = data_in[1668];
     assign  data_out[2752] = data_in[1314];
     assign  data_out[2753] = data_in[886];
     assign  data_out[2754] = data_in[109];
     assign  data_out[2755] = data_in[1449];
     assign  data_out[2756] = data_in[338];
     assign  data_out[2757] = data_in[1177];
     assign  data_out[2758] = data_in[403];
     assign  data_out[2759] = data_in[24];
     assign  data_out[2760] = data_in[817];
     assign  data_out[2761] = data_in[1475];
     assign  data_out[2762] = data_in[789];
     assign  data_out[2763] = data_in[1495];
     assign  data_out[2764] = data_in[209];
     assign  data_out[2765] = data_in[4];
     assign  data_out[2766] = data_in[1102];
     assign  data_out[2767] = data_in[1230];
     assign  data_out[2768] = data_in[1009];
     assign  data_out[2769] = data_in[140];
     assign  data_out[2770] = data_in[971];
     assign  data_out[2771] = data_in[1330];
     assign  data_out[2772] = data_in[7];
     assign  data_out[2773] = data_in[1386];
     assign  data_out[2774] = data_in[306];
     assign  data_out[2775] = data_in[738];
     assign  data_out[2776] = data_in[17];
     assign  data_out[2777] = data_in[676];
     assign  data_out[2778] = data_in[1669];
     assign  data_out[2779] = data_in[449];
     assign  data_out[2780] = data_in[521];
     assign  data_out[2781] = data_in[1666];
     assign  data_out[2782] = data_in[751];
     assign  data_out[2783] = data_in[1192];
     assign  data_out[2784] = data_in[525];
     assign  data_out[2785] = data_in[1192];
     assign  data_out[2786] = data_in[436];
     assign  data_out[2787] = data_in[1185];
     assign  data_out[2788] = data_in[1163];
     assign  data_out[2789] = data_in[674];
     assign  data_out[2790] = data_in[123];
     assign  data_out[2791] = data_in[744];
     assign  data_out[2792] = data_in[1628];
     assign  data_out[2793] = data_in[1275];
     assign  data_out[2794] = data_in[975];
     assign  data_out[2795] = data_in[584];
     assign  data_out[2796] = data_in[135];
     assign  data_out[2797] = data_in[1218];
     assign  data_out[2798] = data_in[1210];
     assign  data_out[2799] = data_in[597];
     assign  data_out[2800] = data_in[409];
     assign  data_out[2801] = data_in[725];
     assign  data_out[2802] = data_in[1381];
     assign  data_out[2803] = data_in[1512];
     assign  data_out[2804] = data_in[862];
     assign  data_out[2805] = data_in[153];
     assign  data_out[2806] = data_in[679];
     assign  data_out[2807] = data_in[656];
     assign  data_out[2808] = data_in[1495];
     assign  data_out[2809] = data_in[240];
     assign  data_out[2810] = data_in[730];
     assign  data_out[2811] = data_in[1506];
     assign  data_out[2812] = data_in[500];
     assign  data_out[2813] = data_in[407];
     assign  data_out[2814] = data_in[1394];
     assign  data_out[2815] = data_in[597];
     assign  data_out[2816] = data_in[64];
     assign  data_out[2817] = data_in[582];
     assign  data_out[2818] = data_in[1571];
     assign  data_out[2819] = data_in[863];
     assign  data_out[2820] = data_in[253];
     assign  data_out[2821] = data_in[749];
     assign  data_out[2822] = data_in[1623];
     assign  data_out[2823] = data_in[1140];
     assign  data_out[2824] = data_in[474];
     assign  data_out[2825] = data_in[239];
     assign  data_out[2826] = data_in[1404];
     assign  data_out[2827] = data_in[557];
     assign  data_out[2828] = data_in[1223];
     assign  data_out[2829] = data_in[1336];
     assign  data_out[2830] = data_in[879];
     assign  data_out[2831] = data_in[353];
     assign  data_out[2832] = data_in[1423];
     assign  data_out[2833] = data_in[207];
     assign  data_out[2834] = data_in[783];
     assign  data_out[2835] = data_in[389];
     assign  data_out[2836] = data_in[1340];
     assign  data_out[2837] = data_in[828];
     assign  data_out[2838] = data_in[1652];
     assign  data_out[2839] = data_in[547];
     assign  data_out[2840] = data_in[1194];
     assign  data_out[2841] = data_in[354];
     assign  data_out[2842] = data_in[409];
     assign  data_out[2843] = data_in[804];
     assign  data_out[2844] = data_in[279];
     assign  data_out[2845] = data_in[631];
     assign  data_out[2846] = data_in[127];
     assign  data_out[2847] = data_in[1562];
     assign  data_out[2848] = data_in[521];
     assign  data_out[2849] = data_in[1181];
     assign  data_out[2850] = data_in[1028];
     assign  data_out[2851] = data_in[1461];
     assign  data_out[2852] = data_in[282];
     assign  data_out[2853] = data_in[727];
     assign  data_out[2854] = data_in[450];
     assign  data_out[2855] = data_in[1173];
     assign  data_out[2856] = data_in[1357];
     assign  data_out[2857] = data_in[614];
     assign  data_out[2858] = data_in[952];
     assign  data_out[2859] = data_in[30];
     assign  data_out[2860] = data_in[1139];
     assign  data_out[2861] = data_in[886];
     assign  data_out[2862] = data_in[693];
     assign  data_out[2863] = data_in[906];
     assign  data_out[2864] = data_in[1536];
     assign  data_out[2865] = data_in[1387];
     assign  data_out[2866] = data_in[1577];
     assign  data_out[2867] = data_in[1563];
     assign  data_out[2868] = data_in[1439];
     assign  data_out[2869] = data_in[384];
     assign  data_out[2870] = data_in[636];
     assign  data_out[2871] = data_in[1697];
     assign  data_out[2872] = data_in[874];
     assign  data_out[2873] = data_in[1349];
     assign  data_out[2874] = data_in[152];
     assign  data_out[2875] = data_in[445];
     assign  data_out[2876] = data_in[896];
     assign  data_out[2877] = data_in[1379];
     assign  data_out[2878] = data_in[263];
     assign  data_out[2879] = data_in[1495];
     assign  data_out[2880] = data_in[1455];
     assign  data_out[2881] = data_in[1279];
     assign  data_out[2882] = data_in[909];
     assign  data_out[2883] = data_in[560];
     assign  data_out[2884] = data_in[304];
     assign  data_out[2885] = data_in[416];
     assign  data_out[2886] = data_in[1064];
     assign  data_out[2887] = data_in[1722];
     assign  data_out[2888] = data_in[343];
     assign  data_out[2889] = data_in[813];
     assign  data_out[2890] = data_in[1357];
     assign  data_out[2891] = data_in[1132];
     assign  data_out[2892] = data_in[841];
     assign  data_out[2893] = data_in[878];
     assign  data_out[2894] = data_in[1506];
     assign  data_out[2895] = data_in[125];
     assign  data_out[2896] = data_in[659];
     assign  data_out[2897] = data_in[1502];
     assign  data_out[2898] = data_in[383];
     assign  data_out[2899] = data_in[47];
     assign  data_out[2900] = data_in[999];
     assign  data_out[2901] = data_in[1467];
     assign  data_out[2902] = data_in[497];
     assign  data_out[2903] = data_in[1123];
     assign  data_out[2904] = data_in[1273];
     assign  data_out[2905] = data_in[1448];
     assign  data_out[2906] = data_in[534];
     assign  data_out[2907] = data_in[855];
     assign  data_out[2908] = data_in[1502];
     assign  data_out[2909] = data_in[449];
     assign  data_out[2910] = data_in[198];
     assign  data_out[2911] = data_in[452];
     assign  data_out[2912] = data_in[1404];
     assign  data_out[2913] = data_in[518];
     assign  data_out[2914] = data_in[996];
     assign  data_out[2915] = data_in[976];
     assign  data_out[2916] = data_in[941];
     assign  data_out[2917] = data_in[112];
     assign  data_out[2918] = data_in[1281];
     assign  data_out[2919] = data_in[1129];
     assign  data_out[2920] = data_in[1111];
     assign  data_out[2921] = data_in[597];
     assign  data_out[2922] = data_in[308];
     assign  data_out[2923] = data_in[862];
     assign  data_out[2924] = data_in[1127];
     assign  data_out[2925] = data_in[1081];
     assign  data_out[2926] = data_in[987];
     assign  data_out[2927] = data_in[253];
     assign  data_out[2928] = data_in[1135];
     assign  data_out[2929] = data_in[868];
     assign  data_out[2930] = data_in[143];
     assign  data_out[2931] = data_in[1277];
     assign  data_out[2932] = data_in[1425];
     assign  data_out[2933] = data_in[296];
     assign  data_out[2934] = data_in[915];
     assign  data_out[2935] = data_in[218];
     assign  data_out[2936] = data_in[372];
     assign  data_out[2937] = data_in[223];
     assign  data_out[2938] = data_in[1540];
     assign  data_out[2939] = data_in[788];
     assign  data_out[2940] = data_in[1086];
     assign  data_out[2941] = data_in[1309];
     assign  data_out[2942] = data_in[329];
     assign  data_out[2943] = data_in[1137];
     assign  data_out[2944] = data_in[1333];
     assign  data_out[2945] = data_in[1616];
     assign  data_out[2946] = data_in[476];
     assign  data_out[2947] = data_in[396];
     assign  data_out[2948] = data_in[925];
     assign  data_out[2949] = data_in[597];
     assign  data_out[2950] = data_in[915];
     assign  data_out[2951] = data_in[382];
     assign  data_out[2952] = data_in[1129];
     assign  data_out[2953] = data_in[1079];
     assign  data_out[2954] = data_in[84];
     assign  data_out[2955] = data_in[1457];
     assign  data_out[2956] = data_in[902];
     assign  data_out[2957] = data_in[22];
     assign  data_out[2958] = data_in[530];
     assign  data_out[2959] = data_in[995];
     assign  data_out[2960] = data_in[825];
     assign  data_out[2961] = data_in[1152];
     assign  data_out[2962] = data_in[1475];
     assign  data_out[2963] = data_in[374];
     assign  data_out[2964] = data_in[502];
     assign  data_out[2965] = data_in[487];
     assign  data_out[2966] = data_in[112];
     assign  data_out[2967] = data_in[1294];
     assign  data_out[2968] = data_in[312];
     assign  data_out[2969] = data_in[328];
     assign  data_out[2970] = data_in[830];
     assign  data_out[2971] = data_in[780];
     assign  data_out[2972] = data_in[200];
     assign  data_out[2973] = data_in[1001];
     assign  data_out[2974] = data_in[1320];
     assign  data_out[2975] = data_in[257];
     assign  data_out[2976] = data_in[1181];
     assign  data_out[2977] = data_in[3];
     assign  data_out[2978] = data_in[1397];
     assign  data_out[2979] = data_in[16];
     assign  data_out[2980] = data_in[553];
     assign  data_out[2981] = data_in[1412];
     assign  data_out[2982] = data_in[53];
     assign  data_out[2983] = data_in[1387];
     assign  data_out[2984] = data_in[297];
     assign  data_out[2985] = data_in[1266];
     assign  data_out[2986] = data_in[641];
     assign  data_out[2987] = data_in[21];
     assign  data_out[2988] = data_in[641];
     assign  data_out[2989] = data_in[171];
     assign  data_out[2990] = data_in[71];
     assign  data_out[2991] = data_in[1246];
     assign  data_out[2992] = data_in[19];
     assign  data_out[2993] = data_in[185];
     assign  data_out[2994] = data_in[946];
     assign  data_out[2995] = data_in[1154];
     assign  data_out[2996] = data_in[1038];
     assign  data_out[2997] = data_in[959];
     assign  data_out[2998] = data_in[35];
     assign  data_out[2999] = data_in[666];
     assign  data_out[3000] = data_in[479];
     assign  data_out[3001] = data_in[579];
     assign  data_out[3002] = data_in[658];
     assign  data_out[3003] = data_in[1420];
     assign  data_out[3004] = data_in[964];
     assign  data_out[3005] = data_in[510];
     assign  data_out[3006] = data_in[650];
     assign  data_out[3007] = data_in[621];
     assign  data_out[3008] = data_in[1590];
     assign  data_out[3009] = data_in[1097];
     assign  data_out[3010] = data_in[31];
     assign  data_out[3011] = data_in[1088];
     assign  data_out[3012] = data_in[1689];
     assign  data_out[3013] = data_in[852];
     assign  data_out[3014] = data_in[776];
     assign  data_out[3015] = data_in[55];
     assign  data_out[3016] = data_in[945];
     assign  data_out[3017] = data_in[1515];
     assign  data_out[3018] = data_in[1341];
     assign  data_out[3019] = data_in[629];
     assign  data_out[3020] = data_in[654];
     assign  data_out[3021] = data_in[1027];
     assign  data_out[3022] = data_in[1544];
     assign  data_out[3023] = data_in[820];
     assign  data_out[3024] = data_in[1439];
     assign  data_out[3025] = data_in[605];
     assign  data_out[3026] = data_in[1442];
     assign  data_out[3027] = data_in[576];
     assign  data_out[3028] = data_in[498];
     assign  data_out[3029] = data_in[1117];
     assign  data_out[3030] = data_in[1175];
     assign  data_out[3031] = data_in[752];
     assign  data_out[3032] = data_in[961];
     assign  data_out[3033] = data_in[1144];
     assign  data_out[3034] = data_in[952];
     assign  data_out[3035] = data_in[1622];
     assign  data_out[3036] = data_in[154];
     assign  data_out[3037] = data_in[1306];
     assign  data_out[3038] = data_in[1254];
     assign  data_out[3039] = data_in[775];
     assign  data_out[3040] = data_in[448];
     assign  data_out[3041] = data_in[1301];
     assign  data_out[3042] = data_in[695];
     assign  data_out[3043] = data_in[1461];
     assign  data_out[3044] = data_in[849];
     assign  data_out[3045] = data_in[1160];
     assign  data_out[3046] = data_in[254];
     assign  data_out[3047] = data_in[127];
     assign  data_out[3048] = data_in[919];
     assign  data_out[3049] = data_in[75];
     assign  data_out[3050] = data_in[954];
     assign  data_out[3051] = data_in[493];
     assign  data_out[3052] = data_in[1089];
     assign  data_out[3053] = data_in[848];
     assign  data_out[3054] = data_in[242];
     assign  data_out[3055] = data_in[447];
     assign  data_out[3056] = data_in[1594];
     assign  data_out[3057] = data_in[1217];
     assign  data_out[3058] = data_in[72];
     assign  data_out[3059] = data_in[836];
     assign  data_out[3060] = data_in[1364];
     assign  data_out[3061] = data_in[851];
     assign  data_out[3062] = data_in[834];
     assign  data_out[3063] = data_in[1435];
     assign  data_out[3064] = data_in[820];
     assign  data_out[3065] = data_in[83];
     assign  data_out[3066] = data_in[1047];
     assign  data_out[3067] = data_in[358];
     assign  data_out[3068] = data_in[1292];
     assign  data_out[3069] = data_in[160];
     assign  data_out[3070] = data_in[1149];
     assign  data_out[3071] = data_in[180];
     assign  data_out[3072] = data_in[1528];
     assign  data_out[3073] = data_in[91];
     assign  data_out[3074] = data_in[200];
     assign  data_out[3075] = data_in[765];
     assign  data_out[3076] = data_in[1302];
     assign  data_out[3077] = data_in[1603];
     assign  data_out[3078] = data_in[1109];
     assign  data_out[3079] = data_in[1080];
     assign  data_out[3080] = data_in[496];
     assign  data_out[3081] = data_in[3];
     assign  data_out[3082] = data_in[1110];
     assign  data_out[3083] = data_in[340];
     assign  data_out[3084] = data_in[206];
     assign  data_out[3085] = data_in[103];
     assign  data_out[3086] = data_in[367];
     assign  data_out[3087] = data_in[49];
     assign  data_out[3088] = data_in[1154];
     assign  data_out[3089] = data_in[445];
     assign  data_out[3090] = data_in[262];
     assign  data_out[3091] = data_in[726];
     assign  data_out[3092] = data_in[775];
     assign  data_out[3093] = data_in[538];
     assign  data_out[3094] = data_in[44];
     assign  data_out[3095] = data_in[56];
     assign  data_out[3096] = data_in[1549];
     assign  data_out[3097] = data_in[266];
     assign  data_out[3098] = data_in[1414];
     assign  data_out[3099] = data_in[105];
     assign  data_out[3100] = data_in[829];
     assign  data_out[3101] = data_in[1244];
     assign  data_out[3102] = data_in[354];
     assign  data_out[3103] = data_in[945];
     assign  data_out[3104] = data_in[666];
     assign  data_out[3105] = data_in[26];
     assign  data_out[3106] = data_in[1674];
     assign  data_out[3107] = data_in[413];
     assign  data_out[3108] = data_in[968];
     assign  data_out[3109] = data_in[210];
     assign  data_out[3110] = data_in[1050];
     assign  data_out[3111] = data_in[1578];
     assign  data_out[3112] = data_in[656];
     assign  data_out[3113] = data_in[522];
     assign  data_out[3114] = data_in[1117];
     assign  data_out[3115] = data_in[946];
     assign  data_out[3116] = data_in[1286];
     assign  data_out[3117] = data_in[1480];
     assign  data_out[3118] = data_in[1208];
     assign  data_out[3119] = data_in[465];
     assign  data_out[3120] = data_in[1490];
     assign  data_out[3121] = data_in[1524];
     assign  data_out[3122] = data_in[1387];
     assign  data_out[3123] = data_in[823];
     assign  data_out[3124] = data_in[892];
     assign  data_out[3125] = data_in[1041];
     assign  data_out[3126] = data_in[103];
     assign  data_out[3127] = data_in[60];
     assign  data_out[3128] = data_in[157];
     assign  data_out[3129] = data_in[725];
     assign  data_out[3130] = data_in[200];
     assign  data_out[3131] = data_in[1670];
     assign  data_out[3132] = data_in[236];
     assign  data_out[3133] = data_in[574];
     assign  data_out[3134] = data_in[884];
     assign  data_out[3135] = data_in[911];
     assign  data_out[3136] = data_in[1313];
     assign  data_out[3137] = data_in[1557];
     assign  data_out[3138] = data_in[742];
     assign  data_out[3139] = data_in[145];
     assign  data_out[3140] = data_in[1063];
     assign  data_out[3141] = data_in[679];
     assign  data_out[3142] = data_in[1511];
     assign  data_out[3143] = data_in[1206];
     assign  data_out[3144] = data_in[1352];
     assign  data_out[3145] = data_in[477];
     assign  data_out[3146] = data_in[1418];
     assign  data_out[3147] = data_in[1416];
     assign  data_out[3148] = data_in[536];
     assign  data_out[3149] = data_in[1236];
     assign  data_out[3150] = data_in[594];
     assign  data_out[3151] = data_in[1724];
     assign  data_out[3152] = data_in[1217];
     assign  data_out[3153] = data_in[393];
     assign  data_out[3154] = data_in[502];
     assign  data_out[3155] = data_in[29];
     assign  data_out[3156] = data_in[257];
     assign  data_out[3157] = data_in[253];
     assign  data_out[3158] = data_in[853];
     assign  data_out[3159] = data_in[626];
     assign  data_out[3160] = data_in[1269];
     assign  data_out[3161] = data_in[115];
     assign  data_out[3162] = data_in[142];
     assign  data_out[3163] = data_in[728];
     assign  data_out[3164] = data_in[823];
     assign  data_out[3165] = data_in[1563];
     assign  data_out[3166] = data_in[1568];
     assign  data_out[3167] = data_in[567];
     assign  data_out[3168] = data_in[706];
     assign  data_out[3169] = data_in[1300];
     assign  data_out[3170] = data_in[1071];
     assign  data_out[3171] = data_in[1480];
     assign  data_out[3172] = data_in[913];
     assign  data_out[3173] = data_in[280];
     assign  data_out[3174] = data_in[743];
     assign  data_out[3175] = data_in[465];
     assign  data_out[3176] = data_in[1512];
     assign  data_out[3177] = data_in[60];
     assign  data_out[3178] = data_in[133];
     assign  data_out[3179] = data_in[909];
     assign  data_out[3180] = data_in[912];
     assign  data_out[3181] = data_in[1302];
     assign  data_out[3182] = data_in[82];
     assign  data_out[3183] = data_in[1316];
     assign  data_out[3184] = data_in[1383];
     assign  data_out[3185] = data_in[1257];
     assign  data_out[3186] = data_in[979];
     assign  data_out[3187] = data_in[755];
     assign  data_out[3188] = data_in[707];
     assign  data_out[3189] = data_in[9];
     assign  data_out[3190] = data_in[679];
     assign  data_out[3191] = data_in[121];
     assign  data_out[3192] = data_in[1571];
     assign  data_out[3193] = data_in[170];
     assign  data_out[3194] = data_in[1656];
     assign  data_out[3195] = data_in[1647];
     assign  data_out[3196] = data_in[283];
     assign  data_out[3197] = data_in[1201];
     assign  data_out[3198] = data_in[1505];
     assign  data_out[3199] = data_in[1318];
     assign  data_out[3200] = data_in[245];
     assign  data_out[3201] = data_in[678];
     assign  data_out[3202] = data_in[554];
     assign  data_out[3203] = data_in[810];
     assign  data_out[3204] = data_in[1409];
     assign  data_out[3205] = data_in[229];
     assign  data_out[3206] = data_in[718];
     assign  data_out[3207] = data_in[775];
     assign  data_out[3208] = data_in[763];
     assign  data_out[3209] = data_in[818];
     assign  data_out[3210] = data_in[1701];
     assign  data_out[3211] = data_in[365];
     assign  data_out[3212] = data_in[26];
     assign  data_out[3213] = data_in[635];
     assign  data_out[3214] = data_in[1499];
     assign  data_out[3215] = data_in[1108];
     assign  data_out[3216] = data_in[279];
     assign  data_out[3217] = data_in[1031];
     assign  data_out[3218] = data_in[411];
     assign  data_out[3219] = data_in[284];
     assign  data_out[3220] = data_in[459];
     assign  data_out[3221] = data_in[900];
     assign  data_out[3222] = data_in[1690];
     assign  data_out[3223] = data_in[1290];
     assign  data_out[3224] = data_in[178];
     assign  data_out[3225] = data_in[518];
     assign  data_out[3226] = data_in[1108];
     assign  data_out[3227] = data_in[212];
     assign  data_out[3228] = data_in[1329];
     assign  data_out[3229] = data_in[416];
     assign  data_out[3230] = data_in[65];
     assign  data_out[3231] = data_in[305];
     assign  data_out[3232] = data_in[301];
     assign  data_out[3233] = data_in[737];
     assign  data_out[3234] = data_in[1670];
     assign  data_out[3235] = data_in[1492];
     assign  data_out[3236] = data_in[1552];
     assign  data_out[3237] = data_in[497];
     assign  data_out[3238] = data_in[227];
     assign  data_out[3239] = data_in[1017];
     assign  data_out[3240] = data_in[1166];
     assign  data_out[3241] = data_in[461];
     assign  data_out[3242] = data_in[1327];
     assign  data_out[3243] = data_in[778];
     assign  data_out[3244] = data_in[510];
     assign  data_out[3245] = data_in[411];
     assign  data_out[3246] = data_in[28];
     assign  data_out[3247] = data_in[425];
     assign  data_out[3248] = data_in[358];
     assign  data_out[3249] = data_in[1434];
     assign  data_out[3250] = data_in[984];
     assign  data_out[3251] = data_in[1136];
     assign  data_out[3252] = data_in[1027];
     assign  data_out[3253] = data_in[550];
     assign  data_out[3254] = data_in[1081];
     assign  data_out[3255] = data_in[879];
     assign  data_out[3256] = data_in[367];
     assign  data_out[3257] = data_in[409];
     assign  data_out[3258] = data_in[1180];
     assign  data_out[3259] = data_in[900];
     assign  data_out[3260] = data_in[1329];
     assign  data_out[3261] = data_in[626];
     assign  data_out[3262] = data_in[343];
     assign  data_out[3263] = data_in[771];
     assign  data_out[3264] = data_in[219];
     assign  data_out[3265] = data_in[415];
     assign  data_out[3266] = data_in[1124];
     assign  data_out[3267] = data_in[24];
     assign  data_out[3268] = data_in[182];
     assign  data_out[3269] = data_in[1541];
     assign  data_out[3270] = data_in[56];
     assign  data_out[3271] = data_in[991];
     assign  data_out[3272] = data_in[297];
     assign  data_out[3273] = data_in[1505];
     assign  data_out[3274] = data_in[533];
     assign  data_out[3275] = data_in[1469];
     assign  data_out[3276] = data_in[1380];
     assign  data_out[3277] = data_in[559];
     assign  data_out[3278] = data_in[1492];
     assign  data_out[3279] = data_in[1242];
     assign  data_out[3280] = data_in[1316];
     assign  data_out[3281] = data_in[352];
     assign  data_out[3282] = data_in[830];
     assign  data_out[3283] = data_in[699];
     assign  data_out[3284] = data_in[305];
     assign  data_out[3285] = data_in[524];
     assign  data_out[3286] = data_in[1503];
     assign  data_out[3287] = data_in[13];
     assign  data_out[3288] = data_in[927];
     assign  data_out[3289] = data_in[440];
     assign  data_out[3290] = data_in[507];
     assign  data_out[3291] = data_in[1329];
     assign  data_out[3292] = data_in[945];
     assign  data_out[3293] = data_in[277];
     assign  data_out[3294] = data_in[520];
     assign  data_out[3295] = data_in[1690];
     assign  data_out[3296] = data_in[48];
     assign  data_out[3297] = data_in[2];
     assign  data_out[3298] = data_in[208];
     assign  data_out[3299] = data_in[1600];
     assign  data_out[3300] = data_in[1160];
     assign  data_out[3301] = data_in[849];
     assign  data_out[3302] = data_in[1261];
     assign  data_out[3303] = data_in[1415];
     assign  data_out[3304] = data_in[1621];
     assign  data_out[3305] = data_in[904];
     assign  data_out[3306] = data_in[247];
     assign  data_out[3307] = data_in[84];
     assign  data_out[3308] = data_in[1487];
     assign  data_out[3309] = data_in[1497];
     assign  data_out[3310] = data_in[1615];
     assign  data_out[3311] = data_in[1266];
     assign  data_out[3312] = data_in[94];
     assign  data_out[3313] = data_in[477];
     assign  data_out[3314] = data_in[946];
     assign  data_out[3315] = data_in[1603];
     assign  data_out[3316] = data_in[1208];
     assign  data_out[3317] = data_in[1144];
     assign  data_out[3318] = data_in[692];
     assign  data_out[3319] = data_in[732];
     assign  data_out[3320] = data_in[1354];
     assign  data_out[3321] = data_in[835];
     assign  data_out[3322] = data_in[585];
     assign  data_out[3323] = data_in[902];
     assign  data_out[3324] = data_in[677];
     assign  data_out[3325] = data_in[29];
     assign  data_out[3326] = data_in[776];
     assign  data_out[3327] = data_in[1230];
     assign  data_out[3328] = data_in[536];
     assign  data_out[3329] = data_in[1136];
     assign  data_out[3330] = data_in[1349];
     assign  data_out[3331] = data_in[1098];
     assign  data_out[3332] = data_in[1274];
     assign  data_out[3333] = data_in[1579];
     assign  data_out[3334] = data_in[1715];
     assign  data_out[3335] = data_in[468];
     assign  data_out[3336] = data_in[661];
     assign  data_out[3337] = data_in[419];
     assign  data_out[3338] = data_in[805];
     assign  data_out[3339] = data_in[1235];
     assign  data_out[3340] = data_in[1252];
     assign  data_out[3341] = data_in[673];
     assign  data_out[3342] = data_in[1576];
     assign  data_out[3343] = data_in[848];
     assign  data_out[3344] = data_in[1251];
     assign  data_out[3345] = data_in[667];
     assign  data_out[3346] = data_in[6];
     assign  data_out[3347] = data_in[1344];
     assign  data_out[3348] = data_in[1309];
     assign  data_out[3349] = data_in[1491];
     assign  data_out[3350] = data_in[109];
     assign  data_out[3351] = data_in[809];
     assign  data_out[3352] = data_in[116];
     assign  data_out[3353] = data_in[1437];
     assign  data_out[3354] = data_in[586];
     assign  data_out[3355] = data_in[802];
     assign  data_out[3356] = data_in[863];
     assign  data_out[3357] = data_in[1027];
     assign  data_out[3358] = data_in[1559];
     assign  data_out[3359] = data_in[201];
     assign  data_out[3360] = data_in[1407];
     assign  data_out[3361] = data_in[1622];
     assign  data_out[3362] = data_in[1196];
     assign  data_out[3363] = data_in[363];
     assign  data_out[3364] = data_in[605];
     assign  data_out[3365] = data_in[463];
     assign  data_out[3366] = data_in[1284];
     assign  data_out[3367] = data_in[703];
     assign  data_out[3368] = data_in[557];
     assign  data_out[3369] = data_in[1433];
     assign  data_out[3370] = data_in[218];
     assign  data_out[3371] = data_in[949];
     assign  data_out[3372] = data_in[931];
     assign  data_out[3373] = data_in[1203];
     assign  data_out[3374] = data_in[1094];
     assign  data_out[3375] = data_in[1262];
     assign  data_out[3376] = data_in[1404];
     assign  data_out[3377] = data_in[1131];
     assign  data_out[3378] = data_in[1274];
     assign  data_out[3379] = data_in[932];
     assign  data_out[3380] = data_in[1470];
     assign  data_out[3381] = data_in[1132];
     assign  data_out[3382] = data_in[1486];
     assign  data_out[3383] = data_in[666];
     assign  data_out[3384] = data_in[1567];
     assign  data_out[3385] = data_in[1710];
     assign  data_out[3386] = data_in[818];
     assign  data_out[3387] = data_in[539];
     assign  data_out[3388] = data_in[1679];
     assign  data_out[3389] = data_in[1450];
     assign  data_out[3390] = data_in[134];
     assign  data_out[3391] = data_in[336];
     assign  data_out[3392] = data_in[1360];
     assign  data_out[3393] = data_in[616];
     assign  data_out[3394] = data_in[989];
     assign  data_out[3395] = data_in[1294];
     assign  data_out[3396] = data_in[800];
     assign  data_out[3397] = data_in[1630];
     assign  data_out[3398] = data_in[109];
     assign  data_out[3399] = data_in[409];
     assign  data_out[3400] = data_in[1694];
     assign  data_out[3401] = data_in[1494];
     assign  data_out[3402] = data_in[1089];
     assign  data_out[3403] = data_in[490];
     assign  data_out[3404] = data_in[619];
     assign  data_out[3405] = data_in[1507];
     assign  data_out[3406] = data_in[161];
     assign  data_out[3407] = data_in[1239];
     assign  data_out[3408] = data_in[1331];
     assign  data_out[3409] = data_in[1697];
     assign  data_out[3410] = data_in[509];
     assign  data_out[3411] = data_in[1426];
     assign  data_out[3412] = data_in[667];
     assign  data_out[3413] = data_in[119];
     assign  data_out[3414] = data_in[1640];
     assign  data_out[3415] = data_in[1642];
     assign  data_out[3416] = data_in[395];
     assign  data_out[3417] = data_in[743];
     assign  data_out[3418] = data_in[995];
     assign  data_out[3419] = data_in[1402];
     assign  data_out[3420] = data_in[1411];
     assign  data_out[3421] = data_in[1686];
     assign  data_out[3422] = data_in[945];
     assign  data_out[3423] = data_in[824];
     assign  data_out[3424] = data_in[1522];
     assign  data_out[3425] = data_in[350];
     assign  data_out[3426] = data_in[1372];
     assign  data_out[3427] = data_in[660];
     assign  data_out[3428] = data_in[1618];
     assign  data_out[3429] = data_in[1056];
     assign  data_out[3430] = data_in[325];
     assign  data_out[3431] = data_in[519];
     assign  data_out[3432] = data_in[1704];
     assign  data_out[3433] = data_in[1229];
     assign  data_out[3434] = data_in[244];
     assign  data_out[3435] = data_in[1177];
     assign  data_out[3436] = data_in[250];
     assign  data_out[3437] = data_in[490];
     assign  data_out[3438] = data_in[763];
     assign  data_out[3439] = data_in[431];
     assign  data_out[3440] = data_in[781];
     assign  data_out[3441] = data_in[91];
     assign  data_out[3442] = data_in[1513];
     assign  data_out[3443] = data_in[489];
     assign  data_out[3444] = data_in[1168];
     assign  data_out[3445] = data_in[720];
     assign  data_out[3446] = data_in[1117];
     assign  data_out[3447] = data_in[809];
     assign  data_out[3448] = data_in[630];
     assign  data_out[3449] = data_in[701];
     assign  data_out[3450] = data_in[236];
     assign  data_out[3451] = data_in[1283];
     assign  data_out[3452] = data_in[1638];
     assign  data_out[3453] = data_in[883];
     assign  data_out[3454] = data_in[68];
     assign  data_out[3455] = data_in[50];
     assign  data_out[3456] = data_in[266];
     assign  data_out[3457] = data_in[952];
     assign  data_out[3458] = data_in[668];
     assign  data_out[3459] = data_in[467];
     assign  data_out[3460] = data_in[925];
     assign  data_out[3461] = data_in[388];
     assign  data_out[3462] = data_in[885];
     assign  data_out[3463] = data_in[1156];
     assign  data_out[3464] = data_in[648];
     assign  data_out[3465] = data_in[885];
     assign  data_out[3466] = data_in[824];
     assign  data_out[3467] = data_in[925];
     assign  data_out[3468] = data_in[1320];
     assign  data_out[3469] = data_in[999];
     assign  data_out[3470] = data_in[1705];
     assign  data_out[3471] = data_in[1135];
     assign  data_out[3472] = data_in[208];
     assign  data_out[3473] = data_in[569];
     assign  data_out[3474] = data_in[586];
     assign  data_out[3475] = data_in[1017];
     assign  data_out[3476] = data_in[1623];
     assign  data_out[3477] = data_in[503];
     assign  data_out[3478] = data_in[729];
     assign  data_out[3479] = data_in[1342];
     assign  data_out[3480] = data_in[93];
     assign  data_out[3481] = data_in[1644];
     assign  data_out[3482] = data_in[524];
     assign  data_out[3483] = data_in[1580];
     assign  data_out[3484] = data_in[323];
     assign  data_out[3485] = data_in[405];
     assign  data_out[3486] = data_in[760];
     assign  data_out[3487] = data_in[768];
     assign  data_out[3488] = data_in[124];
     assign  data_out[3489] = data_in[442];
     assign  data_out[3490] = data_in[63];
     assign  data_out[3491] = data_in[1049];
     assign  data_out[3492] = data_in[1610];
     assign  data_out[3493] = data_in[28];
     assign  data_out[3494] = data_in[1008];
     assign  data_out[3495] = data_in[1635];
     assign  data_out[3496] = data_in[1016];
     assign  data_out[3497] = data_in[334];
     assign  data_out[3498] = data_in[193];
     assign  data_out[3499] = data_in[1162];
     assign  data_out[3500] = data_in[1713];
     assign  data_out[3501] = data_in[1184];
     assign  data_out[3502] = data_in[329];
     assign  data_out[3503] = data_in[1382];
     assign  data_out[3504] = data_in[766];
     assign  data_out[3505] = data_in[101];
     assign  data_out[3506] = data_in[342];
     assign  data_out[3507] = data_in[778];
     assign  data_out[3508] = data_in[520];
     assign  data_out[3509] = data_in[978];
     assign  data_out[3510] = data_in[1559];
     assign  data_out[3511] = data_in[420];
     assign  data_out[3512] = data_in[761];
     assign  data_out[3513] = data_in[1524];
     assign  data_out[3514] = data_in[1516];
     assign  data_out[3515] = data_in[290];
     assign  data_out[3516] = data_in[449];
     assign  data_out[3517] = data_in[371];
     assign  data_out[3518] = data_in[1365];
     assign  data_out[3519] = data_in[1469];
     assign  data_out[3520] = data_in[875];
     assign  data_out[3521] = data_in[1647];
     assign  data_out[3522] = data_in[147];
     assign  data_out[3523] = data_in[1065];
     assign  data_out[3524] = data_in[1218];
     assign  data_out[3525] = data_in[866];
     assign  data_out[3526] = data_in[185];
     assign  data_out[3527] = data_in[458];
     assign  data_out[3528] = data_in[819];
     assign  data_out[3529] = data_in[796];
     assign  data_out[3530] = data_in[307];
     assign  data_out[3531] = data_in[1639];
     assign  data_out[3532] = data_in[875];
     assign  data_out[3533] = data_in[1407];
     assign  data_out[3534] = data_in[1163];
     assign  data_out[3535] = data_in[121];
     assign  data_out[3536] = data_in[856];
     assign  data_out[3537] = data_in[460];
     assign  data_out[3538] = data_in[1078];
     assign  data_out[3539] = data_in[1050];
     assign  data_out[3540] = data_in[1371];
     assign  data_out[3541] = data_in[687];
     assign  data_out[3542] = data_in[1507];
     assign  data_out[3543] = data_in[1328];
     assign  data_out[3544] = data_in[132];
     assign  data_out[3545] = data_in[1374];
     assign  data_out[3546] = data_in[552];
     assign  data_out[3547] = data_in[650];
     assign  data_out[3548] = data_in[1383];
     assign  data_out[3549] = data_in[1388];
     assign  data_out[3550] = data_in[495];
     assign  data_out[3551] = data_in[1561];
     assign  data_out[3552] = data_in[1268];
     assign  data_out[3553] = data_in[104];
     assign  data_out[3554] = data_in[918];
     assign  data_out[3555] = data_in[955];
     assign  data_out[3556] = data_in[585];
     assign  data_out[3557] = data_in[822];
     assign  data_out[3558] = data_in[1634];
     assign  data_out[3559] = data_in[504];
     assign  data_out[3560] = data_in[494];
     assign  data_out[3561] = data_in[1385];
     assign  data_out[3562] = data_in[798];
     assign  data_out[3563] = data_in[435];
     assign  data_out[3564] = data_in[1546];
     assign  data_out[3565] = data_in[790];
     assign  data_out[3566] = data_in[362];
     assign  data_out[3567] = data_in[675];
     assign  data_out[3568] = data_in[1309];
     assign  data_out[3569] = data_in[1313];
     assign  data_out[3570] = data_in[763];
     assign  data_out[3571] = data_in[1437];
     assign  data_out[3572] = data_in[612];
     assign  data_out[3573] = data_in[384];
     assign  data_out[3574] = data_in[468];
     assign  data_out[3575] = data_in[1353];
     assign  data_out[3576] = data_in[1586];
     assign  data_out[3577] = data_in[119];
     assign  data_out[3578] = data_in[1286];
     assign  data_out[3579] = data_in[764];
     assign  data_out[3580] = data_in[600];
     assign  data_out[3581] = data_in[1092];
     assign  data_out[3582] = data_in[489];
     assign  data_out[3583] = data_in[1370];
     assign  data_out[3584] = data_in[759];
     assign  data_out[3585] = data_in[1341];
     assign  data_out[3586] = data_in[50];
     assign  data_out[3587] = data_in[1213];
     assign  data_out[3588] = data_in[387];
     assign  data_out[3589] = data_in[30];
     assign  data_out[3590] = data_in[200];
     assign  data_out[3591] = data_in[384];
     assign  data_out[3592] = data_in[1184];
     assign  data_out[3593] = data_in[839];
     assign  data_out[3594] = data_in[705];
     assign  data_out[3595] = data_in[867];
     assign  data_out[3596] = data_in[1122];
     assign  data_out[3597] = data_in[669];
     assign  data_out[3598] = data_in[1265];
     assign  data_out[3599] = data_in[373];
     assign  data_out[3600] = data_in[201];
     assign  data_out[3601] = data_in[224];
     assign  data_out[3602] = data_in[233];
     assign  data_out[3603] = data_in[1597];
     assign  data_out[3604] = data_in[1428];
     assign  data_out[3605] = data_in[1310];
     assign  data_out[3606] = data_in[335];
     assign  data_out[3607] = data_in[430];
     assign  data_out[3608] = data_in[568];
     assign  data_out[3609] = data_in[1491];
     assign  data_out[3610] = data_in[1596];
     assign  data_out[3611] = data_in[519];
     assign  data_out[3612] = data_in[599];
     assign  data_out[3613] = data_in[1060];
     assign  data_out[3614] = data_in[503];
     assign  data_out[3615] = data_in[412];
     assign  data_out[3616] = data_in[1231];
     assign  data_out[3617] = data_in[138];
     assign  data_out[3618] = data_in[1537];
     assign  data_out[3619] = data_in[662];
     assign  data_out[3620] = data_in[1138];
     assign  data_out[3621] = data_in[838];
     assign  data_out[3622] = data_in[1369];
     assign  data_out[3623] = data_in[1356];
     assign  data_out[3624] = data_in[1275];
     assign  data_out[3625] = data_in[971];
     assign  data_out[3626] = data_in[199];
     assign  data_out[3627] = data_in[1120];
     assign  data_out[3628] = data_in[291];
     assign  data_out[3629] = data_in[1136];
     assign  data_out[3630] = data_in[568];
     assign  data_out[3631] = data_in[920];
     assign  data_out[3632] = data_in[1495];
     assign  data_out[3633] = data_in[1288];
     assign  data_out[3634] = data_in[1455];
     assign  data_out[3635] = data_in[1241];
     assign  data_out[3636] = data_in[1661];
     assign  data_out[3637] = data_in[8];
     assign  data_out[3638] = data_in[1545];
     assign  data_out[3639] = data_in[1140];
     assign  data_out[3640] = data_in[137];
     assign  data_out[3641] = data_in[202];
     assign  data_out[3642] = data_in[494];
     assign  data_out[3643] = data_in[1586];
     assign  data_out[3644] = data_in[258];
     assign  data_out[3645] = data_in[1630];
     assign  data_out[3646] = data_in[1685];
     assign  data_out[3647] = data_in[849];
     assign  data_out[3648] = data_in[86];
     assign  data_out[3649] = data_in[1266];
     assign  data_out[3650] = data_in[138];
     assign  data_out[3651] = data_in[1632];
     assign  data_out[3652] = data_in[1460];
     assign  data_out[3653] = data_in[894];
     assign  data_out[3654] = data_in[528];
     assign  data_out[3655] = data_in[410];
     assign  data_out[3656] = data_in[1585];
     assign  data_out[3657] = data_in[1489];
     assign  data_out[3658] = data_in[589];
     assign  data_out[3659] = data_in[1163];
     assign  data_out[3660] = data_in[1308];
     assign  data_out[3661] = data_in[1042];
     assign  data_out[3662] = data_in[422];
     assign  data_out[3663] = data_in[1478];
     assign  data_out[3664] = data_in[1216];
     assign  data_out[3665] = data_in[1311];
     assign  data_out[3666] = data_in[619];
     assign  data_out[3667] = data_in[136];
     assign  data_out[3668] = data_in[717];
     assign  data_out[3669] = data_in[418];
     assign  data_out[3670] = data_in[1347];
     assign  data_out[3671] = data_in[69];
     assign  data_out[3672] = data_in[596];
     assign  data_out[3673] = data_in[957];
     assign  data_out[3674] = data_in[1581];
     assign  data_out[3675] = data_in[503];
     assign  data_out[3676] = data_in[25];
     assign  data_out[3677] = data_in[168];
     assign  data_out[3678] = data_in[275];
     assign  data_out[3679] = data_in[578];
     assign  data_out[3680] = data_in[610];
     assign  data_out[3681] = data_in[478];
     assign  data_out[3682] = data_in[386];
     assign  data_out[3683] = data_in[1323];
     assign  data_out[3684] = data_in[1544];
     assign  data_out[3685] = data_in[64];
     assign  data_out[3686] = data_in[245];
     assign  data_out[3687] = data_in[642];
     assign  data_out[3688] = data_in[177];
     assign  data_out[3689] = data_in[1725];
     assign  data_out[3690] = data_in[857];
     assign  data_out[3691] = data_in[1018];
     assign  data_out[3692] = data_in[1083];
     assign  data_out[3693] = data_in[1454];
     assign  data_out[3694] = data_in[1518];
     assign  data_out[3695] = data_in[405];
     assign  data_out[3696] = data_in[1274];
     assign  data_out[3697] = data_in[176];
     assign  data_out[3698] = data_in[234];
     assign  data_out[3699] = data_in[1558];
     assign  data_out[3700] = data_in[1295];
     assign  data_out[3701] = data_in[55];
     assign  data_out[3702] = data_in[717];
     assign  data_out[3703] = data_in[1634];
     assign  data_out[3704] = data_in[1223];
     assign  data_out[3705] = data_in[1168];
     assign  data_out[3706] = data_in[952];
     assign  data_out[3707] = data_in[776];
     assign  data_out[3708] = data_in[183];
     assign  data_out[3709] = data_in[1437];
     assign  data_out[3710] = data_in[1418];
     assign  data_out[3711] = data_in[140];
     assign  data_out[3712] = data_in[1611];
     assign  data_out[3713] = data_in[62];
     assign  data_out[3714] = data_in[1035];
     assign  data_out[3715] = data_in[447];
     assign  data_out[3716] = data_in[1417];
     assign  data_out[3717] = data_in[425];
     assign  data_out[3718] = data_in[1631];
     assign  data_out[3719] = data_in[878];
     assign  data_out[3720] = data_in[1000];
     assign  data_out[3721] = data_in[631];
     assign  data_out[3722] = data_in[1123];
     assign  data_out[3723] = data_in[762];
     assign  data_out[3724] = data_in[1546];
     assign  data_out[3725] = data_in[465];
     assign  data_out[3726] = data_in[1363];
     assign  data_out[3727] = data_in[428];
     assign  data_out[3728] = data_in[826];
     assign  data_out[3729] = data_in[847];
     assign  data_out[3730] = data_in[486];
     assign  data_out[3731] = data_in[195];
     assign  data_out[3732] = data_in[752];
     assign  data_out[3733] = data_in[376];
     assign  data_out[3734] = data_in[901];
     assign  data_out[3735] = data_in[801];
     assign  data_out[3736] = data_in[272];
     assign  data_out[3737] = data_in[1328];
     assign  data_out[3738] = data_in[1022];
     assign  data_out[3739] = data_in[779];
     assign  data_out[3740] = data_in[854];
     assign  data_out[3741] = data_in[320];
     assign  data_out[3742] = data_in[166];
     assign  data_out[3743] = data_in[996];
     assign  data_out[3744] = data_in[867];
     assign  data_out[3745] = data_in[197];
     assign  data_out[3746] = data_in[247];
     assign  data_out[3747] = data_in[1496];
     assign  data_out[3748] = data_in[943];
     assign  data_out[3749] = data_in[1084];
     assign  data_out[3750] = data_in[883];
     assign  data_out[3751] = data_in[864];
     assign  data_out[3752] = data_in[65];
     assign  data_out[3753] = data_in[238];
     assign  data_out[3754] = data_in[912];
     assign  data_out[3755] = data_in[525];
     assign  data_out[3756] = data_in[1011];
     assign  data_out[3757] = data_in[114];
     assign  data_out[3758] = data_in[1190];
     assign  data_out[3759] = data_in[11];
     assign  data_out[3760] = data_in[1458];
     assign  data_out[3761] = data_in[722];
     assign  data_out[3762] = data_in[966];
     assign  data_out[3763] = data_in[1161];
     assign  data_out[3764] = data_in[1463];
     assign  data_out[3765] = data_in[1596];
     assign  data_out[3766] = data_in[1686];
     assign  data_out[3767] = data_in[368];
     assign  data_out[3768] = data_in[152];
     assign  data_out[3769] = data_in[1550];
     assign  data_out[3770] = data_in[154];
     assign  data_out[3771] = data_in[672];
     assign  data_out[3772] = data_in[269];
     assign  data_out[3773] = data_in[826];
     assign  data_out[3774] = data_in[475];
     assign  data_out[3775] = data_in[340];
     assign  data_out[3776] = data_in[316];
     assign  data_out[3777] = data_in[688];
     assign  data_out[3778] = data_in[773];
     assign  data_out[3779] = data_in[106];
     assign  data_out[3780] = data_in[1556];
     assign  data_out[3781] = data_in[1635];
     assign  data_out[3782] = data_in[1380];
     assign  data_out[3783] = data_in[1264];
     assign  data_out[3784] = data_in[997];
     assign  data_out[3785] = data_in[469];
     assign  data_out[3786] = data_in[881];
     assign  data_out[3787] = data_in[492];
     assign  data_out[3788] = data_in[1083];
     assign  data_out[3789] = data_in[1196];
     assign  data_out[3790] = data_in[772];
     assign  data_out[3791] = data_in[263];
     assign  data_out[3792] = data_in[276];
     assign  data_out[3793] = data_in[281];
     assign  data_out[3794] = data_in[673];
     assign  data_out[3795] = data_in[981];
     assign  data_out[3796] = data_in[458];
     assign  data_out[3797] = data_in[959];
     assign  data_out[3798] = data_in[1403];
     assign  data_out[3799] = data_in[592];
     assign  data_out[3800] = data_in[518];
     assign  data_out[3801] = data_in[1569];
     assign  data_out[3802] = data_in[1301];
     assign  data_out[3803] = data_in[664];
     assign  data_out[3804] = data_in[1684];
     assign  data_out[3805] = data_in[535];
     assign  data_out[3806] = data_in[1393];
     assign  data_out[3807] = data_in[1467];
     assign  data_out[3808] = data_in[870];
     assign  data_out[3809] = data_in[959];
     assign  data_out[3810] = data_in[1314];
     assign  data_out[3811] = data_in[605];
     assign  data_out[3812] = data_in[1067];
     assign  data_out[3813] = data_in[431];
     assign  data_out[3814] = data_in[1587];
     assign  data_out[3815] = data_in[203];
     assign  data_out[3816] = data_in[1212];
     assign  data_out[3817] = data_in[872];
     assign  data_out[3818] = data_in[1096];
     assign  data_out[3819] = data_in[900];
     assign  data_out[3820] = data_in[1481];
     assign  data_out[3821] = data_in[1535];
     assign  data_out[3822] = data_in[155];
     assign  data_out[3823] = data_in[1483];
     assign  data_out[3824] = data_in[270];
     assign  data_out[3825] = data_in[1350];
     assign  data_out[3826] = data_in[1467];
     assign  data_out[3827] = data_in[1418];
     assign  data_out[3828] = data_in[1518];
     assign  data_out[3829] = data_in[1380];
     assign  data_out[3830] = data_in[379];
     assign  data_out[3831] = data_in[923];
     assign  data_out[3832] = data_in[2];
     assign  data_out[3833] = data_in[743];
     assign  data_out[3834] = data_in[1639];
     assign  data_out[3835] = data_in[1022];
     assign  data_out[3836] = data_in[1277];
     assign  data_out[3837] = data_in[974];
     assign  data_out[3838] = data_in[506];
     assign  data_out[3839] = data_in[1680];
     assign  data_out[3840] = data_in[687];
     assign  data_out[3841] = data_in[57];
     assign  data_out[3842] = data_in[1704];
     assign  data_out[3843] = data_in[464];
     assign  data_out[3844] = data_in[584];
     assign  data_out[3845] = data_in[1492];
     assign  data_out[3846] = data_in[237];
     assign  data_out[3847] = data_in[181];
     assign  data_out[3848] = data_in[554];
     assign  data_out[3849] = data_in[614];
     assign  data_out[3850] = data_in[1026];
     assign  data_out[3851] = data_in[315];
     assign  data_out[3852] = data_in[30];
     assign  data_out[3853] = data_in[1171];
     assign  data_out[3854] = data_in[1379];
     assign  data_out[3855] = data_in[1433];
     assign  data_out[3856] = data_in[1677];
     assign  data_out[3857] = data_in[197];
     assign  data_out[3858] = data_in[1157];
     assign  data_out[3859] = data_in[835];
     assign  data_out[3860] = data_in[1349];
     assign  data_out[3861] = data_in[1075];
     assign  data_out[3862] = data_in[939];
     assign  data_out[3863] = data_in[1727];
     assign  data_out[3864] = data_in[1392];
     assign  data_out[3865] = data_in[1508];
     assign  data_out[3866] = data_in[1205];
     assign  data_out[3867] = data_in[336];
     assign  data_out[3868] = data_in[251];
     assign  data_out[3869] = data_in[696];
     assign  data_out[3870] = data_in[856];
     assign  data_out[3871] = data_in[928];
     assign  data_out[3872] = data_in[354];
     assign  data_out[3873] = data_in[108];
     assign  data_out[3874] = data_in[1186];
     assign  data_out[3875] = data_in[663];
     assign  data_out[3876] = data_in[1054];
     assign  data_out[3877] = data_in[686];
     assign  data_out[3878] = data_in[1521];
     assign  data_out[3879] = data_in[1159];
     assign  data_out[3880] = data_in[1300];
     assign  data_out[3881] = data_in[215];
     assign  data_out[3882] = data_in[1277];
     assign  data_out[3883] = data_in[810];
     assign  data_out[3884] = data_in[1308];
     assign  data_out[3885] = data_in[630];
     assign  data_out[3886] = data_in[1574];
     assign  data_out[3887] = data_in[519];
     assign  data_out[3888] = data_in[251];
     assign  data_out[3889] = data_in[1348];
     assign  data_out[3890] = data_in[416];
     assign  data_out[3891] = data_in[1104];
     assign  data_out[3892] = data_in[1681];
     assign  data_out[3893] = data_in[477];
     assign  data_out[3894] = data_in[497];
     assign  data_out[3895] = data_in[832];
     assign  data_out[3896] = data_in[1265];
     assign  data_out[3897] = data_in[736];
     assign  data_out[3898] = data_in[1171];
     assign  data_out[3899] = data_in[708];
     assign  data_out[3900] = data_in[1373];
     assign  data_out[3901] = data_in[468];
     assign  data_out[3902] = data_in[570];
     assign  data_out[3903] = data_in[75];
     assign  data_out[3904] = data_in[1161];
     assign  data_out[3905] = data_in[1129];
     assign  data_out[3906] = data_in[134];
     assign  data_out[3907] = data_in[510];
     assign  data_out[3908] = data_in[1531];
     assign  data_out[3909] = data_in[1280];
     assign  data_out[3910] = data_in[1257];
     assign  data_out[3911] = data_in[562];
     assign  data_out[3912] = data_in[1241];
     assign  data_out[3913] = data_in[1542];
     assign  data_out[3914] = data_in[131];
     assign  data_out[3915] = data_in[1057];
     assign  data_out[3916] = data_in[1090];
     assign  data_out[3917] = data_in[922];
     assign  data_out[3918] = data_in[1594];
     assign  data_out[3919] = data_in[66];
     assign  data_out[3920] = data_in[1089];
     assign  data_out[3921] = data_in[314];
     assign  data_out[3922] = data_in[1050];
     assign  data_out[3923] = data_in[694];
     assign  data_out[3924] = data_in[622];
     assign  data_out[3925] = data_in[500];
     assign  data_out[3926] = data_in[189];
     assign  data_out[3927] = data_in[441];
     assign  data_out[3928] = data_in[359];
     assign  data_out[3929] = data_in[107];
     assign  data_out[3930] = data_in[387];
     assign  data_out[3931] = data_in[837];
     assign  data_out[3932] = data_in[338];
     assign  data_out[3933] = data_in[1546];
     assign  data_out[3934] = data_in[1501];
     assign  data_out[3935] = data_in[907];
     assign  data_out[3936] = data_in[1644];
     assign  data_out[3937] = data_in[1035];
     assign  data_out[3938] = data_in[57];
     assign  data_out[3939] = data_in[1094];
     assign  data_out[3940] = data_in[908];
     assign  data_out[3941] = data_in[112];
     assign  data_out[3942] = data_in[718];
     assign  data_out[3943] = data_in[186];
     assign  data_out[3944] = data_in[602];
     assign  data_out[3945] = data_in[903];
     assign  data_out[3946] = data_in[461];
     assign  data_out[3947] = data_in[1512];
     assign  data_out[3948] = data_in[173];
     assign  data_out[3949] = data_in[89];
     assign  data_out[3950] = data_in[834];
     assign  data_out[3951] = data_in[590];
     assign  data_out[3952] = data_in[1349];
     assign  data_out[3953] = data_in[866];
     assign  data_out[3954] = data_in[815];
     assign  data_out[3955] = data_in[1585];
     assign  data_out[3956] = data_in[1306];
     assign  data_out[3957] = data_in[821];
     assign  data_out[3958] = data_in[1424];
     assign  data_out[3959] = data_in[219];
     assign  data_out[3960] = data_in[110];
     assign  data_out[3961] = data_in[924];
     assign  data_out[3962] = data_in[564];
     assign  data_out[3963] = data_in[1205];
     assign  data_out[3964] = data_in[1317];
     assign  data_out[3965] = data_in[486];
     assign  data_out[3966] = data_in[588];
     assign  data_out[3967] = data_in[941];
     assign  data_out[3968] = data_in[1040];
     assign  data_out[3969] = data_in[815];
     assign  data_out[3970] = data_in[142];
     assign  data_out[3971] = data_in[101];
     assign  data_out[3972] = data_in[1373];
     assign  data_out[3973] = data_in[1421];
     assign  data_out[3974] = data_in[1446];
     assign  data_out[3975] = data_in[1020];
     assign  data_out[3976] = data_in[307];
     assign  data_out[3977] = data_in[1137];
     assign  data_out[3978] = data_in[1088];
     assign  data_out[3979] = data_in[955];
     assign  data_out[3980] = data_in[919];
     assign  data_out[3981] = data_in[114];
     assign  data_out[3982] = data_in[691];
     assign  data_out[3983] = data_in[67];
     assign  data_out[3984] = data_in[621];
     assign  data_out[3985] = data_in[1216];
     assign  data_out[3986] = data_in[329];
     assign  data_out[3987] = data_in[628];
     assign  data_out[3988] = data_in[1519];
     assign  data_out[3989] = data_in[1599];
     assign  data_out[3990] = data_in[694];
     assign  data_out[3991] = data_in[749];
     assign  data_out[3992] = data_in[931];
     assign  data_out[3993] = data_in[652];
     assign  data_out[3994] = data_in[1091];
     assign  data_out[3995] = data_in[619];
     assign  data_out[3996] = data_in[1409];
     assign  data_out[3997] = data_in[1241];
     assign  data_out[3998] = data_in[225];
     assign  data_out[3999] = data_in[342];
     assign  data_out[4000] = data_in[1016];
     assign  data_out[4001] = data_in[1084];
     assign  data_out[4002] = data_in[710];
     assign  data_out[4003] = data_in[457];
     assign  data_out[4004] = data_in[1496];
     assign  data_out[4005] = data_in[1290];
     assign  data_out[4006] = data_in[70];
     assign  data_out[4007] = data_in[1513];
     assign  data_out[4008] = data_in[255];
     assign  data_out[4009] = data_in[1252];
     assign  data_out[4010] = data_in[243];
     assign  data_out[4011] = data_in[1676];
     assign  data_out[4012] = data_in[346];
     assign  data_out[4013] = data_in[10];
     assign  data_out[4014] = data_in[1099];
     assign  data_out[4015] = data_in[849];
     assign  data_out[4016] = data_in[923];
     assign  data_out[4017] = data_in[922];
     assign  data_out[4018] = data_in[1343];
     assign  data_out[4019] = data_in[1637];
     assign  data_out[4020] = data_in[614];
     assign  data_out[4021] = data_in[26];
     assign  data_out[4022] = data_in[1677];
     assign  data_out[4023] = data_in[75];
     assign  data_out[4024] = data_in[481];
     assign  data_out[4025] = data_in[1566];
     assign  data_out[4026] = data_in[765];
     assign  data_out[4027] = data_in[1396];
     assign  data_out[4028] = data_in[1005];
     assign  data_out[4029] = data_in[1341];
     assign  data_out[4030] = data_in[1347];
     assign  data_out[4031] = data_in[191];
     assign  data_out[4032] = data_in[488];
     assign  data_out[4033] = data_in[347];
     assign  data_out[4034] = data_in[1489];
     assign  data_out[4035] = data_in[1684];
     assign  data_out[4036] = data_in[1412];
     assign  data_out[4037] = data_in[1474];
     assign  data_out[4038] = data_in[401];
     assign  data_out[4039] = data_in[1032];
     assign  data_out[4040] = data_in[1048];
     assign  data_out[4041] = data_in[1604];
     assign  data_out[4042] = data_in[742];
     assign  data_out[4043] = data_in[835];
     assign  data_out[4044] = data_in[493];
     assign  data_out[4045] = data_in[1005];
     assign  data_out[4046] = data_in[536];
     assign  data_out[4047] = data_in[1022];
     assign  data_out[4048] = data_in[1520];
     assign  data_out[4049] = data_in[896];
     assign  data_out[4050] = data_in[1561];
     assign  data_out[4051] = data_in[1571];
     assign  data_out[4052] = data_in[1236];
     assign  data_out[4053] = data_in[690];
     assign  data_out[4054] = data_in[1405];
     assign  data_out[4055] = data_in[615];
     assign  data_out[4056] = data_in[575];
     assign  data_out[4057] = data_in[378];
     assign  data_out[4058] = data_in[1243];
     assign  data_out[4059] = data_in[724];
     assign  data_out[4060] = data_in[335];
     assign  data_out[4061] = data_in[527];
     assign  data_out[4062] = data_in[1704];
     assign  data_out[4063] = data_in[761];
     assign  data_out[4064] = data_in[797];
     assign  data_out[4065] = data_in[191];
     assign  data_out[4066] = data_in[1611];
     assign  data_out[4067] = data_in[1630];
     assign  data_out[4068] = data_in[1094];
     assign  data_out[4069] = data_in[755];
     assign  data_out[4070] = data_in[1337];
     assign  data_out[4071] = data_in[1591];
     assign  data_out[4072] = data_in[533];
     assign  data_out[4073] = data_in[442];
     assign  data_out[4074] = data_in[1355];
     assign  data_out[4075] = data_in[830];
     assign  data_out[4076] = data_in[1507];
     assign  data_out[4077] = data_in[1355];
     assign  data_out[4078] = data_in[1209];
     assign  data_out[4079] = data_in[1315];
     assign  data_out[4080] = data_in[650];
     assign  data_out[4081] = data_in[1667];
     assign  data_out[4082] = data_in[1546];
     assign  data_out[4083] = data_in[898];
     assign  data_out[4084] = data_in[687];
     assign  data_out[4085] = data_in[26];
     assign  data_out[4086] = data_in[639];
     assign  data_out[4087] = data_in[522];
     assign  data_out[4088] = data_in[276];
     assign  data_out[4089] = data_in[332];
     assign  data_out[4090] = data_in[131];
     assign  data_out[4091] = data_in[1028];
     assign  data_out[4092] = data_in[1195];
     assign  data_out[4093] = data_in[755];
     assign  data_out[4094] = data_in[1042];
     assign  data_out[4095] = data_in[1514];
     assign  data_out[4096] = data_in[535];
     assign  data_out[4097] = data_in[94];
     assign  data_out[4098] = data_in[1343];
     assign  data_out[4099] = data_in[1656];
     assign  data_out[4100] = data_in[354];
     assign  data_out[4101] = data_in[132];
     assign  data_out[4102] = data_in[315];
     assign  data_out[4103] = data_in[938];
     assign  data_out[4104] = data_in[715];
     assign  data_out[4105] = data_in[825];
     assign  data_out[4106] = data_in[257];
     assign  data_out[4107] = data_in[659];
     assign  data_out[4108] = data_in[1650];
     assign  data_out[4109] = data_in[1532];
     assign  data_out[4110] = data_in[405];
     assign  data_out[4111] = data_in[1650];
     assign  data_out[4112] = data_in[710];
     assign  data_out[4113] = data_in[1664];
     assign  data_out[4114] = data_in[1267];
     assign  data_out[4115] = data_in[140];
     assign  data_out[4116] = data_in[1289];
     assign  data_out[4117] = data_in[139];
     assign  data_out[4118] = data_in[409];
     assign  data_out[4119] = data_in[595];
     assign  data_out[4120] = data_in[1076];
     assign  data_out[4121] = data_in[840];
     assign  data_out[4122] = data_in[1357];
     assign  data_out[4123] = data_in[1332];
     assign  data_out[4124] = data_in[35];
     assign  data_out[4125] = data_in[1013];
     assign  data_out[4126] = data_in[1108];
     assign  data_out[4127] = data_in[1101];
     assign  data_out[4128] = data_in[720];
     assign  data_out[4129] = data_in[885];
     assign  data_out[4130] = data_in[359];
     assign  data_out[4131] = data_in[1445];
     assign  data_out[4132] = data_in[570];
     assign  data_out[4133] = data_in[1088];
     assign  data_out[4134] = data_in[228];
     assign  data_out[4135] = data_in[1195];
     assign  data_out[4136] = data_in[846];
     assign  data_out[4137] = data_in[245];
     assign  data_out[4138] = data_in[211];
     assign  data_out[4139] = data_in[1099];
     assign  data_out[4140] = data_in[744];
     assign  data_out[4141] = data_in[766];
     assign  data_out[4142] = data_in[871];
     assign  data_out[4143] = data_in[1139];
     assign  data_out[4144] = data_in[1343];
     assign  data_out[4145] = data_in[662];
     assign  data_out[4146] = data_in[102];
     assign  data_out[4147] = data_in[1600];
     assign  data_out[4148] = data_in[17];
     assign  data_out[4149] = data_in[163];
     assign  data_out[4150] = data_in[285];
     assign  data_out[4151] = data_in[823];
     assign  data_out[4152] = data_in[1713];
     assign  data_out[4153] = data_in[936];
     assign  data_out[4154] = data_in[1338];
     assign  data_out[4155] = data_in[712];
     assign  data_out[4156] = data_in[56];
     assign  data_out[4157] = data_in[771];
     assign  data_out[4158] = data_in[459];
     assign  data_out[4159] = data_in[822];
     assign  data_out[4160] = data_in[1347];
     assign  data_out[4161] = data_in[1286];
     assign  data_out[4162] = data_in[1193];
     assign  data_out[4163] = data_in[737];
     assign  data_out[4164] = data_in[1227];
     assign  data_out[4165] = data_in[409];
     assign  data_out[4166] = data_in[784];
     assign  data_out[4167] = data_in[216];
     assign  data_out[4168] = data_in[878];
     assign  data_out[4169] = data_in[1004];
     assign  data_out[4170] = data_in[1661];
     assign  data_out[4171] = data_in[1254];
     assign  data_out[4172] = data_in[181];
     assign  data_out[4173] = data_in[498];
     assign  data_out[4174] = data_in[436];
     assign  data_out[4175] = data_in[1538];
     assign  data_out[4176] = data_in[1165];
     assign  data_out[4177] = data_in[1514];
     assign  data_out[4178] = data_in[289];
     assign  data_out[4179] = data_in[724];
     assign  data_out[4180] = data_in[600];
     assign  data_out[4181] = data_in[1447];
     assign  data_out[4182] = data_in[111];
     assign  data_out[4183] = data_in[384];
     assign  data_out[4184] = data_in[1628];
     assign  data_out[4185] = data_in[1003];
     assign  data_out[4186] = data_in[1086];
     assign  data_out[4187] = data_in[29];
     assign  data_out[4188] = data_in[838];
     assign  data_out[4189] = data_in[1716];
     assign  data_out[4190] = data_in[1382];
     assign  data_out[4191] = data_in[1164];
     assign  data_out[4192] = data_in[1382];
     assign  data_out[4193] = data_in[1372];
     assign  data_out[4194] = data_in[602];
     assign  data_out[4195] = data_in[1053];
     assign  data_out[4196] = data_in[1653];
     assign  data_out[4197] = data_in[551];
     assign  data_out[4198] = data_in[231];
     assign  data_out[4199] = data_in[232];
     assign  data_out[4200] = data_in[1466];
     assign  data_out[4201] = data_in[1569];
     assign  data_out[4202] = data_in[998];
     assign  data_out[4203] = data_in[284];
     assign  data_out[4204] = data_in[1191];
     assign  data_out[4205] = data_in[932];
     assign  data_out[4206] = data_in[656];
     assign  data_out[4207] = data_in[338];
     assign  data_out[4208] = data_in[1223];
     assign  data_out[4209] = data_in[1513];
     assign  data_out[4210] = data_in[14];
     assign  data_out[4211] = data_in[1652];
     assign  data_out[4212] = data_in[1416];
     assign  data_out[4213] = data_in[642];
     assign  data_out[4214] = data_in[1725];
     assign  data_out[4215] = data_in[1102];
     assign  data_out[4216] = data_in[961];
     assign  data_out[4217] = data_in[1047];
     assign  data_out[4218] = data_in[1015];
     assign  data_out[4219] = data_in[195];
     assign  data_out[4220] = data_in[73];
     assign  data_out[4221] = data_in[837];
     assign  data_out[4222] = data_in[1248];
     assign  data_out[4223] = data_in[77];
     assign  data_out[4224] = data_in[497];
     assign  data_out[4225] = data_in[837];
     assign  data_out[4226] = data_in[1662];
     assign  data_out[4227] = data_in[510];
     assign  data_out[4228] = data_in[1010];
     assign  data_out[4229] = data_in[1000];
     assign  data_out[4230] = data_in[544];
     assign  data_out[4231] = data_in[934];
     assign  data_out[4232] = data_in[512];
     assign  data_out[4233] = data_in[27];
     assign  data_out[4234] = data_in[934];
     assign  data_out[4235] = data_in[856];
     assign  data_out[4236] = data_in[1384];
     assign  data_out[4237] = data_in[1025];
     assign  data_out[4238] = data_in[1630];
     assign  data_out[4239] = data_in[1133];
     assign  data_out[4240] = data_in[1538];
     assign  data_out[4241] = data_in[1028];
     assign  data_out[4242] = data_in[329];
     assign  data_out[4243] = data_in[1666];
     assign  data_out[4244] = data_in[685];
     assign  data_out[4245] = data_in[69];
     assign  data_out[4246] = data_in[325];
     assign  data_out[4247] = data_in[537];
     assign  data_out[4248] = data_in[559];
     assign  data_out[4249] = data_in[695];
     assign  data_out[4250] = data_in[948];
     assign  data_out[4251] = data_in[450];
     assign  data_out[4252] = data_in[477];
     assign  data_out[4253] = data_in[792];
     assign  data_out[4254] = data_in[1155];
     assign  data_out[4255] = data_in[1613];
     assign  data_out[4256] = data_in[789];
     assign  data_out[4257] = data_in[725];
     assign  data_out[4258] = data_in[1669];
     assign  data_out[4259] = data_in[739];
     assign  data_out[4260] = data_in[29];
     assign  data_out[4261] = data_in[1726];
     assign  data_out[4262] = data_in[511];
     assign  data_out[4263] = data_in[1205];
     assign  data_out[4264] = data_in[75];
     assign  data_out[4265] = data_in[1001];
     assign  data_out[4266] = data_in[130];
     assign  data_out[4267] = data_in[509];
     assign  data_out[4268] = data_in[1664];
     assign  data_out[4269] = data_in[223];
     assign  data_out[4270] = data_in[271];
     assign  data_out[4271] = data_in[1521];
     assign  data_out[4272] = data_in[1105];
     assign  data_out[4273] = data_in[52];
     assign  data_out[4274] = data_in[1689];
     assign  data_out[4275] = data_in[1558];
     assign  data_out[4276] = data_in[1646];
     assign  data_out[4277] = data_in[806];
     assign  data_out[4278] = data_in[20];
     assign  data_out[4279] = data_in[620];
     assign  data_out[4280] = data_in[238];
     assign  data_out[4281] = data_in[924];
     assign  data_out[4282] = data_in[110];
     assign  data_out[4283] = data_in[87];
     assign  data_out[4284] = data_in[1144];
     assign  data_out[4285] = data_in[1269];
     assign  data_out[4286] = data_in[740];
     assign  data_out[4287] = data_in[375];
     assign  data_out[4288] = data_in[1605];
     assign  data_out[4289] = data_in[1705];
     assign  data_out[4290] = data_in[784];
     assign  data_out[4291] = data_in[1694];
     assign  data_out[4292] = data_in[1003];
     assign  data_out[4293] = data_in[1461];
     assign  data_out[4294] = data_in[920];
     assign  data_out[4295] = data_in[842];
     assign  data_out[4296] = data_in[1188];
     assign  data_out[4297] = data_in[96];
     assign  data_out[4298] = data_in[106];
     assign  data_out[4299] = data_in[292];
     assign  data_out[4300] = data_in[1047];
     assign  data_out[4301] = data_in[186];
     assign  data_out[4302] = data_in[671];
     assign  data_out[4303] = data_in[20];
     assign  data_out[4304] = data_in[1347];
     assign  data_out[4305] = data_in[1655];
     assign  data_out[4306] = data_in[501];
     assign  data_out[4307] = data_in[446];
     assign  data_out[4308] = data_in[467];
     assign  data_out[4309] = data_in[962];
     assign  data_out[4310] = data_in[4];
     assign  data_out[4311] = data_in[747];
     assign  data_out[4312] = data_in[519];
     assign  data_out[4313] = data_in[607];
     assign  data_out[4314] = data_in[593];
     assign  data_out[4315] = data_in[182];
     assign  data_out[4316] = data_in[1009];
     assign  data_out[4317] = data_in[714];
     assign  data_out[4318] = data_in[1643];
     assign  data_out[4319] = data_in[523];
     assign  data_out[4320] = data_in[1266];
     assign  data_out[4321] = data_in[608];
     assign  data_out[4322] = data_in[298];
     assign  data_out[4323] = data_in[1656];
     assign  data_out[4324] = data_in[883];
     assign  data_out[4325] = data_in[1147];
     assign  data_out[4326] = data_in[1100];
     assign  data_out[4327] = data_in[565];
     assign  data_out[4328] = data_in[402];
     assign  data_out[4329] = data_in[1178];
     assign  data_out[4330] = data_in[65];
     assign  data_out[4331] = data_in[1305];
     assign  data_out[4332] = data_in[115];
     assign  data_out[4333] = data_in[1330];
     assign  data_out[4334] = data_in[284];
     assign  data_out[4335] = data_in[1250];
     assign  data_out[4336] = data_in[936];
     assign  data_out[4337] = data_in[1617];
     assign  data_out[4338] = data_in[1215];
     assign  data_out[4339] = data_in[958];
     assign  data_out[4340] = data_in[63];
     assign  data_out[4341] = data_in[860];
     assign  data_out[4342] = data_in[1467];
     assign  data_out[4343] = data_in[1230];
     assign  data_out[4344] = data_in[896];
     assign  data_out[4345] = data_in[1692];
     assign  data_out[4346] = data_in[436];
     assign  data_out[4347] = data_in[136];
     assign  data_out[4348] = data_in[571];
     assign  data_out[4349] = data_in[1515];
     assign  data_out[4350] = data_in[585];
     assign  data_out[4351] = data_in[222];
     assign  data_out[4352] = data_in[519];
     assign  data_out[4353] = data_in[802];
     assign  data_out[4354] = data_in[910];
     assign  data_out[4355] = data_in[687];
     assign  data_out[4356] = data_in[1641];
     assign  data_out[4357] = data_in[487];
     assign  data_out[4358] = data_in[648];
     assign  data_out[4359] = data_in[280];
     assign  data_out[4360] = data_in[155];
     assign  data_out[4361] = data_in[823];
     assign  data_out[4362] = data_in[341];
     assign  data_out[4363] = data_in[1251];
     assign  data_out[4364] = data_in[1012];
     assign  data_out[4365] = data_in[1103];
     assign  data_out[4366] = data_in[289];
     assign  data_out[4367] = data_in[378];
     assign  data_out[4368] = data_in[973];
     assign  data_out[4369] = data_in[523];
     assign  data_out[4370] = data_in[780];
     assign  data_out[4371] = data_in[590];
     assign  data_out[4372] = data_in[1462];
     assign  data_out[4373] = data_in[1309];
     assign  data_out[4374] = data_in[687];
     assign  data_out[4375] = data_in[1572];
     assign  data_out[4376] = data_in[1565];
     assign  data_out[4377] = data_in[567];
     assign  data_out[4378] = data_in[539];
     assign  data_out[4379] = data_in[1132];
     assign  data_out[4380] = data_in[169];
     assign  data_out[4381] = data_in[1363];
     assign  data_out[4382] = data_in[1473];
     assign  data_out[4383] = data_in[285];
     assign  data_out[4384] = data_in[817];
     assign  data_out[4385] = data_in[92];
     assign  data_out[4386] = data_in[998];
     assign  data_out[4387] = data_in[633];
     assign  data_out[4388] = data_in[1629];
     assign  data_out[4389] = data_in[1396];
     assign  data_out[4390] = data_in[1162];
     assign  data_out[4391] = data_in[813];
     assign  data_out[4392] = data_in[130];
     assign  data_out[4393] = data_in[414];
     assign  data_out[4394] = data_in[673];
     assign  data_out[4395] = data_in[1339];
     assign  data_out[4396] = data_in[542];
     assign  data_out[4397] = data_in[895];
     assign  data_out[4398] = data_in[404];
     assign  data_out[4399] = data_in[404];
     assign  data_out[4400] = data_in[1532];
     assign  data_out[4401] = data_in[310];
     assign  data_out[4402] = data_in[730];
     assign  data_out[4403] = data_in[352];
     assign  data_out[4404] = data_in[343];
     assign  data_out[4405] = data_in[146];
     assign  data_out[4406] = data_in[1126];
     assign  data_out[4407] = data_in[465];
     assign  data_out[4408] = data_in[1697];
     assign  data_out[4409] = data_in[154];
     assign  data_out[4410] = data_in[1211];
     assign  data_out[4411] = data_in[952];
     assign  data_out[4412] = data_in[1706];
     assign  data_out[4413] = data_in[162];
     assign  data_out[4414] = data_in[1570];
     assign  data_out[4415] = data_in[714];
     assign  data_out[4416] = data_in[859];
     assign  data_out[4417] = data_in[1089];
     assign  data_out[4418] = data_in[73];
     assign  data_out[4419] = data_in[1665];
     assign  data_out[4420] = data_in[766];
     assign  data_out[4421] = data_in[1092];
     assign  data_out[4422] = data_in[1053];
     assign  data_out[4423] = data_in[453];
     assign  data_out[4424] = data_in[711];
     assign  data_out[4425] = data_in[956];
     assign  data_out[4426] = data_in[210];
     assign  data_out[4427] = data_in[1106];
     assign  data_out[4428] = data_in[526];
     assign  data_out[4429] = data_in[851];
     assign  data_out[4430] = data_in[621];
     assign  data_out[4431] = data_in[61];
     assign  data_out[4432] = data_in[1661];
     assign  data_out[4433] = data_in[807];
     assign  data_out[4434] = data_in[279];
     assign  data_out[4435] = data_in[1306];
     assign  data_out[4436] = data_in[865];
     assign  data_out[4437] = data_in[882];
     assign  data_out[4438] = data_in[1327];
     assign  data_out[4439] = data_in[976];
     assign  data_out[4440] = data_in[1163];
     assign  data_out[4441] = data_in[1268];
     assign  data_out[4442] = data_in[438];
     assign  data_out[4443] = data_in[887];
     assign  data_out[4444] = data_in[12];
     assign  data_out[4445] = data_in[31];
     assign  data_out[4446] = data_in[136];
     assign  data_out[4447] = data_in[700];
     assign  data_out[4448] = data_in[42];
     assign  data_out[4449] = data_in[842];
     assign  data_out[4450] = data_in[508];
     assign  data_out[4451] = data_in[550];
     assign  data_out[4452] = data_in[540];
     assign  data_out[4453] = data_in[734];
     assign  data_out[4454] = data_in[729];
     assign  data_out[4455] = data_in[131];
     assign  data_out[4456] = data_in[1258];
     assign  data_out[4457] = data_in[1347];
     assign  data_out[4458] = data_in[958];
     assign  data_out[4459] = data_in[141];
     assign  data_out[4460] = data_in[897];
     assign  data_out[4461] = data_in[1606];
     assign  data_out[4462] = data_in[1200];
     assign  data_out[4463] = data_in[729];
     assign  data_out[4464] = data_in[1112];
     assign  data_out[4465] = data_in[1467];
     assign  data_out[4466] = data_in[1504];
     assign  data_out[4467] = data_in[1110];
     assign  data_out[4468] = data_in[113];
     assign  data_out[4469] = data_in[599];
     assign  data_out[4470] = data_in[108];
     assign  data_out[4471] = data_in[177];
     assign  data_out[4472] = data_in[538];
     assign  data_out[4473] = data_in[890];
     assign  data_out[4474] = data_in[795];
     assign  data_out[4475] = data_in[554];
     assign  data_out[4476] = data_in[123];
     assign  data_out[4477] = data_in[116];
     assign  data_out[4478] = data_in[160];
     assign  data_out[4479] = data_in[355];
     assign  data_out[4480] = data_in[198];
     assign  data_out[4481] = data_in[1206];
     assign  data_out[4482] = data_in[626];
     assign  data_out[4483] = data_in[1026];
     assign  data_out[4484] = data_in[544];
     assign  data_out[4485] = data_in[241];
     assign  data_out[4486] = data_in[870];
     assign  data_out[4487] = data_in[1701];
     assign  data_out[4488] = data_in[104];
     assign  data_out[4489] = data_in[108];
     assign  data_out[4490] = data_in[878];
     assign  data_out[4491] = data_in[1546];
     assign  data_out[4492] = data_in[1427];
     assign  data_out[4493] = data_in[823];
     assign  data_out[4494] = data_in[943];
     assign  data_out[4495] = data_in[1248];
     assign  data_out[4496] = data_in[337];
     assign  data_out[4497] = data_in[1364];
     assign  data_out[4498] = data_in[703];
     assign  data_out[4499] = data_in[935];
     assign  data_out[4500] = data_in[192];
     assign  data_out[4501] = data_in[321];
     assign  data_out[4502] = data_in[10];
     assign  data_out[4503] = data_in[1244];
     assign  data_out[4504] = data_in[1099];
     assign  data_out[4505] = data_in[808];
     assign  data_out[4506] = data_in[806];
     assign  data_out[4507] = data_in[1353];
     assign  data_out[4508] = data_in[2];
     assign  data_out[4509] = data_in[53];
     assign  data_out[4510] = data_in[1442];
     assign  data_out[4511] = data_in[707];
     assign  data_out[4512] = data_in[401];
     assign  data_out[4513] = data_in[201];
     assign  data_out[4514] = data_in[1612];
     assign  data_out[4515] = data_in[1695];
     assign  data_out[4516] = data_in[212];
     assign  data_out[4517] = data_in[16];
     assign  data_out[4518] = data_in[696];
     assign  data_out[4519] = data_in[1020];
     assign  data_out[4520] = data_in[1469];
     assign  data_out[4521] = data_in[564];
     assign  data_out[4522] = data_in[789];
     assign  data_out[4523] = data_in[1562];
     assign  data_out[4524] = data_in[1724];
     assign  data_out[4525] = data_in[106];
     assign  data_out[4526] = data_in[650];
     assign  data_out[4527] = data_in[1378];
     assign  data_out[4528] = data_in[491];
     assign  data_out[4529] = data_in[921];
     assign  data_out[4530] = data_in[492];
     assign  data_out[4531] = data_in[277];
     assign  data_out[4532] = data_in[1319];
     assign  data_out[4533] = data_in[1559];
     assign  data_out[4534] = data_in[388];
     assign  data_out[4535] = data_in[1356];
     assign  data_out[4536] = data_in[1366];
     assign  data_out[4537] = data_in[704];
     assign  data_out[4538] = data_in[133];
     assign  data_out[4539] = data_in[1281];
     assign  data_out[4540] = data_in[903];
     assign  data_out[4541] = data_in[1690];
     assign  data_out[4542] = data_in[599];
     assign  data_out[4543] = data_in[244];
     assign  data_out[4544] = data_in[429];
     assign  data_out[4545] = data_in[655];
     assign  data_out[4546] = data_in[601];
     assign  data_out[4547] = data_in[1217];
     assign  data_out[4548] = data_in[544];
     assign  data_out[4549] = data_in[949];
     assign  data_out[4550] = data_in[1425];
     assign  data_out[4551] = data_in[47];
     assign  data_out[4552] = data_in[1633];
     assign  data_out[4553] = data_in[481];
     assign  data_out[4554] = data_in[918];
     assign  data_out[4555] = data_in[1671];
     assign  data_out[4556] = data_in[1235];
     assign  data_out[4557] = data_in[1548];
     assign  data_out[4558] = data_in[1392];
     assign  data_out[4559] = data_in[67];
     assign  data_out[4560] = data_in[1702];
     assign  data_out[4561] = data_in[185];
     assign  data_out[4562] = data_in[1164];
     assign  data_out[4563] = data_in[413];
     assign  data_out[4564] = data_in[93];
     assign  data_out[4565] = data_in[1126];
     assign  data_out[4566] = data_in[869];
     assign  data_out[4567] = data_in[341];
     assign  data_out[4568] = data_in[564];
     assign  data_out[4569] = data_in[1609];
     assign  data_out[4570] = data_in[1296];
     assign  data_out[4571] = data_in[118];
     assign  data_out[4572] = data_in[466];
     assign  data_out[4573] = data_in[449];
     assign  data_out[4574] = data_in[1426];
     assign  data_out[4575] = data_in[104];
     assign  data_out[4576] = data_in[763];
     assign  data_out[4577] = data_in[1561];
     assign  data_out[4578] = data_in[1046];
     assign  data_out[4579] = data_in[32];
     assign  data_out[4580] = data_in[650];
     assign  data_out[4581] = data_in[959];
     assign  data_out[4582] = data_in[1091];
     assign  data_out[4583] = data_in[1660];
     assign  data_out[4584] = data_in[1035];
     assign  data_out[4585] = data_in[701];
     assign  data_out[4586] = data_in[897];
     assign  data_out[4587] = data_in[1678];
     assign  data_out[4588] = data_in[974];
     assign  data_out[4589] = data_in[813];
     assign  data_out[4590] = data_in[1054];
     assign  data_out[4591] = data_in[639];
     assign  data_out[4592] = data_in[1345];
     assign  data_out[4593] = data_in[551];
     assign  data_out[4594] = data_in[692];
     assign  data_out[4595] = data_in[948];
     assign  data_out[4596] = data_in[1590];
     assign  data_out[4597] = data_in[1505];
     assign  data_out[4598] = data_in[1348];
     assign  data_out[4599] = data_in[671];
     assign  data_out[4600] = data_in[348];
     assign  data_out[4601] = data_in[720];
     assign  data_out[4602] = data_in[1040];
     assign  data_out[4603] = data_in[1152];
     assign  data_out[4604] = data_in[1349];
     assign  data_out[4605] = data_in[879];
     assign  data_out[4606] = data_in[1080];
     assign  data_out[4607] = data_in[613];
     assign  data_out[4608] = data_in[855];
     assign  data_out[4609] = data_in[1534];
     assign  data_out[4610] = data_in[622];
     assign  data_out[4611] = data_in[365];
     assign  data_out[4612] = data_in[1203];
     assign  data_out[4613] = data_in[181];
     assign  data_out[4614] = data_in[1453];
     assign  data_out[4615] = data_in[1014];
     assign  data_out[4616] = data_in[818];
     assign  data_out[4617] = data_in[1689];
     assign  data_out[4618] = data_in[1494];
     assign  data_out[4619] = data_in[1444];
     assign  data_out[4620] = data_in[62];
     assign  data_out[4621] = data_in[965];
     assign  data_out[4622] = data_in[1244];
     assign  data_out[4623] = data_in[423];
     assign  data_out[4624] = data_in[953];
     assign  data_out[4625] = data_in[1310];
     assign  data_out[4626] = data_in[1638];
     assign  data_out[4627] = data_in[1539];
     assign  data_out[4628] = data_in[357];
     assign  data_out[4629] = data_in[481];
     assign  data_out[4630] = data_in[263];
     assign  data_out[4631] = data_in[552];
     assign  data_out[4632] = data_in[1346];
     assign  data_out[4633] = data_in[42];
     assign  data_out[4634] = data_in[696];
     assign  data_out[4635] = data_in[816];
     assign  data_out[4636] = data_in[867];
     assign  data_out[4637] = data_in[1100];
     assign  data_out[4638] = data_in[441];
     assign  data_out[4639] = data_in[1286];
     assign  data_out[4640] = data_in[862];
     assign  data_out[4641] = data_in[539];
     assign  data_out[4642] = data_in[1594];
     assign  data_out[4643] = data_in[1034];
     assign  data_out[4644] = data_in[991];
     assign  data_out[4645] = data_in[961];
     assign  data_out[4646] = data_in[1083];
     assign  data_out[4647] = data_in[1095];
     assign  data_out[4648] = data_in[1095];
     assign  data_out[4649] = data_in[74];
     assign  data_out[4650] = data_in[1152];
     assign  data_out[4651] = data_in[883];
     assign  data_out[4652] = data_in[918];
     assign  data_out[4653] = data_in[369];
     assign  data_out[4654] = data_in[388];
     assign  data_out[4655] = data_in[1122];
     assign  data_out[4656] = data_in[1033];
     assign  data_out[4657] = data_in[1373];
     assign  data_out[4658] = data_in[786];
     assign  data_out[4659] = data_in[170];
     assign  data_out[4660] = data_in[1146];
     assign  data_out[4661] = data_in[1507];
     assign  data_out[4662] = data_in[1507];
     assign  data_out[4663] = data_in[838];
     assign  data_out[4664] = data_in[1432];
     assign  data_out[4665] = data_in[1198];
     assign  data_out[4666] = data_in[1006];
     assign  data_out[4667] = data_in[778];
     assign  data_out[4668] = data_in[1356];
     assign  data_out[4669] = data_in[1451];
     assign  data_out[4670] = data_in[662];
     assign  data_out[4671] = data_in[830];
     assign  data_out[4672] = data_in[1640];
     assign  data_out[4673] = data_in[1618];
     assign  data_out[4674] = data_in[449];
     assign  data_out[4675] = data_in[917];
     assign  data_out[4676] = data_in[364];
     assign  data_out[4677] = data_in[951];
     assign  data_out[4678] = data_in[552];
     assign  data_out[4679] = data_in[624];
     assign  data_out[4680] = data_in[957];
     assign  data_out[4681] = data_in[750];
     assign  data_out[4682] = data_in[1178];
     assign  data_out[4683] = data_in[1691];
     assign  data_out[4684] = data_in[611];
     assign  data_out[4685] = data_in[1332];
     assign  data_out[4686] = data_in[637];
     assign  data_out[4687] = data_in[173];
     assign  data_out[4688] = data_in[1065];
     assign  data_out[4689] = data_in[1002];
     assign  data_out[4690] = data_in[1238];
     assign  data_out[4691] = data_in[63];
     assign  data_out[4692] = data_in[1635];
     assign  data_out[4693] = data_in[1613];
     assign  data_out[4694] = data_in[600];
     assign  data_out[4695] = data_in[1570];
     assign  data_out[4696] = data_in[909];
     assign  data_out[4697] = data_in[254];
     assign  data_out[4698] = data_in[387];
     assign  data_out[4699] = data_in[1034];
     assign  data_out[4700] = data_in[1533];
     assign  data_out[4701] = data_in[1025];
     assign  data_out[4702] = data_in[1434];
     assign  data_out[4703] = data_in[597];
     assign  data_out[4704] = data_in[1295];
     assign  data_out[4705] = data_in[525];
     assign  data_out[4706] = data_in[1720];
     assign  data_out[4707] = data_in[668];
     assign  data_out[4708] = data_in[1240];
     assign  data_out[4709] = data_in[13];
     assign  data_out[4710] = data_in[700];
     assign  data_out[4711] = data_in[964];
     assign  data_out[4712] = data_in[194];
     assign  data_out[4713] = data_in[1318];
     assign  data_out[4714] = data_in[557];
     assign  data_out[4715] = data_in[435];
     assign  data_out[4716] = data_in[1235];
     assign  data_out[4717] = data_in[1464];
     assign  data_out[4718] = data_in[953];
     assign  data_out[4719] = data_in[1116];
     assign  data_out[4720] = data_in[1231];
     assign  data_out[4721] = data_in[82];
     assign  data_out[4722] = data_in[318];
     assign  data_out[4723] = data_in[1039];
     assign  data_out[4724] = data_in[1068];
     assign  data_out[4725] = data_in[42];
     assign  data_out[4726] = data_in[246];
     assign  data_out[4727] = data_in[254];
     assign  data_out[4728] = data_in[785];
     assign  data_out[4729] = data_in[1534];
     assign  data_out[4730] = data_in[117];
     assign  data_out[4731] = data_in[1634];
     assign  data_out[4732] = data_in[1683];
     assign  data_out[4733] = data_in[1130];
     assign  data_out[4734] = data_in[995];
     assign  data_out[4735] = data_in[1128];
     assign  data_out[4736] = data_in[358];
     assign  data_out[4737] = data_in[1275];
     assign  data_out[4738] = data_in[707];
     assign  data_out[4739] = data_in[999];
     assign  data_out[4740] = data_in[190];
     assign  data_out[4741] = data_in[225];
     assign  data_out[4742] = data_in[912];
     assign  data_out[4743] = data_in[945];
     assign  data_out[4744] = data_in[1027];
     assign  data_out[4745] = data_in[733];
     assign  data_out[4746] = data_in[1135];
     assign  data_out[4747] = data_in[648];
     assign  data_out[4748] = data_in[1265];
     assign  data_out[4749] = data_in[587];
     assign  data_out[4750] = data_in[572];
     assign  data_out[4751] = data_in[1494];
     assign  data_out[4752] = data_in[689];
     assign  data_out[4753] = data_in[1575];
     assign  data_out[4754] = data_in[1668];
     assign  data_out[4755] = data_in[1241];
     assign  data_out[4756] = data_in[257];
     assign  data_out[4757] = data_in[1707];
     assign  data_out[4758] = data_in[1692];
     assign  data_out[4759] = data_in[495];
     assign  data_out[4760] = data_in[1039];
     assign  data_out[4761] = data_in[345];
     assign  data_out[4762] = data_in[884];
     assign  data_out[4763] = data_in[952];
     assign  data_out[4764] = data_in[199];
     assign  data_out[4765] = data_in[104];
     assign  data_out[4766] = data_in[1304];
     assign  data_out[4767] = data_in[429];
     assign  data_out[4768] = data_in[67];
     assign  data_out[4769] = data_in[592];
     assign  data_out[4770] = data_in[754];
     assign  data_out[4771] = data_in[948];
     assign  data_out[4772] = data_in[535];
     assign  data_out[4773] = data_in[695];
     assign  data_out[4774] = data_in[839];
     assign  data_out[4775] = data_in[311];
     assign  data_out[4776] = data_in[1196];
     assign  data_out[4777] = data_in[1022];
     assign  data_out[4778] = data_in[708];
     assign  data_out[4779] = data_in[731];
     assign  data_out[4780] = data_in[742];
     assign  data_out[4781] = data_in[738];
     assign  data_out[4782] = data_in[726];
     assign  data_out[4783] = data_in[1500];
     assign  data_out[4784] = data_in[1025];
     assign  data_out[4785] = data_in[1152];
     assign  data_out[4786] = data_in[1424];
     assign  data_out[4787] = data_in[600];
     assign  data_out[4788] = data_in[1577];
     assign  data_out[4789] = data_in[1637];
     assign  data_out[4790] = data_in[1268];
     assign  data_out[4791] = data_in[1636];
     assign  data_out[4792] = data_in[625];
     assign  data_out[4793] = data_in[259];
     assign  data_out[4794] = data_in[1050];
     assign  data_out[4795] = data_in[874];
     assign  data_out[4796] = data_in[498];
     assign  data_out[4797] = data_in[228];
     assign  data_out[4798] = data_in[1138];
     assign  data_out[4799] = data_in[877];
     assign  data_out[4800] = data_in[631];
     assign  data_out[4801] = data_in[8];
     assign  data_out[4802] = data_in[1156];
     assign  data_out[4803] = data_in[1332];
     assign  data_out[4804] = data_in[252];
     assign  data_out[4805] = data_in[1017];
     assign  data_out[4806] = data_in[404];
     assign  data_out[4807] = data_in[1454];
     assign  data_out[4808] = data_in[870];
     assign  data_out[4809] = data_in[385];
     assign  data_out[4810] = data_in[1665];
     assign  data_out[4811] = data_in[869];
     assign  data_out[4812] = data_in[1272];
     assign  data_out[4813] = data_in[986];
     assign  data_out[4814] = data_in[1188];
     assign  data_out[4815] = data_in[514];
     assign  data_out[4816] = data_in[1072];
     assign  data_out[4817] = data_in[1019];
     assign  data_out[4818] = data_in[312];
     assign  data_out[4819] = data_in[824];
     assign  data_out[4820] = data_in[332];
     assign  data_out[4821] = data_in[535];
     assign  data_out[4822] = data_in[762];
     assign  data_out[4823] = data_in[477];
     assign  data_out[4824] = data_in[928];
     assign  data_out[4825] = data_in[1009];
     assign  data_out[4826] = data_in[112];
     assign  data_out[4827] = data_in[1611];
     assign  data_out[4828] = data_in[649];
     assign  data_out[4829] = data_in[812];
     assign  data_out[4830] = data_in[1269];
     assign  data_out[4831] = data_in[585];
     assign  data_out[4832] = data_in[1233];
     assign  data_out[4833] = data_in[676];
     assign  data_out[4834] = data_in[615];
     assign  data_out[4835] = data_in[1296];
     assign  data_out[4836] = data_in[609];
     assign  data_out[4837] = data_in[1271];
     assign  data_out[4838] = data_in[1528];
     assign  data_out[4839] = data_in[772];
     assign  data_out[4840] = data_in[920];
     assign  data_out[4841] = data_in[94];
     assign  data_out[4842] = data_in[612];
     assign  data_out[4843] = data_in[1300];
     assign  data_out[4844] = data_in[845];
     assign  data_out[4845] = data_in[884];
     assign  data_out[4846] = data_in[277];
     assign  data_out[4847] = data_in[564];
     assign  data_out[4848] = data_in[365];
     assign  data_out[4849] = data_in[1277];
     assign  data_out[4850] = data_in[192];
     assign  data_out[4851] = data_in[221];
     assign  data_out[4852] = data_in[301];
     assign  data_out[4853] = data_in[1313];
     assign  data_out[4854] = data_in[500];
     assign  data_out[4855] = data_in[1653];
     assign  data_out[4856] = data_in[578];
     assign  data_out[4857] = data_in[225];
     assign  data_out[4858] = data_in[431];
     assign  data_out[4859] = data_in[1701];
     assign  data_out[4860] = data_in[288];
     assign  data_out[4861] = data_in[1653];
     assign  data_out[4862] = data_in[1013];
     assign  data_out[4863] = data_in[310];
     assign  data_out[4864] = data_in[31];
     assign  data_out[4865] = data_in[1642];
     assign  data_out[4866] = data_in[694];
     assign  data_out[4867] = data_in[41];
     assign  data_out[4868] = data_in[986];
     assign  data_out[4869] = data_in[293];
     assign  data_out[4870] = data_in[1218];
     assign  data_out[4871] = data_in[764];
     assign  data_out[4872] = data_in[1191];
     assign  data_out[4873] = data_in[1046];
     assign  data_out[4874] = data_in[476];
     assign  data_out[4875] = data_in[589];
     assign  data_out[4876] = data_in[743];
     assign  data_out[4877] = data_in[470];
     assign  data_out[4878] = data_in[33];
     assign  data_out[4879] = data_in[1139];
     assign  data_out[4880] = data_in[867];
     assign  data_out[4881] = data_in[1647];
     assign  data_out[4882] = data_in[603];
     assign  data_out[4883] = data_in[609];
     assign  data_out[4884] = data_in[1646];
     assign  data_out[4885] = data_in[463];
     assign  data_out[4886] = data_in[1081];
     assign  data_out[4887] = data_in[345];
     assign  data_out[4888] = data_in[635];
     assign  data_out[4889] = data_in[343];
     assign  data_out[4890] = data_in[316];
     assign  data_out[4891] = data_in[1464];
     assign  data_out[4892] = data_in[618];
     assign  data_out[4893] = data_in[1303];
     assign  data_out[4894] = data_in[1683];
     assign  data_out[4895] = data_in[0];
     assign  data_out[4896] = data_in[1069];
     assign  data_out[4897] = data_in[1576];
     assign  data_out[4898] = data_in[632];
     assign  data_out[4899] = data_in[273];
     assign  data_out[4900] = data_in[601];
     assign  data_out[4901] = data_in[865];
     assign  data_out[4902] = data_in[206];
     assign  data_out[4903] = data_in[1393];
     assign  data_out[4904] = data_in[503];
     assign  data_out[4905] = data_in[304];
     assign  data_out[4906] = data_in[134];
     assign  data_out[4907] = data_in[810];
     assign  data_out[4908] = data_in[360];
     assign  data_out[4909] = data_in[269];
     assign  data_out[4910] = data_in[1041];
     assign  data_out[4911] = data_in[918];
     assign  data_out[4912] = data_in[63];
     assign  data_out[4913] = data_in[1474];
     assign  data_out[4914] = data_in[487];
     assign  data_out[4915] = data_in[405];
     assign  data_out[4916] = data_in[913];
     assign  data_out[4917] = data_in[141];
     assign  data_out[4918] = data_in[1644];
     assign  data_out[4919] = data_in[1293];
     assign  data_out[4920] = data_in[1134];
     assign  data_out[4921] = data_in[1692];
     assign  data_out[4922] = data_in[939];
     assign  data_out[4923] = data_in[1271];
     assign  data_out[4924] = data_in[949];
     assign  data_out[4925] = data_in[533];
     assign  data_out[4926] = data_in[1406];
     assign  data_out[4927] = data_in[522];
     assign  data_out[4928] = data_in[452];
     assign  data_out[4929] = data_in[497];
     assign  data_out[4930] = data_in[807];
     assign  data_out[4931] = data_in[1301];
     assign  data_out[4932] = data_in[236];
     assign  data_out[4933] = data_in[1067];
     assign  data_out[4934] = data_in[1224];
     assign  data_out[4935] = data_in[81];
     assign  data_out[4936] = data_in[104];
     assign  data_out[4937] = data_in[1465];
     assign  data_out[4938] = data_in[1325];
     assign  data_out[4939] = data_in[635];
     assign  data_out[4940] = data_in[654];
     assign  data_out[4941] = data_in[1294];
     assign  data_out[4942] = data_in[699];
     assign  data_out[4943] = data_in[1226];
     assign  data_out[4944] = data_in[1320];
     assign  data_out[4945] = data_in[1451];
     assign  data_out[4946] = data_in[1653];
     assign  data_out[4947] = data_in[1533];
     assign  data_out[4948] = data_in[1396];
     assign  data_out[4949] = data_in[1265];
     assign  data_out[4950] = data_in[1599];
     assign  data_out[4951] = data_in[1518];
     assign  data_out[4952] = data_in[1081];
     assign  data_out[4953] = data_in[769];
     assign  data_out[4954] = data_in[1148];
     assign  data_out[4955] = data_in[1552];
     assign  data_out[4956] = data_in[433];
     assign  data_out[4957] = data_in[595];
     assign  data_out[4958] = data_in[309];
     assign  data_out[4959] = data_in[204];
     assign  data_out[4960] = data_in[172];
     assign  data_out[4961] = data_in[1501];
     assign  data_out[4962] = data_in[998];
     assign  data_out[4963] = data_in[757];
     assign  data_out[4964] = data_in[513];
     assign  data_out[4965] = data_in[1195];
     assign  data_out[4966] = data_in[361];
     assign  data_out[4967] = data_in[354];
     assign  data_out[4968] = data_in[218];
     assign  data_out[4969] = data_in[834];
     assign  data_out[4970] = data_in[9];
     assign  data_out[4971] = data_in[519];
     assign  data_out[4972] = data_in[694];
     assign  data_out[4973] = data_in[1585];
     assign  data_out[4974] = data_in[132];
     assign  data_out[4975] = data_in[849];
     assign  data_out[4976] = data_in[69];
     assign  data_out[4977] = data_in[166];
     assign  data_out[4978] = data_in[126];
     assign  data_out[4979] = data_in[790];
     assign  data_out[4980] = data_in[1043];
     assign  data_out[4981] = data_in[53];
     assign  data_out[4982] = data_in[626];
     assign  data_out[4983] = data_in[683];
     assign  data_out[4984] = data_in[188];
     assign  data_out[4985] = data_in[601];
     assign  data_out[4986] = data_in[928];
     assign  data_out[4987] = data_in[1058];
     assign  data_out[4988] = data_in[1512];
     assign  data_out[4989] = data_in[1502];
     assign  data_out[4990] = data_in[513];
     assign  data_out[4991] = data_in[20];
     assign  data_out[4992] = data_in[1196];
     assign  data_out[4993] = data_in[396];
     assign  data_out[4994] = data_in[392];
     assign  data_out[4995] = data_in[1512];
     assign  data_out[4996] = data_in[164];
     assign  data_out[4997] = data_in[304];
     assign  data_out[4998] = data_in[886];
     assign  data_out[4999] = data_in[1472];
     assign  data_out[5000] = data_in[41];
     assign  data_out[5001] = data_in[1253];
     assign  data_out[5002] = data_in[193];
     assign  data_out[5003] = data_in[970];
     assign  data_out[5004] = data_in[1115];
     assign  data_out[5005] = data_in[1397];
     assign  data_out[5006] = data_in[733];
     assign  data_out[5007] = data_in[1222];
     assign  data_out[5008] = data_in[1083];
     assign  data_out[5009] = data_in[1013];
     assign  data_out[5010] = data_in[1710];
     assign  data_out[5011] = data_in[210];
     assign  data_out[5012] = data_in[1096];
     assign  data_out[5013] = data_in[123];
     assign  data_out[5014] = data_in[403];
     assign  data_out[5015] = data_in[1099];
     assign  data_out[5016] = data_in[595];
     assign  data_out[5017] = data_in[385];
     assign  data_out[5018] = data_in[1396];
     assign  data_out[5019] = data_in[326];
     assign  data_out[5020] = data_in[1285];
     assign  data_out[5021] = data_in[297];
     assign  data_out[5022] = data_in[956];
     assign  data_out[5023] = data_in[134];
     assign  data_out[5024] = data_in[5];
     assign  data_out[5025] = data_in[1250];
     assign  data_out[5026] = data_in[1040];
     assign  data_out[5027] = data_in[1306];
     assign  data_out[5028] = data_in[1214];
     assign  data_out[5029] = data_in[1389];
     assign  data_out[5030] = data_in[1157];
     assign  data_out[5031] = data_in[157];
     assign  data_out[5032] = data_in[1202];
     assign  data_out[5033] = data_in[1727];
     assign  data_out[5034] = data_in[104];
     assign  data_out[5035] = data_in[822];
     assign  data_out[5036] = data_in[662];
     assign  data_out[5037] = data_in[1472];
     assign  data_out[5038] = data_in[712];
     assign  data_out[5039] = data_in[1239];
     assign  data_out[5040] = data_in[1196];
     assign  data_out[5041] = data_in[97];
     assign  data_out[5042] = data_in[1244];
     assign  data_out[5043] = data_in[152];
     assign  data_out[5044] = data_in[908];
     assign  data_out[5045] = data_in[393];
     assign  data_out[5046] = data_in[1149];
     assign  data_out[5047] = data_in[810];
     assign  data_out[5048] = data_in[1688];
     assign  data_out[5049] = data_in[667];
     assign  data_out[5050] = data_in[1348];
     assign  data_out[5051] = data_in[1673];
     assign  data_out[5052] = data_in[144];
     assign  data_out[5053] = data_in[1419];
     assign  data_out[5054] = data_in[846];
     assign  data_out[5055] = data_in[1628];
     assign  data_out[5056] = data_in[699];
     assign  data_out[5057] = data_in[843];
     assign  data_out[5058] = data_in[939];
     assign  data_out[5059] = data_in[1391];
     assign  data_out[5060] = data_in[342];
     assign  data_out[5061] = data_in[1019];
     assign  data_out[5062] = data_in[1528];
     assign  data_out[5063] = data_in[959];
     assign  data_out[5064] = data_in[845];
     assign  data_out[5065] = data_in[886];
     assign  data_out[5066] = data_in[835];
     assign  data_out[5067] = data_in[693];
     assign  data_out[5068] = data_in[1375];
     assign  data_out[5069] = data_in[1309];
     assign  data_out[5070] = data_in[275];
     assign  data_out[5071] = data_in[714];
     assign  data_out[5072] = data_in[1402];
     assign  data_out[5073] = data_in[55];
     assign  data_out[5074] = data_in[1615];
     assign  data_out[5075] = data_in[1031];
     assign  data_out[5076] = data_in[1398];
     assign  data_out[5077] = data_in[267];
     assign  data_out[5078] = data_in[1626];
     assign  data_out[5079] = data_in[507];
     assign  data_out[5080] = data_in[99];
     assign  data_out[5081] = data_in[1613];
     assign  data_out[5082] = data_in[713];
     assign  data_out[5083] = data_in[558];
     assign  data_out[5084] = data_in[47];
     assign  data_out[5085] = data_in[1155];
     assign  data_out[5086] = data_in[1388];
     assign  data_out[5087] = data_in[1318];
     assign  data_out[5088] = data_in[1164];
     assign  data_out[5089] = data_in[759];
     assign  data_out[5090] = data_in[951];
     assign  data_out[5091] = data_in[1344];
     assign  data_out[5092] = data_in[979];
     assign  data_out[5093] = data_in[1434];
     assign  data_out[5094] = data_in[897];
     assign  data_out[5095] = data_in[710];
     assign  data_out[5096] = data_in[273];
     assign  data_out[5097] = data_in[435];
     assign  data_out[5098] = data_in[1152];
     assign  data_out[5099] = data_in[1251];
     assign  data_out[5100] = data_in[1673];
     assign  data_out[5101] = data_in[894];
     assign  data_out[5102] = data_in[1625];
     assign  data_out[5103] = data_in[377];
     assign  data_out[5104] = data_in[1667];
     assign  data_out[5105] = data_in[1420];
     assign  data_out[5106] = data_in[1659];
     assign  data_out[5107] = data_in[1585];
     assign  data_out[5108] = data_in[1594];
     assign  data_out[5109] = data_in[1365];
     assign  data_out[5110] = data_in[866];
     assign  data_out[5111] = data_in[71];
     assign  data_out[5112] = data_in[74];
     assign  data_out[5113] = data_in[1285];
     assign  data_out[5114] = data_in[555];
     assign  data_out[5115] = data_in[1135];
     assign  data_out[5116] = data_in[1061];
     assign  data_out[5117] = data_in[1462];
     assign  data_out[5118] = data_in[601];
     assign  data_out[5119] = data_in[394];
     assign  data_out[5120] = data_in[1719];
     assign  data_out[5121] = data_in[478];
     assign  data_out[5122] = data_in[1342];
     assign  data_out[5123] = data_in[795];
     assign  data_out[5124] = data_in[1206];
     assign  data_out[5125] = data_in[176];
     assign  data_out[5126] = data_in[159];
     assign  data_out[5127] = data_in[611];
     assign  data_out[5128] = data_in[1492];
     assign  data_out[5129] = data_in[1703];
     assign  data_out[5130] = data_in[959];
     assign  data_out[5131] = data_in[1494];
     assign  data_out[5132] = data_in[1544];
     assign  data_out[5133] = data_in[696];
     assign  data_out[5134] = data_in[326];
     assign  data_out[5135] = data_in[149];
     assign  data_out[5136] = data_in[931];
     assign  data_out[5137] = data_in[888];
     assign  data_out[5138] = data_in[1345];
     assign  data_out[5139] = data_in[610];
     assign  data_out[5140] = data_in[361];
     assign  data_out[5141] = data_in[607];
     assign  data_out[5142] = data_in[1628];
     assign  data_out[5143] = data_in[301];
     assign  data_out[5144] = data_in[1377];
     assign  data_out[5145] = data_in[823];
     assign  data_out[5146] = data_in[1343];
     assign  data_out[5147] = data_in[699];
     assign  data_out[5148] = data_in[1365];
     assign  data_out[5149] = data_in[1324];
     assign  data_out[5150] = data_in[231];
     assign  data_out[5151] = data_in[965];
     assign  data_out[5152] = data_in[1655];
     assign  data_out[5153] = data_in[828];
     assign  data_out[5154] = data_in[59];
     assign  data_out[5155] = data_in[1158];
     assign  data_out[5156] = data_in[674];
     assign  data_out[5157] = data_in[458];
     assign  data_out[5158] = data_in[477];
     assign  data_out[5159] = data_in[1058];
     assign  data_out[5160] = data_in[296];
     assign  data_out[5161] = data_in[457];
     assign  data_out[5162] = data_in[1293];
     assign  data_out[5163] = data_in[472];
     assign  data_out[5164] = data_in[812];
     assign  data_out[5165] = data_in[1675];
     assign  data_out[5166] = data_in[848];
     assign  data_out[5167] = data_in[871];
     assign  data_out[5168] = data_in[565];
     assign  data_out[5169] = data_in[1693];
     assign  data_out[5170] = data_in[50];
     assign  data_out[5171] = data_in[409];
     assign  data_out[5172] = data_in[1590];
     assign  data_out[5173] = data_in[584];
     assign  data_out[5174] = data_in[26];
     assign  data_out[5175] = data_in[1184];
     assign  data_out[5176] = data_in[1019];
     assign  data_out[5177] = data_in[989];
     assign  data_out[5178] = data_in[1225];
     assign  data_out[5179] = data_in[55];
     assign  data_out[5180] = data_in[702];
     assign  data_out[5181] = data_in[215];
     assign  data_out[5182] = data_in[564];
     assign  data_out[5183] = data_in[872];
     assign  data_out[5184] = data_in[966];
     assign  data_out[5185] = data_in[533];
     assign  data_out[5186] = data_in[1363];
     assign  data_out[5187] = data_in[442];
     assign  data_out[5188] = data_in[598];
     assign  data_out[5189] = data_in[791];
     assign  data_out[5190] = data_in[1559];
     assign  data_out[5191] = data_in[1632];
     assign  data_out[5192] = data_in[95];
     assign  data_out[5193] = data_in[726];
     assign  data_out[5194] = data_in[868];
     assign  data_out[5195] = data_in[745];
     assign  data_out[5196] = data_in[870];
     assign  data_out[5197] = data_in[88];
     assign  data_out[5198] = data_in[1024];
     assign  data_out[5199] = data_in[842];
     assign  data_out[5200] = data_in[914];
     assign  data_out[5201] = data_in[1504];
     assign  data_out[5202] = data_in[11];
     assign  data_out[5203] = data_in[1611];
     assign  data_out[5204] = data_in[365];
     assign  data_out[5205] = data_in[916];
     assign  data_out[5206] = data_in[1086];
     assign  data_out[5207] = data_in[172];
     assign  data_out[5208] = data_in[168];
     assign  data_out[5209] = data_in[437];
     assign  data_out[5210] = data_in[1210];
     assign  data_out[5211] = data_in[63];
     assign  data_out[5212] = data_in[383];
     assign  data_out[5213] = data_in[1549];
     assign  data_out[5214] = data_in[431];
     assign  data_out[5215] = data_in[604];
     assign  data_out[5216] = data_in[347];
     assign  data_out[5217] = data_in[1394];
     assign  data_out[5218] = data_in[285];
     assign  data_out[5219] = data_in[169];
     assign  data_out[5220] = data_in[304];
     assign  data_out[5221] = data_in[178];
     assign  data_out[5222] = data_in[1653];
     assign  data_out[5223] = data_in[1110];
     assign  data_out[5224] = data_in[1545];
     assign  data_out[5225] = data_in[975];
     assign  data_out[5226] = data_in[1260];
     assign  data_out[5227] = data_in[1472];
     assign  data_out[5228] = data_in[1217];
     assign  data_out[5229] = data_in[1321];
     assign  data_out[5230] = data_in[680];
     assign  data_out[5231] = data_in[1010];
     assign  data_out[5232] = data_in[1297];
     assign  data_out[5233] = data_in[1070];
     assign  data_out[5234] = data_in[1145];
     assign  data_out[5235] = data_in[1445];
     assign  data_out[5236] = data_in[252];
     assign  data_out[5237] = data_in[1711];
     assign  data_out[5238] = data_in[1465];
     assign  data_out[5239] = data_in[817];
     assign  data_out[5240] = data_in[693];
     assign  data_out[5241] = data_in[901];
     assign  data_out[5242] = data_in[1715];
     assign  data_out[5243] = data_in[1635];
     assign  data_out[5244] = data_in[1555];
     assign  data_out[5245] = data_in[586];
     assign  data_out[5246] = data_in[658];
     assign  data_out[5247] = data_in[1566];
     assign  data_out[5248] = data_in[1197];
     assign  data_out[5249] = data_in[1376];
     assign  data_out[5250] = data_in[1626];
     assign  data_out[5251] = data_in[186];
     assign  data_out[5252] = data_in[683];
     assign  data_out[5253] = data_in[1558];
     assign  data_out[5254] = data_in[1007];
     assign  data_out[5255] = data_in[908];
     assign  data_out[5256] = data_in[818];
     assign  data_out[5257] = data_in[1021];
     assign  data_out[5258] = data_in[1724];
     assign  data_out[5259] = data_in[136];
     assign  data_out[5260] = data_in[1192];
     assign  data_out[5261] = data_in[878];
     assign  data_out[5262] = data_in[1644];
     assign  data_out[5263] = data_in[1512];
     assign  data_out[5264] = data_in[6];
     assign  data_out[5265] = data_in[759];
     assign  data_out[5266] = data_in[1046];
     assign  data_out[5267] = data_in[649];
     assign  data_out[5268] = data_in[1197];
     assign  data_out[5269] = data_in[105];
     assign  data_out[5270] = data_in[1543];
     assign  data_out[5271] = data_in[678];
     assign  data_out[5272] = data_in[1712];
     assign  data_out[5273] = data_in[280];
     assign  data_out[5274] = data_in[831];
     assign  data_out[5275] = data_in[557];
     assign  data_out[5276] = data_in[20];
     assign  data_out[5277] = data_in[1712];
     assign  data_out[5278] = data_in[614];
     assign  data_out[5279] = data_in[900];
     assign  data_out[5280] = data_in[430];
     assign  data_out[5281] = data_in[1527];
     assign  data_out[5282] = data_in[957];
     assign  data_out[5283] = data_in[394];
     assign  data_out[5284] = data_in[736];
     assign  data_out[5285] = data_in[1447];
     assign  data_out[5286] = data_in[138];
     assign  data_out[5287] = data_in[1638];
     assign  data_out[5288] = data_in[1701];
     assign  data_out[5289] = data_in[302];
     assign  data_out[5290] = data_in[920];
     assign  data_out[5291] = data_in[1189];
     assign  data_out[5292] = data_in[1701];
     assign  data_out[5293] = data_in[1659];
     assign  data_out[5294] = data_in[827];
     assign  data_out[5295] = data_in[1675];
     assign  data_out[5296] = data_in[1220];
     assign  data_out[5297] = data_in[565];
     assign  data_out[5298] = data_in[170];
     assign  data_out[5299] = data_in[14];
     assign  data_out[5300] = data_in[1256];
     assign  data_out[5301] = data_in[633];
     assign  data_out[5302] = data_in[246];
     assign  data_out[5303] = data_in[1687];
     assign  data_out[5304] = data_in[1314];
     assign  data_out[5305] = data_in[1281];
     assign  data_out[5306] = data_in[1244];
     assign  data_out[5307] = data_in[1303];
     assign  data_out[5308] = data_in[58];
     assign  data_out[5309] = data_in[1159];
     assign  data_out[5310] = data_in[1668];
     assign  data_out[5311] = data_in[118];
     assign  data_out[5312] = data_in[849];
     assign  data_out[5313] = data_in[783];
     assign  data_out[5314] = data_in[163];
     assign  data_out[5315] = data_in[748];
     assign  data_out[5316] = data_in[1031];
     assign  data_out[5317] = data_in[305];
     assign  data_out[5318] = data_in[1559];
     assign  data_out[5319] = data_in[1371];
     assign  data_out[5320] = data_in[44];
     assign  data_out[5321] = data_in[1336];
     assign  data_out[5322] = data_in[372];
     assign  data_out[5323] = data_in[495];
     assign  data_out[5324] = data_in[30];
     assign  data_out[5325] = data_in[141];
     assign  data_out[5326] = data_in[596];
     assign  data_out[5327] = data_in[17];
     assign  data_out[5328] = data_in[1179];
     assign  data_out[5329] = data_in[101];
     assign  data_out[5330] = data_in[107];
     assign  data_out[5331] = data_in[386];
     assign  data_out[5332] = data_in[52];
     assign  data_out[5333] = data_in[1404];
     assign  data_out[5334] = data_in[222];
     assign  data_out[5335] = data_in[1511];
     assign  data_out[5336] = data_in[19];
     assign  data_out[5337] = data_in[1047];
     assign  data_out[5338] = data_in[1587];
     assign  data_out[5339] = data_in[1495];
     assign  data_out[5340] = data_in[604];
     assign  data_out[5341] = data_in[830];
     assign  data_out[5342] = data_in[272];
     assign  data_out[5343] = data_in[1654];
     assign  data_out[5344] = data_in[772];
     assign  data_out[5345] = data_in[1163];
     assign  data_out[5346] = data_in[539];
     assign  data_out[5347] = data_in[1255];
     assign  data_out[5348] = data_in[245];
     assign  data_out[5349] = data_in[801];
     assign  data_out[5350] = data_in[1144];
     assign  data_out[5351] = data_in[825];
     assign  data_out[5352] = data_in[1037];
     assign  data_out[5353] = data_in[1076];
     assign  data_out[5354] = data_in[1007];
     assign  data_out[5355] = data_in[884];
     assign  data_out[5356] = data_in[217];
     assign  data_out[5357] = data_in[195];
     assign  data_out[5358] = data_in[131];
     assign  data_out[5359] = data_in[1156];
     assign  data_out[5360] = data_in[283];
     assign  data_out[5361] = data_in[331];
     assign  data_out[5362] = data_in[125];
     assign  data_out[5363] = data_in[937];
     assign  data_out[5364] = data_in[501];
     assign  data_out[5365] = data_in[1012];
     assign  data_out[5366] = data_in[935];
     assign  data_out[5367] = data_in[463];
     assign  data_out[5368] = data_in[778];
     assign  data_out[5369] = data_in[1526];
     assign  data_out[5370] = data_in[1626];
     assign  data_out[5371] = data_in[534];
     assign  data_out[5372] = data_in[428];
     assign  data_out[5373] = data_in[1386];
     assign  data_out[5374] = data_in[61];
     assign  data_out[5375] = data_in[216];
     assign  data_out[5376] = data_in[951];
     assign  data_out[5377] = data_in[850];
     assign  data_out[5378] = data_in[1055];
     assign  data_out[5379] = data_in[252];
     assign  data_out[5380] = data_in[350];
     assign  data_out[5381] = data_in[910];
     assign  data_out[5382] = data_in[219];
     assign  data_out[5383] = data_in[1634];
     assign  data_out[5384] = data_in[207];
     assign  data_out[5385] = data_in[1284];
     assign  data_out[5386] = data_in[1432];
     assign  data_out[5387] = data_in[56];
     assign  data_out[5388] = data_in[951];
     assign  data_out[5389] = data_in[997];
     assign  data_out[5390] = data_in[611];
     assign  data_out[5391] = data_in[261];
     assign  data_out[5392] = data_in[1360];
     assign  data_out[5393] = data_in[113];
     assign  data_out[5394] = data_in[625];
     assign  data_out[5395] = data_in[893];
     assign  data_out[5396] = data_in[174];
     assign  data_out[5397] = data_in[266];
     assign  data_out[5398] = data_in[392];
     assign  data_out[5399] = data_in[1501];
     assign  data_out[5400] = data_in[331];
     assign  data_out[5401] = data_in[835];
     assign  data_out[5402] = data_in[536];
     assign  data_out[5403] = data_in[1330];
     assign  data_out[5404] = data_in[1597];
     assign  data_out[5405] = data_in[515];
     assign  data_out[5406] = data_in[1485];
     assign  data_out[5407] = data_in[74];
     assign  data_out[5408] = data_in[1108];
     assign  data_out[5409] = data_in[1103];
     assign  data_out[5410] = data_in[89];
     assign  data_out[5411] = data_in[1311];
     assign  data_out[5412] = data_in[1427];
     assign  data_out[5413] = data_in[820];
     assign  data_out[5414] = data_in[382];
     assign  data_out[5415] = data_in[1170];
     assign  data_out[5416] = data_in[691];
     assign  data_out[5417] = data_in[1613];
     assign  data_out[5418] = data_in[1388];
     assign  data_out[5419] = data_in[949];
     assign  data_out[5420] = data_in[763];
     assign  data_out[5421] = data_in[481];
     assign  data_out[5422] = data_in[28];
     assign  data_out[5423] = data_in[332];
     assign  data_out[5424] = data_in[1028];
     assign  data_out[5425] = data_in[1383];
     assign  data_out[5426] = data_in[1417];
     assign  data_out[5427] = data_in[1262];
     assign  data_out[5428] = data_in[1663];
     assign  data_out[5429] = data_in[460];
     assign  data_out[5430] = data_in[324];
     assign  data_out[5431] = data_in[1590];
     assign  data_out[5432] = data_in[1304];
     assign  data_out[5433] = data_in[167];
     assign  data_out[5434] = data_in[353];
     assign  data_out[5435] = data_in[1666];
     assign  data_out[5436] = data_in[831];
     assign  data_out[5437] = data_in[1579];
     assign  data_out[5438] = data_in[80];
     assign  data_out[5439] = data_in[1230];
     assign  data_out[5440] = data_in[1670];
     assign  data_out[5441] = data_in[1080];
     assign  data_out[5442] = data_in[606];
     assign  data_out[5443] = data_in[1147];
     assign  data_out[5444] = data_in[1667];
     assign  data_out[5445] = data_in[1205];
     assign  data_out[5446] = data_in[43];
     assign  data_out[5447] = data_in[1175];
     assign  data_out[5448] = data_in[1148];
     assign  data_out[5449] = data_in[1340];
     assign  data_out[5450] = data_in[22];
     assign  data_out[5451] = data_in[1373];
     assign  data_out[5452] = data_in[1475];
     assign  data_out[5453] = data_in[522];
     assign  data_out[5454] = data_in[99];
     assign  data_out[5455] = data_in[102];
     assign  data_out[5456] = data_in[65];
     assign  data_out[5457] = data_in[515];
     assign  data_out[5458] = data_in[1714];
     assign  data_out[5459] = data_in[1377];
     assign  data_out[5460] = data_in[486];
     assign  data_out[5461] = data_in[1648];
     assign  data_out[5462] = data_in[1004];
     assign  data_out[5463] = data_in[340];
     assign  data_out[5464] = data_in[112];
     assign  data_out[5465] = data_in[338];
     assign  data_out[5466] = data_in[789];
     assign  data_out[5467] = data_in[1104];
     assign  data_out[5468] = data_in[1600];
     assign  data_out[5469] = data_in[1511];
     assign  data_out[5470] = data_in[289];
     assign  data_out[5471] = data_in[1147];
     assign  data_out[5472] = data_in[307];
     assign  data_out[5473] = data_in[1283];
     assign  data_out[5474] = data_in[1525];
     assign  data_out[5475] = data_in[1713];
     assign  data_out[5476] = data_in[829];
     assign  data_out[5477] = data_in[1495];
     assign  data_out[5478] = data_in[1339];
     assign  data_out[5479] = data_in[854];
     assign  data_out[5480] = data_in[936];
     assign  data_out[5481] = data_in[1091];
     assign  data_out[5482] = data_in[1069];
     assign  data_out[5483] = data_in[918];
     assign  data_out[5484] = data_in[1292];
     assign  data_out[5485] = data_in[25];
     assign  data_out[5486] = data_in[1086];
     assign  data_out[5487] = data_in[950];
     assign  data_out[5488] = data_in[1676];
     assign  data_out[5489] = data_in[418];
     assign  data_out[5490] = data_in[136];
     assign  data_out[5491] = data_in[627];
     assign  data_out[5492] = data_in[640];
     assign  data_out[5493] = data_in[913];
     assign  data_out[5494] = data_in[1249];
     assign  data_out[5495] = data_in[8];
     assign  data_out[5496] = data_in[787];
     assign  data_out[5497] = data_in[56];
     assign  data_out[5498] = data_in[965];
     assign  data_out[5499] = data_in[989];
     assign  data_out[5500] = data_in[300];
     assign  data_out[5501] = data_in[1188];
     assign  data_out[5502] = data_in[1646];
     assign  data_out[5503] = data_in[1663];
     assign  data_out[5504] = data_in[578];
     assign  data_out[5505] = data_in[113];
     assign  data_out[5506] = data_in[1168];
     assign  data_out[5507] = data_in[1560];
     assign  data_out[5508] = data_in[234];
     assign  data_out[5509] = data_in[1610];
     assign  data_out[5510] = data_in[1493];
     assign  data_out[5511] = data_in[333];
     assign  data_out[5512] = data_in[117];
     assign  data_out[5513] = data_in[1116];
     assign  data_out[5514] = data_in[760];
     assign  data_out[5515] = data_in[955];
     assign  data_out[5516] = data_in[1712];
     assign  data_out[5517] = data_in[109];
     assign  data_out[5518] = data_in[63];
     assign  data_out[5519] = data_in[1716];
     assign  data_out[5520] = data_in[1131];
     assign  data_out[5521] = data_in[164];
     assign  data_out[5522] = data_in[1621];
     assign  data_out[5523] = data_in[181];
     assign  data_out[5524] = data_in[776];
     assign  data_out[5525] = data_in[1006];
     assign  data_out[5526] = data_in[145];
     assign  data_out[5527] = data_in[313];
     assign  data_out[5528] = data_in[1149];
     assign  data_out[5529] = data_in[1111];
     assign  data_out[5530] = data_in[1133];
     assign  data_out[5531] = data_in[995];
     assign  data_out[5532] = data_in[76];
     assign  data_out[5533] = data_in[245];
     assign  data_out[5534] = data_in[495];
     assign  data_out[5535] = data_in[352];
     assign  data_out[5536] = data_in[1558];
     assign  data_out[5537] = data_in[774];
     assign  data_out[5538] = data_in[721];
     assign  data_out[5539] = data_in[1020];
     assign  data_out[5540] = data_in[1046];
     assign  data_out[5541] = data_in[224];
     assign  data_out[5542] = data_in[1453];
     assign  data_out[5543] = data_in[651];
     assign  data_out[5544] = data_in[1182];
     assign  data_out[5545] = data_in[1284];
     assign  data_out[5546] = data_in[1644];
     assign  data_out[5547] = data_in[1183];
     assign  data_out[5548] = data_in[618];
     assign  data_out[5549] = data_in[652];
     assign  data_out[5550] = data_in[1285];
     assign  data_out[5551] = data_in[433];
     assign  data_out[5552] = data_in[1312];
     assign  data_out[5553] = data_in[179];
     assign  data_out[5554] = data_in[145];
     assign  data_out[5555] = data_in[1264];
     assign  data_out[5556] = data_in[1109];
     assign  data_out[5557] = data_in[1711];
     assign  data_out[5558] = data_in[503];
     assign  data_out[5559] = data_in[163];
     assign  data_out[5560] = data_in[1447];
     assign  data_out[5561] = data_in[1454];
     assign  data_out[5562] = data_in[954];
     assign  data_out[5563] = data_in[844];
     assign  data_out[5564] = data_in[456];
     assign  data_out[5565] = data_in[528];
     assign  data_out[5566] = data_in[363];
     assign  data_out[5567] = data_in[886];
     assign  data_out[5568] = data_in[1297];
     assign  data_out[5569] = data_in[909];
     assign  data_out[5570] = data_in[774];
     assign  data_out[5571] = data_in[480];
     assign  data_out[5572] = data_in[806];
     assign  data_out[5573] = data_in[1683];
     assign  data_out[5574] = data_in[711];
     assign  data_out[5575] = data_in[313];
     assign  data_out[5576] = data_in[412];
     assign  data_out[5577] = data_in[1088];
     assign  data_out[5578] = data_in[492];
     assign  data_out[5579] = data_in[1355];
     assign  data_out[5580] = data_in[911];
     assign  data_out[5581] = data_in[288];
     assign  data_out[5582] = data_in[640];
     assign  data_out[5583] = data_in[1232];
     assign  data_out[5584] = data_in[621];
     assign  data_out[5585] = data_in[507];
     assign  data_out[5586] = data_in[1187];
     assign  data_out[5587] = data_in[1696];
     assign  data_out[5588] = data_in[1694];
     assign  data_out[5589] = data_in[1569];
     assign  data_out[5590] = data_in[221];
     assign  data_out[5591] = data_in[1113];
     assign  data_out[5592] = data_in[906];
     assign  data_out[5593] = data_in[389];
     assign  data_out[5594] = data_in[1221];
     assign  data_out[5595] = data_in[318];
     assign  data_out[5596] = data_in[807];
     assign  data_out[5597] = data_in[918];
     assign  data_out[5598] = data_in[1591];
     assign  data_out[5599] = data_in[946];
     assign  data_out[5600] = data_in[274];
     assign  data_out[5601] = data_in[1240];
     assign  data_out[5602] = data_in[1325];
     assign  data_out[5603] = data_in[382];
     assign  data_out[5604] = data_in[353];
     assign  data_out[5605] = data_in[452];
     assign  data_out[5606] = data_in[755];
     assign  data_out[5607] = data_in[469];
     assign  data_out[5608] = data_in[1701];
     assign  data_out[5609] = data_in[1371];
     assign  data_out[5610] = data_in[392];
     assign  data_out[5611] = data_in[1277];
     assign  data_out[5612] = data_in[149];
     assign  data_out[5613] = data_in[1596];
     assign  data_out[5614] = data_in[1195];
     assign  data_out[5615] = data_in[526];
     assign  data_out[5616] = data_in[1614];
     assign  data_out[5617] = data_in[818];
     assign  data_out[5618] = data_in[989];
     assign  data_out[5619] = data_in[1083];
     assign  data_out[5620] = data_in[696];
     assign  data_out[5621] = data_in[1334];
     assign  data_out[5622] = data_in[922];
     assign  data_out[5623] = data_in[451];
     assign  data_out[5624] = data_in[1180];
     assign  data_out[5625] = data_in[299];
     assign  data_out[5626] = data_in[405];
     assign  data_out[5627] = data_in[977];
     assign  data_out[5628] = data_in[332];
     assign  data_out[5629] = data_in[777];
     assign  data_out[5630] = data_in[1336];
     assign  data_out[5631] = data_in[858];
     assign  data_out[5632] = data_in[1399];
     assign  data_out[5633] = data_in[381];
     assign  data_out[5634] = data_in[49];
     assign  data_out[5635] = data_in[1220];
     assign  data_out[5636] = data_in[362];
     assign  data_out[5637] = data_in[119];
     assign  data_out[5638] = data_in[1616];
     assign  data_out[5639] = data_in[1458];
     assign  data_out[5640] = data_in[1008];
     assign  data_out[5641] = data_in[868];
     assign  data_out[5642] = data_in[382];
     assign  data_out[5643] = data_in[809];
     assign  data_out[5644] = data_in[910];
     assign  data_out[5645] = data_in[725];
     assign  data_out[5646] = data_in[1105];
     assign  data_out[5647] = data_in[828];
     assign  data_out[5648] = data_in[642];
     assign  data_out[5649] = data_in[400];
     assign  data_out[5650] = data_in[388];
     assign  data_out[5651] = data_in[809];
     assign  data_out[5652] = data_in[1301];
     assign  data_out[5653] = data_in[518];
     assign  data_out[5654] = data_in[1045];
     assign  data_out[5655] = data_in[1569];
     assign  data_out[5656] = data_in[1169];
     assign  data_out[5657] = data_in[1458];
     assign  data_out[5658] = data_in[1569];
     assign  data_out[5659] = data_in[981];
     assign  data_out[5660] = data_in[1530];
     assign  data_out[5661] = data_in[1684];
     assign  data_out[5662] = data_in[477];
     assign  data_out[5663] = data_in[138];
     assign  data_out[5664] = data_in[1373];
     assign  data_out[5665] = data_in[25];
     assign  data_out[5666] = data_in[938];
     assign  data_out[5667] = data_in[87];
     assign  data_out[5668] = data_in[1347];
     assign  data_out[5669] = data_in[1305];
     assign  data_out[5670] = data_in[138];
     assign  data_out[5671] = data_in[1081];
     assign  data_out[5672] = data_in[176];
     assign  data_out[5673] = data_in[1395];
     assign  data_out[5674] = data_in[636];
     assign  data_out[5675] = data_in[1594];
     assign  data_out[5676] = data_in[428];
     assign  data_out[5677] = data_in[1226];
     assign  data_out[5678] = data_in[523];
     assign  data_out[5679] = data_in[383];
     assign  data_out[5680] = data_in[1668];
     assign  data_out[5681] = data_in[1623];
     assign  data_out[5682] = data_in[1349];
     assign  data_out[5683] = data_in[587];
     assign  data_out[5684] = data_in[1349];
     assign  data_out[5685] = data_in[850];
     assign  data_out[5686] = data_in[1026];
     assign  data_out[5687] = data_in[134];
     assign  data_out[5688] = data_in[475];
     assign  data_out[5689] = data_in[308];
     assign  data_out[5690] = data_in[267];
     assign  data_out[5691] = data_in[271];
     assign  data_out[5692] = data_in[1552];
     assign  data_out[5693] = data_in[519];
     assign  data_out[5694] = data_in[168];
     assign  data_out[5695] = data_in[949];
     assign  data_out[5696] = data_in[1052];
     assign  data_out[5697] = data_in[1488];
     assign  data_out[5698] = data_in[479];
     assign  data_out[5699] = data_in[1042];
     assign  data_out[5700] = data_in[203];
     assign  data_out[5701] = data_in[1659];
     assign  data_out[5702] = data_in[349];
     assign  data_out[5703] = data_in[1515];
     assign  data_out[5704] = data_in[21];
     assign  data_out[5705] = data_in[932];
     assign  data_out[5706] = data_in[731];
     assign  data_out[5707] = data_in[144];
     assign  data_out[5708] = data_in[957];
     assign  data_out[5709] = data_in[221];
     assign  data_out[5710] = data_in[1597];
     assign  data_out[5711] = data_in[87];
     assign  data_out[5712] = data_in[714];
     assign  data_out[5713] = data_in[1291];
     assign  data_out[5714] = data_in[64];
     assign  data_out[5715] = data_in[183];
     assign  data_out[5716] = data_in[247];
     assign  data_out[5717] = data_in[1084];
     assign  data_out[5718] = data_in[1570];
     assign  data_out[5719] = data_in[1374];
     assign  data_out[5720] = data_in[1131];
     assign  data_out[5721] = data_in[1552];
     assign  data_out[5722] = data_in[101];
     assign  data_out[5723] = data_in[570];
     assign  data_out[5724] = data_in[844];
     assign  data_out[5725] = data_in[1561];
     assign  data_out[5726] = data_in[100];
     assign  data_out[5727] = data_in[1185];
     assign  data_out[5728] = data_in[268];
     assign  data_out[5729] = data_in[521];
     assign  data_out[5730] = data_in[1479];
     assign  data_out[5731] = data_in[1285];
     assign  data_out[5732] = data_in[574];
     assign  data_out[5733] = data_in[1045];
     assign  data_out[5734] = data_in[1362];
     assign  data_out[5735] = data_in[669];
     assign  data_out[5736] = data_in[335];
     assign  data_out[5737] = data_in[537];
     assign  data_out[5738] = data_in[1380];
     assign  data_out[5739] = data_in[1665];
     assign  data_out[5740] = data_in[1135];
     assign  data_out[5741] = data_in[505];
     assign  data_out[5742] = data_in[1566];
     assign  data_out[5743] = data_in[21];
     assign  data_out[5744] = data_in[1421];
     assign  data_out[5745] = data_in[1018];
     assign  data_out[5746] = data_in[769];
     assign  data_out[5747] = data_in[1144];
     assign  data_out[5748] = data_in[696];
     assign  data_out[5749] = data_in[465];
     assign  data_out[5750] = data_in[197];
     assign  data_out[5751] = data_in[1064];
     assign  data_out[5752] = data_in[687];
     assign  data_out[5753] = data_in[876];
     assign  data_out[5754] = data_in[623];
     assign  data_out[5755] = data_in[200];
     assign  data_out[5756] = data_in[1418];
     assign  data_out[5757] = data_in[934];
     assign  data_out[5758] = data_in[237];
     assign  data_out[5759] = data_in[1391];
     assign  data_out[5760] = data_in[1283];
     assign  data_out[5761] = data_in[1141];
     assign  data_out[5762] = data_in[963];
     assign  data_out[5763] = data_in[1528];
     assign  data_out[5764] = data_in[762];
     assign  data_out[5765] = data_in[1541];
     assign  data_out[5766] = data_in[830];
     assign  data_out[5767] = data_in[825];
     assign  data_out[5768] = data_in[1611];
     assign  data_out[5769] = data_in[891];
     assign  data_out[5770] = data_in[974];
     assign  data_out[5771] = data_in[1050];
     assign  data_out[5772] = data_in[1163];
     assign  data_out[5773] = data_in[171];
     assign  data_out[5774] = data_in[1390];
     assign  data_out[5775] = data_in[1187];
     assign  data_out[5776] = data_in[1217];
     assign  data_out[5777] = data_in[308];
     assign  data_out[5778] = data_in[193];
     assign  data_out[5779] = data_in[1616];
     assign  data_out[5780] = data_in[49];
     assign  data_out[5781] = data_in[449];
     assign  data_out[5782] = data_in[1608];
     assign  data_out[5783] = data_in[1084];
     assign  data_out[5784] = data_in[850];
     assign  data_out[5785] = data_in[500];
     assign  data_out[5786] = data_in[790];
     assign  data_out[5787] = data_in[992];
     assign  data_out[5788] = data_in[1668];
     assign  data_out[5789] = data_in[431];
     assign  data_out[5790] = data_in[813];
     assign  data_out[5791] = data_in[1297];
     assign  data_out[5792] = data_in[149];
     assign  data_out[5793] = data_in[72];
     assign  data_out[5794] = data_in[549];
     assign  data_out[5795] = data_in[807];
     assign  data_out[5796] = data_in[630];
     assign  data_out[5797] = data_in[526];
     assign  data_out[5798] = data_in[136];
     assign  data_out[5799] = data_in[3];
     assign  data_out[5800] = data_in[1589];
     assign  data_out[5801] = data_in[569];
     assign  data_out[5802] = data_in[765];
     assign  data_out[5803] = data_in[157];
     assign  data_out[5804] = data_in[1084];
     assign  data_out[5805] = data_in[1258];
     assign  data_out[5806] = data_in[575];
     assign  data_out[5807] = data_in[319];
     assign  data_out[5808] = data_in[1689];
     assign  data_out[5809] = data_in[19];
     assign  data_out[5810] = data_in[1385];
     assign  data_out[5811] = data_in[1527];
     assign  data_out[5812] = data_in[683];
     assign  data_out[5813] = data_in[1250];
     assign  data_out[5814] = data_in[408];
     assign  data_out[5815] = data_in[774];
     assign  data_out[5816] = data_in[576];
     assign  data_out[5817] = data_in[536];
     assign  data_out[5818] = data_in[694];
     assign  data_out[5819] = data_in[1376];
     assign  data_out[5820] = data_in[1553];
     assign  data_out[5821] = data_in[606];
     assign  data_out[5822] = data_in[602];
     assign  data_out[5823] = data_in[1554];
     assign  data_out[5824] = data_in[530];
     assign  data_out[5825] = data_in[574];
     assign  data_out[5826] = data_in[1260];
     assign  data_out[5827] = data_in[1670];
     assign  data_out[5828] = data_in[1612];
     assign  data_out[5829] = data_in[1051];
     assign  data_out[5830] = data_in[929];
     assign  data_out[5831] = data_in[594];
     assign  data_out[5832] = data_in[436];
     assign  data_out[5833] = data_in[1222];
     assign  data_out[5834] = data_in[1412];
     assign  data_out[5835] = data_in[898];
     assign  data_out[5836] = data_in[777];
     assign  data_out[5837] = data_in[1104];
     assign  data_out[5838] = data_in[622];
     assign  data_out[5839] = data_in[256];
     assign  data_out[5840] = data_in[1669];
     assign  data_out[5841] = data_in[627];
     assign  data_out[5842] = data_in[1614];
     assign  data_out[5843] = data_in[859];
     assign  data_out[5844] = data_in[1356];
     assign  data_out[5845] = data_in[114];
     assign  data_out[5846] = data_in[111];
     assign  data_out[5847] = data_in[393];
     assign  data_out[5848] = data_in[1247];
     assign  data_out[5849] = data_in[721];
     assign  data_out[5850] = data_in[1560];
     assign  data_out[5851] = data_in[1563];
     assign  data_out[5852] = data_in[873];
     assign  data_out[5853] = data_in[768];
     assign  data_out[5854] = data_in[379];
     assign  data_out[5855] = data_in[273];
     assign  data_out[5856] = data_in[1612];
     assign  data_out[5857] = data_in[342];
     assign  data_out[5858] = data_in[69];
     assign  data_out[5859] = data_in[1532];
     assign  data_out[5860] = data_in[1519];
     assign  data_out[5861] = data_in[1466];
     assign  data_out[5862] = data_in[1675];
     assign  data_out[5863] = data_in[723];
     assign  data_out[5864] = data_in[753];
     assign  data_out[5865] = data_in[669];
     assign  data_out[5866] = data_in[1251];
     assign  data_out[5867] = data_in[56];
     assign  data_out[5868] = data_in[1685];
     assign  data_out[5869] = data_in[992];
     assign  data_out[5870] = data_in[1577];
     assign  data_out[5871] = data_in[1296];
     assign  data_out[5872] = data_in[692];
     assign  data_out[5873] = data_in[505];
     assign  data_out[5874] = data_in[1013];
     assign  data_out[5875] = data_in[1376];
     assign  data_out[5876] = data_in[666];
     assign  data_out[5877] = data_in[1683];
     assign  data_out[5878] = data_in[1044];
     assign  data_out[5879] = data_in[1117];
     assign  data_out[5880] = data_in[1495];
     assign  data_out[5881] = data_in[412];
     assign  data_out[5882] = data_in[564];
     assign  data_out[5883] = data_in[89];
     assign  data_out[5884] = data_in[990];
     assign  data_out[5885] = data_in[714];
     assign  data_out[5886] = data_in[1185];
     assign  data_out[5887] = data_in[1670];
     assign  data_out[5888] = data_in[1552];
     assign  data_out[5889] = data_in[152];
     assign  data_out[5890] = data_in[267];
     assign  data_out[5891] = data_in[1322];
     assign  data_out[5892] = data_in[1459];
     assign  data_out[5893] = data_in[610];
     assign  data_out[5894] = data_in[1108];
     assign  data_out[5895] = data_in[1162];
     assign  data_out[5896] = data_in[657];
     assign  data_out[5897] = data_in[1536];
     assign  data_out[5898] = data_in[1482];
     assign  data_out[5899] = data_in[1380];
     assign  data_out[5900] = data_in[1636];
     assign  data_out[5901] = data_in[959];
     assign  data_out[5902] = data_in[296];
     assign  data_out[5903] = data_in[1200];
     assign  data_out[5904] = data_in[723];
     assign  data_out[5905] = data_in[1103];
     assign  data_out[5906] = data_in[848];
     assign  data_out[5907] = data_in[1440];
     assign  data_out[5908] = data_in[502];
     assign  data_out[5909] = data_in[717];
     assign  data_out[5910] = data_in[348];
     assign  data_out[5911] = data_in[1585];
     assign  data_out[5912] = data_in[652];
     assign  data_out[5913] = data_in[315];
     assign  data_out[5914] = data_in[1199];
     assign  data_out[5915] = data_in[732];
     assign  data_out[5916] = data_in[1380];
     assign  data_out[5917] = data_in[726];
     assign  data_out[5918] = data_in[880];
     assign  data_out[5919] = data_in[507];
     assign  data_out[5920] = data_in[936];
     assign  data_out[5921] = data_in[402];
     assign  data_out[5922] = data_in[1095];
     assign  data_out[5923] = data_in[292];
     assign  data_out[5924] = data_in[651];
     assign  data_out[5925] = data_in[1263];
     assign  data_out[5926] = data_in[1689];
     assign  data_out[5927] = data_in[144];
     assign  data_out[5928] = data_in[695];
     assign  data_out[5929] = data_in[884];
     assign  data_out[5930] = data_in[979];
     assign  data_out[5931] = data_in[30];
     assign  data_out[5932] = data_in[23];
     assign  data_out[5933] = data_in[1532];
     assign  data_out[5934] = data_in[821];
     assign  data_out[5935] = data_in[376];
     assign  data_out[5936] = data_in[972];
     assign  data_out[5937] = data_in[37];
     assign  data_out[5938] = data_in[63];
     assign  data_out[5939] = data_in[1194];
     assign  data_out[5940] = data_in[865];
     assign  data_out[5941] = data_in[1104];
     assign  data_out[5942] = data_in[621];
     assign  data_out[5943] = data_in[1353];
     assign  data_out[5944] = data_in[479];
     assign  data_out[5945] = data_in[762];
     assign  data_out[5946] = data_in[1182];
     assign  data_out[5947] = data_in[407];
     assign  data_out[5948] = data_in[1352];
     assign  data_out[5949] = data_in[1572];
     assign  data_out[5950] = data_in[1045];
     assign  data_out[5951] = data_in[1108];
     assign  data_out[5952] = data_in[1056];
     assign  data_out[5953] = data_in[1110];
     assign  data_out[5954] = data_in[1199];
     assign  data_out[5955] = data_in[1204];
     assign  data_out[5956] = data_in[1604];
     assign  data_out[5957] = data_in[1506];
     assign  data_out[5958] = data_in[965];
     assign  data_out[5959] = data_in[278];
     assign  data_out[5960] = data_in[387];
     assign  data_out[5961] = data_in[581];
     assign  data_out[5962] = data_in[1483];
     assign  data_out[5963] = data_in[1593];
     assign  data_out[5964] = data_in[1260];
     assign  data_out[5965] = data_in[265];
     assign  data_out[5966] = data_in[550];
     assign  data_out[5967] = data_in[148];
     assign  data_out[5968] = data_in[1352];
     assign  data_out[5969] = data_in[1457];
     assign  data_out[5970] = data_in[463];
     assign  data_out[5971] = data_in[837];
     assign  data_out[5972] = data_in[1592];
     assign  data_out[5973] = data_in[305];
     assign  data_out[5974] = data_in[1271];
     assign  data_out[5975] = data_in[897];
     assign  data_out[5976] = data_in[1713];
     assign  data_out[5977] = data_in[1703];
     assign  data_out[5978] = data_in[1089];
     assign  data_out[5979] = data_in[1271];
     assign  data_out[5980] = data_in[58];
     assign  data_out[5981] = data_in[1051];
     assign  data_out[5982] = data_in[79];
     assign  data_out[5983] = data_in[72];
     assign  data_out[5984] = data_in[446];
     assign  data_out[5985] = data_in[189];
     assign  data_out[5986] = data_in[362];
     assign  data_out[5987] = data_in[1692];
     assign  data_out[5988] = data_in[1486];
     assign  data_out[5989] = data_in[1634];
     assign  data_out[5990] = data_in[209];
     assign  data_out[5991] = data_in[1632];
     assign  data_out[5992] = data_in[1686];
     assign  data_out[5993] = data_in[391];
     assign  data_out[5994] = data_in[681];
     assign  data_out[5995] = data_in[1338];
     assign  data_out[5996] = data_in[962];
     assign  data_out[5997] = data_in[384];
     assign  data_out[5998] = data_in[607];
     assign  data_out[5999] = data_in[1031];
     assign  data_out[6000] = data_in[749];
     assign  data_out[6001] = data_in[495];
     assign  data_out[6002] = data_in[1533];
     assign  data_out[6003] = data_in[620];
     assign  data_out[6004] = data_in[634];
     assign  data_out[6005] = data_in[1449];
     assign  data_out[6006] = data_in[250];
     assign  data_out[6007] = data_in[1609];
     assign  data_out[6008] = data_in[608];
     assign  data_out[6009] = data_in[984];
     assign  data_out[6010] = data_in[904];
     assign  data_out[6011] = data_in[348];
     assign  data_out[6012] = data_in[1670];
     assign  data_out[6013] = data_in[902];
     assign  data_out[6014] = data_in[104];
     assign  data_out[6015] = data_in[101];
     assign  data_out[6016] = data_in[72];
     assign  data_out[6017] = data_in[358];
     assign  data_out[6018] = data_in[1226];
     assign  data_out[6019] = data_in[1170];
     assign  data_out[6020] = data_in[754];
     assign  data_out[6021] = data_in[702];
     assign  data_out[6022] = data_in[964];
     assign  data_out[6023] = data_in[11];
     assign  data_out[6024] = data_in[332];
     assign  data_out[6025] = data_in[1426];
     assign  data_out[6026] = data_in[853];
     assign  data_out[6027] = data_in[1501];
     assign  data_out[6028] = data_in[1490];
     assign  data_out[6029] = data_in[416];
     assign  data_out[6030] = data_in[658];
     assign  data_out[6031] = data_in[1003];
     assign  data_out[6032] = data_in[481];
     assign  data_out[6033] = data_in[544];
     assign  data_out[6034] = data_in[435];
     assign  data_out[6035] = data_in[849];
     assign  data_out[6036] = data_in[960];
     assign  data_out[6037] = data_in[1242];
     assign  data_out[6038] = data_in[965];
     assign  data_out[6039] = data_in[615];
     assign  data_out[6040] = data_in[1032];
     assign  data_out[6041] = data_in[1256];
     assign  data_out[6042] = data_in[17];
     assign  data_out[6043] = data_in[1630];
     assign  data_out[6044] = data_in[1556];
     assign  data_out[6045] = data_in[1624];
     assign  data_out[6046] = data_in[57];
     assign  data_out[6047] = data_in[1360];
     assign  data_out[6048] = data_in[1603];
     assign  data_out[6049] = data_in[501];
     assign  data_out[6050] = data_in[657];
     assign  data_out[6051] = data_in[836];
     assign  data_out[6052] = data_in[1435];
     assign  data_out[6053] = data_in[1706];
     assign  data_out[6054] = data_in[1585];
     assign  data_out[6055] = data_in[775];
     assign  data_out[6056] = data_in[1409];
     assign  data_out[6057] = data_in[963];
     assign  data_out[6058] = data_in[226];
     assign  data_out[6059] = data_in[918];
     assign  data_out[6060] = data_in[1589];
     assign  data_out[6061] = data_in[1102];
     assign  data_out[6062] = data_in[640];
     assign  data_out[6063] = data_in[687];
     assign  data_out[6064] = data_in[838];
     assign  data_out[6065] = data_in[1165];
     assign  data_out[6066] = data_in[650];
     assign  data_out[6067] = data_in[156];
     assign  data_out[6068] = data_in[194];
     assign  data_out[6069] = data_in[331];
     assign  data_out[6070] = data_in[178];
     assign  data_out[6071] = data_in[1144];
     assign  data_out[6072] = data_in[644];
     assign  data_out[6073] = data_in[1337];
     assign  data_out[6074] = data_in[679];
     assign  data_out[6075] = data_in[523];
     assign  data_out[6076] = data_in[111];
     assign  data_out[6077] = data_in[745];
     assign  data_out[6078] = data_in[875];
     assign  data_out[6079] = data_in[1474];
     assign  data_out[6080] = data_in[495];
     assign  data_out[6081] = data_in[855];
     assign  data_out[6082] = data_in[108];
     assign  data_out[6083] = data_in[212];
     assign  data_out[6084] = data_in[208];
     assign  data_out[6085] = data_in[1215];
     assign  data_out[6086] = data_in[701];
     assign  data_out[6087] = data_in[1565];
     assign  data_out[6088] = data_in[334];
     assign  data_out[6089] = data_in[1089];
     assign  data_out[6090] = data_in[1619];
     assign  data_out[6091] = data_in[203];
     assign  data_out[6092] = data_in[1572];
     assign  data_out[6093] = data_in[213];
     assign  data_out[6094] = data_in[759];
     assign  data_out[6095] = data_in[1624];
     assign  data_out[6096] = data_in[1085];
     assign  data_out[6097] = data_in[1540];
     assign  data_out[6098] = data_in[1606];
     assign  data_out[6099] = data_in[682];
     assign  data_out[6100] = data_in[982];
     assign  data_out[6101] = data_in[1575];
     assign  data_out[6102] = data_in[109];
     assign  data_out[6103] = data_in[430];
     assign  data_out[6104] = data_in[1259];
     assign  data_out[6105] = data_in[1394];
     assign  data_out[6106] = data_in[1092];
     assign  data_out[6107] = data_in[1125];
     assign  data_out[6108] = data_in[1018];
     assign  data_out[6109] = data_in[1463];
     assign  data_out[6110] = data_in[306];
     assign  data_out[6111] = data_in[716];
     assign  data_out[6112] = data_in[1548];
     assign  data_out[6113] = data_in[1277];
     assign  data_out[6114] = data_in[442];
     assign  data_out[6115] = data_in[602];
     assign  data_out[6116] = data_in[502];
     assign  data_out[6117] = data_in[1468];
     assign  data_out[6118] = data_in[664];
     assign  data_out[6119] = data_in[938];
     assign  data_out[6120] = data_in[137];
     assign  data_out[6121] = data_in[53];
     assign  data_out[6122] = data_in[345];
     assign  data_out[6123] = data_in[29];
     assign  data_out[6124] = data_in[1585];
     assign  data_out[6125] = data_in[1191];
     assign  data_out[6126] = data_in[1492];
     assign  data_out[6127] = data_in[1089];
     assign  data_out[6128] = data_in[1188];
     assign  data_out[6129] = data_in[473];
     assign  data_out[6130] = data_in[412];
     assign  data_out[6131] = data_in[1169];
     assign  data_out[6132] = data_in[627];
     assign  data_out[6133] = data_in[1411];
     assign  data_out[6134] = data_in[1515];
     assign  data_out[6135] = data_in[83];
     assign  data_out[6136] = data_in[212];
     assign  data_out[6137] = data_in[1216];
     assign  data_out[6138] = data_in[590];
     assign  data_out[6139] = data_in[678];
     assign  data_out[6140] = data_in[890];
     assign  data_out[6141] = data_in[551];
     assign  data_out[6142] = data_in[1554];
     assign  data_out[6143] = data_in[276];
     assign  data_out[6144] = data_in[1624];
     assign  data_out[6145] = data_in[1244];
     assign  data_out[6146] = data_in[197];
     assign  data_out[6147] = data_in[1639];
     assign  data_out[6148] = data_in[401];
     assign  data_out[6149] = data_in[8];
     assign  data_out[6150] = data_in[640];
     assign  data_out[6151] = data_in[98];
     assign  data_out[6152] = data_in[1097];
     assign  data_out[6153] = data_in[911];
     assign  data_out[6154] = data_in[1490];
     assign  data_out[6155] = data_in[1118];
     assign  data_out[6156] = data_in[1617];
     assign  data_out[6157] = data_in[1052];
     assign  data_out[6158] = data_in[127];
     assign  data_out[6159] = data_in[731];
     assign  data_out[6160] = data_in[88];
     assign  data_out[6161] = data_in[1574];
     assign  data_out[6162] = data_in[494];
     assign  data_out[6163] = data_in[409];
     assign  data_out[6164] = data_in[1449];
     assign  data_out[6165] = data_in[214];
     assign  data_out[6166] = data_in[245];
     assign  data_out[6167] = data_in[901];
     assign  data_out[6168] = data_in[722];
     assign  data_out[6169] = data_in[216];
     assign  data_out[6170] = data_in[1373];
     assign  data_out[6171] = data_in[1662];
     assign  data_out[6172] = data_in[1362];
     assign  data_out[6173] = data_in[451];
     assign  data_out[6174] = data_in[1180];
     assign  data_out[6175] = data_in[534];
     assign  data_out[6176] = data_in[15];
     assign  data_out[6177] = data_in[1586];
     assign  data_out[6178] = data_in[775];
     assign  data_out[6179] = data_in[1278];
     assign  data_out[6180] = data_in[1282];
     assign  data_out[6181] = data_in[47];
     assign  data_out[6182] = data_in[67];
     assign  data_out[6183] = data_in[1167];
     assign  data_out[6184] = data_in[735];
     assign  data_out[6185] = data_in[1159];
     assign  data_out[6186] = data_in[907];
     assign  data_out[6187] = data_in[794];
     assign  data_out[6188] = data_in[1492];
     assign  data_out[6189] = data_in[751];
     assign  data_out[6190] = data_in[1139];
     assign  data_out[6191] = data_in[1389];
     assign  data_out[6192] = data_in[884];
     assign  data_out[6193] = data_in[1162];
     assign  data_out[6194] = data_in[1229];
     assign  data_out[6195] = data_in[706];
     assign  data_out[6196] = data_in[425];
     assign  data_out[6197] = data_in[576];
     assign  data_out[6198] = data_in[1052];
     assign  data_out[6199] = data_in[1144];
     assign  data_out[6200] = data_in[1529];
     assign  data_out[6201] = data_in[883];
     assign  data_out[6202] = data_in[1587];
     assign  data_out[6203] = data_in[1426];
     assign  data_out[6204] = data_in[448];
     assign  data_out[6205] = data_in[635];
     assign  data_out[6206] = data_in[1200];
     assign  data_out[6207] = data_in[1060];
     assign  data_out[6208] = data_in[170];
     assign  data_out[6209] = data_in[1026];
     assign  data_out[6210] = data_in[1254];
     assign  data_out[6211] = data_in[987];
     assign  data_out[6212] = data_in[904];
     assign  data_out[6213] = data_in[97];
     assign  data_out[6214] = data_in[379];
     assign  data_out[6215] = data_in[271];
     assign  data_out[6216] = data_in[734];
     assign  data_out[6217] = data_in[1368];
     assign  data_out[6218] = data_in[767];
     assign  data_out[6219] = data_in[1616];
     assign  data_out[6220] = data_in[873];
     assign  data_out[6221] = data_in[5];
     assign  data_out[6222] = data_in[629];
     assign  data_out[6223] = data_in[1364];
     assign  data_out[6224] = data_in[464];
     assign  data_out[6225] = data_in[364];
     assign  data_out[6226] = data_in[1398];
     assign  data_out[6227] = data_in[963];
     assign  data_out[6228] = data_in[1281];
     assign  data_out[6229] = data_in[389];
     assign  data_out[6230] = data_in[323];
     assign  data_out[6231] = data_in[1719];
     assign  data_out[6232] = data_in[344];
     assign  data_out[6233] = data_in[144];
     assign  data_out[6234] = data_in[514];
     assign  data_out[6235] = data_in[829];
     assign  data_out[6236] = data_in[1187];
     assign  data_out[6237] = data_in[1061];
     assign  data_out[6238] = data_in[441];
     assign  data_out[6239] = data_in[614];
     assign  data_out[6240] = data_in[1057];
     assign  data_out[6241] = data_in[1365];
     assign  data_out[6242] = data_in[119];
     assign  data_out[6243] = data_in[558];
     assign  data_out[6244] = data_in[322];
     assign  data_out[6245] = data_in[887];
     assign  data_out[6246] = data_in[1554];
     assign  data_out[6247] = data_in[1369];
     assign  data_out[6248] = data_in[21];
     assign  data_out[6249] = data_in[6];
     assign  data_out[6250] = data_in[917];
     assign  data_out[6251] = data_in[1016];
     assign  data_out[6252] = data_in[989];
     assign  data_out[6253] = data_in[742];
     assign  data_out[6254] = data_in[154];
     assign  data_out[6255] = data_in[1604];
     assign  data_out[6256] = data_in[1604];
     assign  data_out[6257] = data_in[1656];
     assign  data_out[6258] = data_in[916];
     assign  data_out[6259] = data_in[135];
     assign  data_out[6260] = data_in[671];
     assign  data_out[6261] = data_in[1488];
     assign  data_out[6262] = data_in[1626];
     assign  data_out[6263] = data_in[994];
     assign  data_out[6264] = data_in[766];
     assign  data_out[6265] = data_in[1460];
     assign  data_out[6266] = data_in[298];
     assign  data_out[6267] = data_in[784];
     assign  data_out[6268] = data_in[1271];
     assign  data_out[6269] = data_in[445];
     assign  data_out[6270] = data_in[1461];
     assign  data_out[6271] = data_in[602];
     assign  data_out[6272] = data_in[618];
     assign  data_out[6273] = data_in[570];
     assign  data_out[6274] = data_in[446];
     assign  data_out[6275] = data_in[1567];
     assign  data_out[6276] = data_in[426];
     assign  data_out[6277] = data_in[175];
     assign  data_out[6278] = data_in[381];
     assign  data_out[6279] = data_in[696];
     assign  data_out[6280] = data_in[1680];
     assign  data_out[6281] = data_in[344];
     assign  data_out[6282] = data_in[613];
     assign  data_out[6283] = data_in[1661];
     assign  data_out[6284] = data_in[1179];
     assign  data_out[6285] = data_in[194];
     assign  data_out[6286] = data_in[1539];
     assign  data_out[6287] = data_in[518];
     assign  data_out[6288] = data_in[867];
     assign  data_out[6289] = data_in[223];
     assign  data_out[6290] = data_in[836];
     assign  data_out[6291] = data_in[687];
     assign  data_out[6292] = data_in[268];
     assign  data_out[6293] = data_in[1009];
     assign  data_out[6294] = data_in[159];
     assign  data_out[6295] = data_in[1713];
     assign  data_out[6296] = data_in[182];
     assign  data_out[6297] = data_in[1003];
     assign  data_out[6298] = data_in[759];
     assign  data_out[6299] = data_in[531];
     assign  data_out[6300] = data_in[1686];
     assign  data_out[6301] = data_in[1447];
     assign  data_out[6302] = data_in[172];
     assign  data_out[6303] = data_in[1621];
     assign  data_out[6304] = data_in[952];
     assign  data_out[6305] = data_in[1413];
     assign  data_out[6306] = data_in[1260];
     assign  data_out[6307] = data_in[458];
     assign  data_out[6308] = data_in[219];
     assign  data_out[6309] = data_in[1388];
     assign  data_out[6310] = data_in[834];
     assign  data_out[6311] = data_in[590];
     assign  data_out[6312] = data_in[860];
     assign  data_out[6313] = data_in[93];
     assign  data_out[6314] = data_in[243];
     assign  data_out[6315] = data_in[1090];
     assign  data_out[6316] = data_in[621];
     assign  data_out[6317] = data_in[1263];
     assign  data_out[6318] = data_in[1697];
     assign  data_out[6319] = data_in[888];
     assign  data_out[6320] = data_in[704];
     assign  data_out[6321] = data_in[1242];
     assign  data_out[6322] = data_in[1611];
     assign  data_out[6323] = data_in[1685];
     assign  data_out[6324] = data_in[1585];
     assign  data_out[6325] = data_in[32];
     assign  data_out[6326] = data_in[29];
     assign  data_out[6327] = data_in[624];
     assign  data_out[6328] = data_in[139];
     assign  data_out[6329] = data_in[1479];
     assign  data_out[6330] = data_in[1126];
     assign  data_out[6331] = data_in[1092];
     assign  data_out[6332] = data_in[1527];
     assign  data_out[6333] = data_in[297];
     assign  data_out[6334] = data_in[1397];
     assign  data_out[6335] = data_in[0];
     assign  data_out[6336] = data_in[1405];
     assign  data_out[6337] = data_in[1107];
     assign  data_out[6338] = data_in[991];
     assign  data_out[6339] = data_in[642];
     assign  data_out[6340] = data_in[266];
     assign  data_out[6341] = data_in[1528];
     assign  data_out[6342] = data_in[243];
     assign  data_out[6343] = data_in[851];
     assign  data_out[6344] = data_in[320];
     assign  data_out[6345] = data_in[42];
     assign  data_out[6346] = data_in[1329];
     assign  data_out[6347] = data_in[351];
     assign  data_out[6348] = data_in[56];
     assign  data_out[6349] = data_in[422];
     assign  data_out[6350] = data_in[1267];
     assign  data_out[6351] = data_in[1232];
     assign  data_out[6352] = data_in[813];
     assign  data_out[6353] = data_in[871];
     assign  data_out[6354] = data_in[1377];
     assign  data_out[6355] = data_in[517];
     assign  data_out[6356] = data_in[788];
     assign  data_out[6357] = data_in[121];
     assign  data_out[6358] = data_in[430];
     assign  data_out[6359] = data_in[578];
     assign  data_out[6360] = data_in[1156];
     assign  data_out[6361] = data_in[32];
     assign  data_out[6362] = data_in[32];
     assign  data_out[6363] = data_in[85];
     assign  data_out[6364] = data_in[1457];
     assign  data_out[6365] = data_in[626];
     assign  data_out[6366] = data_in[1590];
     assign  data_out[6367] = data_in[1627];
     assign  data_out[6368] = data_in[296];
     assign  data_out[6369] = data_in[1668];
     assign  data_out[6370] = data_in[933];
     assign  data_out[6371] = data_in[400];
     assign  data_out[6372] = data_in[974];
     assign  data_out[6373] = data_in[1538];
     assign  data_out[6374] = data_in[1394];
     assign  data_out[6375] = data_in[467];
     assign  data_out[6376] = data_in[69];
     assign  data_out[6377] = data_in[601];
     assign  data_out[6378] = data_in[1345];
     assign  data_out[6379] = data_in[546];
     assign  data_out[6380] = data_in[66];
     assign  data_out[6381] = data_in[1547];
     assign  data_out[6382] = data_in[1156];
     assign  data_out[6383] = data_in[985];
     assign  data_out[6384] = data_in[1591];
     assign  data_out[6385] = data_in[73];
     assign  data_out[6386] = data_in[1130];
     assign  data_out[6387] = data_in[1540];
     assign  data_out[6388] = data_in[794];
     assign  data_out[6389] = data_in[1599];
     assign  data_out[6390] = data_in[825];
     assign  data_out[6391] = data_in[158];
     assign  data_out[6392] = data_in[1001];
     assign  data_out[6393] = data_in[337];
     assign  data_out[6394] = data_in[701];
     assign  data_out[6395] = data_in[368];
     assign  data_out[6396] = data_in[248];
     assign  data_out[6397] = data_in[1367];
     assign  data_out[6398] = data_in[930];
     assign  data_out[6399] = data_in[1213];
     assign  data_out[6400] = data_in[104];
     assign  data_out[6401] = data_in[1279];
     assign  data_out[6402] = data_in[56];
     assign  data_out[6403] = data_in[1522];
     assign  data_out[6404] = data_in[858];
     assign  data_out[6405] = data_in[1121];
     assign  data_out[6406] = data_in[428];
     assign  data_out[6407] = data_in[1075];
     assign  data_out[6408] = data_in[815];
     assign  data_out[6409] = data_in[74];
     assign  data_out[6410] = data_in[624];
     assign  data_out[6411] = data_in[1105];
     assign  data_out[6412] = data_in[1069];
     assign  data_out[6413] = data_in[355];
     assign  data_out[6414] = data_in[816];
     assign  data_out[6415] = data_in[499];
     assign  data_out[6416] = data_in[684];
     assign  data_out[6417] = data_in[1163];
     assign  data_out[6418] = data_in[1271];
     assign  data_out[6419] = data_in[524];
     assign  data_out[6420] = data_in[901];
     assign  data_out[6421] = data_in[90];
     assign  data_out[6422] = data_in[950];
     assign  data_out[6423] = data_in[596];
     assign  data_out[6424] = data_in[1598];
     assign  data_out[6425] = data_in[512];
     assign  data_out[6426] = data_in[578];
     assign  data_out[6427] = data_in[1396];
     assign  data_out[6428] = data_in[1692];
     assign  data_out[6429] = data_in[210];
     assign  data_out[6430] = data_in[1595];
     assign  data_out[6431] = data_in[1299];
     assign  data_out[6432] = data_in[552];
     assign  data_out[6433] = data_in[1200];
     assign  data_out[6434] = data_in[195];
     assign  data_out[6435] = data_in[670];
     assign  data_out[6436] = data_in[0];
     assign  data_out[6437] = data_in[464];
     assign  data_out[6438] = data_in[672];
     assign  data_out[6439] = data_in[45];
     assign  data_out[6440] = data_in[514];
     assign  data_out[6441] = data_in[1573];
     assign  data_out[6442] = data_in[635];
     assign  data_out[6443] = data_in[1508];
     assign  data_out[6444] = data_in[1595];
     assign  data_out[6445] = data_in[1692];
     assign  data_out[6446] = data_in[1693];
     assign  data_out[6447] = data_in[1047];
     assign  data_out[6448] = data_in[1621];
     assign  data_out[6449] = data_in[893];
     assign  data_out[6450] = data_in[1608];
     assign  data_out[6451] = data_in[203];
     assign  data_out[6452] = data_in[246];
     assign  data_out[6453] = data_in[345];
     assign  data_out[6454] = data_in[807];
     assign  data_out[6455] = data_in[585];
     assign  data_out[6456] = data_in[387];
     assign  data_out[6457] = data_in[22];
     assign  data_out[6458] = data_in[1698];
     assign  data_out[6459] = data_in[952];
     assign  data_out[6460] = data_in[784];
     assign  data_out[6461] = data_in[514];
     assign  data_out[6462] = data_in[847];
     assign  data_out[6463] = data_in[156];
     assign  data_out[6464] = data_in[338];
     assign  data_out[6465] = data_in[587];
     assign  data_out[6466] = data_in[859];
     assign  data_out[6467] = data_in[1471];
     assign  data_out[6468] = data_in[47];
     assign  data_out[6469] = data_in[241];
     assign  data_out[6470] = data_in[535];
     assign  data_out[6471] = data_in[847];
     assign  data_out[6472] = data_in[1278];
     assign  data_out[6473] = data_in[917];
     assign  data_out[6474] = data_in[526];
     assign  data_out[6475] = data_in[1294];
     assign  data_out[6476] = data_in[11];
     assign  data_out[6477] = data_in[521];
     assign  data_out[6478] = data_in[323];
     assign  data_out[6479] = data_in[1361];
     assign  data_out[6480] = data_in[1725];
     assign  data_out[6481] = data_in[820];
     assign  data_out[6482] = data_in[1356];
     assign  data_out[6483] = data_in[1641];
     assign  data_out[6484] = data_in[1258];
     assign  data_out[6485] = data_in[690];
     assign  data_out[6486] = data_in[671];
     assign  data_out[6487] = data_in[1462];
     assign  data_out[6488] = data_in[698];
     assign  data_out[6489] = data_in[1409];
     assign  data_out[6490] = data_in[320];
     assign  data_out[6491] = data_in[325];
     assign  data_out[6492] = data_in[991];
     assign  data_out[6493] = data_in[943];
     assign  data_out[6494] = data_in[1404];
     assign  data_out[6495] = data_in[435];
     assign  data_out[6496] = data_in[589];
     assign  data_out[6497] = data_in[1674];
     assign  data_out[6498] = data_in[966];
     assign  data_out[6499] = data_in[693];
     assign  data_out[6500] = data_in[756];
     assign  data_out[6501] = data_in[1612];
     assign  data_out[6502] = data_in[427];
     assign  data_out[6503] = data_in[960];
     assign  data_out[6504] = data_in[739];
     assign  data_out[6505] = data_in[461];
     assign  data_out[6506] = data_in[575];
     assign  data_out[6507] = data_in[51];
     assign  data_out[6508] = data_in[1433];
     assign  data_out[6509] = data_in[932];
     assign  data_out[6510] = data_in[422];
     assign  data_out[6511] = data_in[1093];
     assign  data_out[6512] = data_in[745];
     assign  data_out[6513] = data_in[397];
     assign  data_out[6514] = data_in[863];
     assign  data_out[6515] = data_in[769];
     assign  data_out[6516] = data_in[1023];
     assign  data_out[6517] = data_in[1662];
     assign  data_out[6518] = data_in[1084];
     assign  data_out[6519] = data_in[301];
     assign  data_out[6520] = data_in[1377];
     assign  data_out[6521] = data_in[1656];
     assign  data_out[6522] = data_in[747];
     assign  data_out[6523] = data_in[861];
     assign  data_out[6524] = data_in[439];
     assign  data_out[6525] = data_in[644];
     assign  data_out[6526] = data_in[1070];
     assign  data_out[6527] = data_in[518];
     assign  data_out[6528] = data_in[1407];
     assign  data_out[6529] = data_in[1129];
     assign  data_out[6530] = data_in[566];
     assign  data_out[6531] = data_in[343];
     assign  data_out[6532] = data_in[1723];
     assign  data_out[6533] = data_in[1038];
     assign  data_out[6534] = data_in[1026];
     assign  data_out[6535] = data_in[506];
     assign  data_out[6536] = data_in[687];
     assign  data_out[6537] = data_in[454];
     assign  data_out[6538] = data_in[470];
     assign  data_out[6539] = data_in[880];
     assign  data_out[6540] = data_in[448];
     assign  data_out[6541] = data_in[588];
     assign  data_out[6542] = data_in[792];
     assign  data_out[6543] = data_in[811];
     assign  data_out[6544] = data_in[862];
     assign  data_out[6545] = data_in[425];
     assign  data_out[6546] = data_in[1610];
     assign  data_out[6547] = data_in[484];
     assign  data_out[6548] = data_in[1647];
     assign  data_out[6549] = data_in[831];
     assign  data_out[6550] = data_in[1134];
     assign  data_out[6551] = data_in[276];
     assign  data_out[6552] = data_in[244];
     assign  data_out[6553] = data_in[822];
     assign  data_out[6554] = data_in[1504];
     assign  data_out[6555] = data_in[505];
     assign  data_out[6556] = data_in[544];
     assign  data_out[6557] = data_in[979];
     assign  data_out[6558] = data_in[1373];
     assign  data_out[6559] = data_in[1431];
     assign  data_out[6560] = data_in[140];
     assign  data_out[6561] = data_in[432];
     assign  data_out[6562] = data_in[846];
     assign  data_out[6563] = data_in[754];
     assign  data_out[6564] = data_in[654];
     assign  data_out[6565] = data_in[651];
     assign  data_out[6566] = data_in[1553];
     assign  data_out[6567] = data_in[529];
     assign  data_out[6568] = data_in[156];
     assign  data_out[6569] = data_in[765];
     assign  data_out[6570] = data_in[1032];
     assign  data_out[6571] = data_in[25];
     assign  data_out[6572] = data_in[122];
     assign  data_out[6573] = data_in[1093];
     assign  data_out[6574] = data_in[506];
     assign  data_out[6575] = data_in[274];
     assign  data_out[6576] = data_in[1503];
     assign  data_out[6577] = data_in[1329];
     assign  data_out[6578] = data_in[1030];
     assign  data_out[6579] = data_in[283];
     assign  data_out[6580] = data_in[1618];
     assign  data_out[6581] = data_in[1435];
     assign  data_out[6582] = data_in[175];
     assign  data_out[6583] = data_in[296];
     assign  data_out[6584] = data_in[1005];
     assign  data_out[6585] = data_in[316];
     assign  data_out[6586] = data_in[523];
     assign  data_out[6587] = data_in[708];
     assign  data_out[6588] = data_in[836];
     assign  data_out[6589] = data_in[342];
     assign  data_out[6590] = data_in[656];
     assign  data_out[6591] = data_in[1665];
     assign  data_out[6592] = data_in[21];
     assign  data_out[6593] = data_in[681];
     assign  data_out[6594] = data_in[668];
     assign  data_out[6595] = data_in[585];
     assign  data_out[6596] = data_in[275];
     assign  data_out[6597] = data_in[1341];
     assign  data_out[6598] = data_in[1499];
     assign  data_out[6599] = data_in[1259];
     assign  data_out[6600] = data_in[611];
     assign  data_out[6601] = data_in[888];
     assign  data_out[6602] = data_in[759];
     assign  data_out[6603] = data_in[692];
     assign  data_out[6604] = data_in[1629];
     assign  data_out[6605] = data_in[1084];
     assign  data_out[6606] = data_in[633];
     assign  data_out[6607] = data_in[160];
     assign  data_out[6608] = data_in[1068];
     assign  data_out[6609] = data_in[1427];
     assign  data_out[6610] = data_in[1145];
     assign  data_out[6611] = data_in[1444];
     assign  data_out[6612] = data_in[990];
     assign  data_out[6613] = data_in[287];
     assign  data_out[6614] = data_in[1290];
     assign  data_out[6615] = data_in[187];
     assign  data_out[6616] = data_in[1157];
     assign  data_out[6617] = data_in[1171];
     assign  data_out[6618] = data_in[325];
     assign  data_out[6619] = data_in[1251];
     assign  data_out[6620] = data_in[679];
     assign  data_out[6621] = data_in[1065];
     assign  data_out[6622] = data_in[990];
     assign  data_out[6623] = data_in[630];
     assign  data_out[6624] = data_in[1530];
     assign  data_out[6625] = data_in[868];
     assign  data_out[6626] = data_in[29];
     assign  data_out[6627] = data_in[276];
     assign  data_out[6628] = data_in[1424];
     assign  data_out[6629] = data_in[1028];
     assign  data_out[6630] = data_in[624];
     assign  data_out[6631] = data_in[389];
     assign  data_out[6632] = data_in[764];
     assign  data_out[6633] = data_in[1665];
     assign  data_out[6634] = data_in[1011];
     assign  data_out[6635] = data_in[961];
     assign  data_out[6636] = data_in[798];
     assign  data_out[6637] = data_in[1409];
     assign  data_out[6638] = data_in[787];
     assign  data_out[6639] = data_in[336];
     assign  data_out[6640] = data_in[388];
     assign  data_out[6641] = data_in[386];
     assign  data_out[6642] = data_in[1655];
     assign  data_out[6643] = data_in[115];
     assign  data_out[6644] = data_in[1385];
     assign  data_out[6645] = data_in[1597];
     assign  data_out[6646] = data_in[918];
     assign  data_out[6647] = data_in[694];
     assign  data_out[6648] = data_in[624];
     assign  data_out[6649] = data_in[582];
     assign  data_out[6650] = data_in[1111];
     assign  data_out[6651] = data_in[239];
     assign  data_out[6652] = data_in[1007];
     assign  data_out[6653] = data_in[786];
     assign  data_out[6654] = data_in[1258];
     assign  data_out[6655] = data_in[377];
     assign  data_out[6656] = data_in[665];
     assign  data_out[6657] = data_in[1337];
     assign  data_out[6658] = data_in[60];
     assign  data_out[6659] = data_in[324];
     assign  data_out[6660] = data_in[1320];
     assign  data_out[6661] = data_in[1572];
     assign  data_out[6662] = data_in[688];
     assign  data_out[6663] = data_in[1716];
     assign  data_out[6664] = data_in[28];
     assign  data_out[6665] = data_in[105];
     assign  data_out[6666] = data_in[827];
     assign  data_out[6667] = data_in[691];
     assign  data_out[6668] = data_in[208];
     assign  data_out[6669] = data_in[1676];
     assign  data_out[6670] = data_in[848];
     assign  data_out[6671] = data_in[1586];
     assign  data_out[6672] = data_in[996];
     assign  data_out[6673] = data_in[952];
     assign  data_out[6674] = data_in[1665];
     assign  data_out[6675] = data_in[1136];
     assign  data_out[6676] = data_in[804];
     assign  data_out[6677] = data_in[1423];
     assign  data_out[6678] = data_in[953];
     assign  data_out[6679] = data_in[24];
     assign  data_out[6680] = data_in[37];
     assign  data_out[6681] = data_in[555];
     assign  data_out[6682] = data_in[757];
     assign  data_out[6683] = data_in[1015];
     assign  data_out[6684] = data_in[860];
     assign  data_out[6685] = data_in[1082];
     assign  data_out[6686] = data_in[612];
     assign  data_out[6687] = data_in[425];
     assign  data_out[6688] = data_in[1037];
     assign  data_out[6689] = data_in[325];
     assign  data_out[6690] = data_in[1298];
     assign  data_out[6691] = data_in[1276];
     assign  data_out[6692] = data_in[478];
     assign  data_out[6693] = data_in[139];
     assign  data_out[6694] = data_in[264];
     assign  data_out[6695] = data_in[1314];
     assign  data_out[6696] = data_in[246];
     assign  data_out[6697] = data_in[1477];
     assign  data_out[6698] = data_in[380];
     assign  data_out[6699] = data_in[1526];
     assign  data_out[6700] = data_in[549];
     assign  data_out[6701] = data_in[250];
     assign  data_out[6702] = data_in[970];
     assign  data_out[6703] = data_in[431];
     assign  data_out[6704] = data_in[1671];
     assign  data_out[6705] = data_in[310];
     assign  data_out[6706] = data_in[1416];
     assign  data_out[6707] = data_in[765];
     assign  data_out[6708] = data_in[544];
     assign  data_out[6709] = data_in[1492];
     assign  data_out[6710] = data_in[103];
     assign  data_out[6711] = data_in[757];
     assign  data_out[6712] = data_in[724];
     assign  data_out[6713] = data_in[986];
     assign  data_out[6714] = data_in[3];
     assign  data_out[6715] = data_in[64];
     assign  data_out[6716] = data_in[847];
     assign  data_out[6717] = data_in[562];
     assign  data_out[6718] = data_in[204];
     assign  data_out[6719] = data_in[1206];
     assign  data_out[6720] = data_in[48];
     assign  data_out[6721] = data_in[875];
     assign  data_out[6722] = data_in[230];
     assign  data_out[6723] = data_in[279];
     assign  data_out[6724] = data_in[976];
     assign  data_out[6725] = data_in[1290];
     assign  data_out[6726] = data_in[1649];
     assign  data_out[6727] = data_in[1357];
     assign  data_out[6728] = data_in[507];
     assign  data_out[6729] = data_in[307];
     assign  data_out[6730] = data_in[976];
     assign  data_out[6731] = data_in[1705];
     assign  data_out[6732] = data_in[618];
     assign  data_out[6733] = data_in[1166];
     assign  data_out[6734] = data_in[1576];
     assign  data_out[6735] = data_in[1219];
     assign  data_out[6736] = data_in[165];
     assign  data_out[6737] = data_in[450];
     assign  data_out[6738] = data_in[555];
     assign  data_out[6739] = data_in[495];
     assign  data_out[6740] = data_in[11];
     assign  data_out[6741] = data_in[559];
     assign  data_out[6742] = data_in[802];
     assign  data_out[6743] = data_in[1208];
     assign  data_out[6744] = data_in[1262];
     assign  data_out[6745] = data_in[1396];
     assign  data_out[6746] = data_in[723];
     assign  data_out[6747] = data_in[838];
     assign  data_out[6748] = data_in[1413];
     assign  data_out[6749] = data_in[49];
     assign  data_out[6750] = data_in[1455];
     assign  data_out[6751] = data_in[617];
     assign  data_out[6752] = data_in[986];
     assign  data_out[6753] = data_in[467];
     assign  data_out[6754] = data_in[1389];
     assign  data_out[6755] = data_in[1446];
     assign  data_out[6756] = data_in[1276];
     assign  data_out[6757] = data_in[1432];
     assign  data_out[6758] = data_in[501];
     assign  data_out[6759] = data_in[1483];
     assign  data_out[6760] = data_in[602];
     assign  data_out[6761] = data_in[1109];
     assign  data_out[6762] = data_in[1599];
     assign  data_out[6763] = data_in[1251];
     assign  data_out[6764] = data_in[781];
     assign  data_out[6765] = data_in[305];
     assign  data_out[6766] = data_in[1628];
     assign  data_out[6767] = data_in[576];
     assign  data_out[6768] = data_in[116];
     assign  data_out[6769] = data_in[1255];
     assign  data_out[6770] = data_in[1588];
     assign  data_out[6771] = data_in[146];
     assign  data_out[6772] = data_in[178];
     assign  data_out[6773] = data_in[1324];
     assign  data_out[6774] = data_in[569];
     assign  data_out[6775] = data_in[609];
     assign  data_out[6776] = data_in[930];
     assign  data_out[6777] = data_in[924];
     assign  data_out[6778] = data_in[740];
     assign  data_out[6779] = data_in[1659];
     assign  data_out[6780] = data_in[1115];
     assign  data_out[6781] = data_in[849];
     assign  data_out[6782] = data_in[873];
     assign  data_out[6783] = data_in[928];
     assign  data_out[6784] = data_in[928];
     assign  data_out[6785] = data_in[1389];
     assign  data_out[6786] = data_in[75];
     assign  data_out[6787] = data_in[305];
     assign  data_out[6788] = data_in[1405];
     assign  data_out[6789] = data_in[916];
     assign  data_out[6790] = data_in[1387];
     assign  data_out[6791] = data_in[521];
     assign  data_out[6792] = data_in[1024];
     assign  data_out[6793] = data_in[1107];
     assign  data_out[6794] = data_in[641];
     assign  data_out[6795] = data_in[240];
     assign  data_out[6796] = data_in[1240];
     assign  data_out[6797] = data_in[947];
     assign  data_out[6798] = data_in[362];
     assign  data_out[6799] = data_in[1234];
     assign  data_out[6800] = data_in[682];
     assign  data_out[6801] = data_in[503];
     assign  data_out[6802] = data_in[1246];
     assign  data_out[6803] = data_in[1319];
     assign  data_out[6804] = data_in[127];
     assign  data_out[6805] = data_in[59];
     assign  data_out[6806] = data_in[651];
     assign  data_out[6807] = data_in[839];
     assign  data_out[6808] = data_in[1435];
     assign  data_out[6809] = data_in[63];
     assign  data_out[6810] = data_in[739];
     assign  data_out[6811] = data_in[901];
     assign  data_out[6812] = data_in[75];
     assign  data_out[6813] = data_in[1302];
     assign  data_out[6814] = data_in[419];
     assign  data_out[6815] = data_in[143];
     assign  data_out[6816] = data_in[1111];
     assign  data_out[6817] = data_in[366];
     assign  data_out[6818] = data_in[1360];
     assign  data_out[6819] = data_in[1075];
     assign  data_out[6820] = data_in[1228];
     assign  data_out[6821] = data_in[576];
     assign  data_out[6822] = data_in[503];
     assign  data_out[6823] = data_in[1671];
     assign  data_out[6824] = data_in[1242];
     assign  data_out[6825] = data_in[604];
     assign  data_out[6826] = data_in[1082];
     assign  data_out[6827] = data_in[531];
     assign  data_out[6828] = data_in[310];
     assign  data_out[6829] = data_in[1673];
     assign  data_out[6830] = data_in[738];
     assign  data_out[6831] = data_in[1653];
     assign  data_out[6832] = data_in[1722];
     assign  data_out[6833] = data_in[779];
     assign  data_out[6834] = data_in[850];
     assign  data_out[6835] = data_in[487];
     assign  data_out[6836] = data_in[507];
     assign  data_out[6837] = data_in[435];
     assign  data_out[6838] = data_in[834];
     assign  data_out[6839] = data_in[1238];
     assign  data_out[6840] = data_in[3];
     assign  data_out[6841] = data_in[655];
     assign  data_out[6842] = data_in[813];
     assign  data_out[6843] = data_in[451];
     assign  data_out[6844] = data_in[1708];
     assign  data_out[6845] = data_in[231];
     assign  data_out[6846] = data_in[597];
     assign  data_out[6847] = data_in[640];
     assign  data_out[6848] = data_in[15];
     assign  data_out[6849] = data_in[656];
     assign  data_out[6850] = data_in[1084];
     assign  data_out[6851] = data_in[1120];
     assign  data_out[6852] = data_in[450];
     assign  data_out[6853] = data_in[7];
     assign  data_out[6854] = data_in[1228];
     assign  data_out[6855] = data_in[413];
     assign  data_out[6856] = data_in[1423];
     assign  data_out[6857] = data_in[1252];
     assign  data_out[6858] = data_in[123];
     assign  data_out[6859] = data_in[580];
     assign  data_out[6860] = data_in[1324];
     assign  data_out[6861] = data_in[1550];
     assign  data_out[6862] = data_in[802];
     assign  data_out[6863] = data_in[1216];
     assign  data_out[6864] = data_in[339];
     assign  data_out[6865] = data_in[832];
     assign  data_out[6866] = data_in[1124];
     assign  data_out[6867] = data_in[1087];
     assign  data_out[6868] = data_in[76];
     assign  data_out[6869] = data_in[1425];
     assign  data_out[6870] = data_in[1178];
     assign  data_out[6871] = data_in[338];
     assign  data_out[6872] = data_in[1475];
     assign  data_out[6873] = data_in[707];
     assign  data_out[6874] = data_in[459];
     assign  data_out[6875] = data_in[518];
     assign  data_out[6876] = data_in[628];
     assign  data_out[6877] = data_in[404];
     assign  data_out[6878] = data_in[450];
     assign  data_out[6879] = data_in[532];
     assign  data_out[6880] = data_in[281];
     assign  data_out[6881] = data_in[1685];
     assign  data_out[6882] = data_in[1402];
     assign  data_out[6883] = data_in[1313];
     assign  data_out[6884] = data_in[339];
     assign  data_out[6885] = data_in[1017];
     assign  data_out[6886] = data_in[300];
     assign  data_out[6887] = data_in[57];
     assign  data_out[6888] = data_in[711];
     assign  data_out[6889] = data_in[870];
     assign  data_out[6890] = data_in[1287];
     assign  data_out[6891] = data_in[625];
     assign  data_out[6892] = data_in[543];
     assign  data_out[6893] = data_in[131];
     assign  data_out[6894] = data_in[598];
     assign  data_out[6895] = data_in[222];
     assign  data_out[6896] = data_in[1252];
     assign  data_out[6897] = data_in[763];
     assign  data_out[6898] = data_in[474];
     assign  data_out[6899] = data_in[1428];
     assign  data_out[6900] = data_in[886];
     assign  data_out[6901] = data_in[759];
     assign  data_out[6902] = data_in[281];
     assign  data_out[6903] = data_in[1043];
     assign  data_out[6904] = data_in[1025];
     assign  data_out[6905] = data_in[1304];
     assign  data_out[6906] = data_in[308];
     assign  data_out[6907] = data_in[1370];
     assign  data_out[6908] = data_in[1656];
     assign  data_out[6909] = data_in[1616];
     assign  data_out[6910] = data_in[1024];
     assign  data_out[6911] = data_in[576];
     assign  data_out[6912] = data_in[65];
     assign  data_out[6913] = data_in[772];
     assign  data_out[6914] = data_in[424];
     assign  data_out[6915] = data_in[852];
     assign  data_out[6916] = data_in[275];
     assign  data_out[6917] = data_in[715];
     assign  data_out[6918] = data_in[1636];
     assign  data_out[6919] = data_in[1374];
     assign  data_out[6920] = data_in[680];
     assign  data_out[6921] = data_in[355];
     assign  data_out[6922] = data_in[587];
     assign  data_out[6923] = data_in[959];
     assign  data_out[6924] = data_in[979];
     assign  data_out[6925] = data_in[912];
     assign  data_out[6926] = data_in[441];
     assign  data_out[6927] = data_in[1615];
     assign  data_out[6928] = data_in[1243];
     assign  data_out[6929] = data_in[293];
     assign  data_out[6930] = data_in[165];
     assign  data_out[6931] = data_in[1599];
     assign  data_out[6932] = data_in[1372];
     assign  data_out[6933] = data_in[111];
     assign  data_out[6934] = data_in[470];
     assign  data_out[6935] = data_in[263];
     assign  data_out[6936] = data_in[1441];
     assign  data_out[6937] = data_in[1425];
     assign  data_out[6938] = data_in[399];
     assign  data_out[6939] = data_in[1596];
     assign  data_out[6940] = data_in[808];
     assign  data_out[6941] = data_in[693];
     assign  data_out[6942] = data_in[175];
     assign  data_out[6943] = data_in[720];
     assign  data_out[6944] = data_in[1685];
     assign  data_out[6945] = data_in[41];
     assign  data_out[6946] = data_in[845];
     assign  data_out[6947] = data_in[719];
     assign  data_out[6948] = data_in[1203];
     assign  data_out[6949] = data_in[152];
     assign  data_out[6950] = data_in[786];
     assign  data_out[6951] = data_in[870];
     assign  data_out[6952] = data_in[148];
     assign  data_out[6953] = data_in[224];
     assign  data_out[6954] = data_in[356];
     assign  data_out[6955] = data_in[199];
     assign  data_out[6956] = data_in[296];
     assign  data_out[6957] = data_in[962];
     assign  data_out[6958] = data_in[915];
     assign  data_out[6959] = data_in[620];
     assign  data_out[6960] = data_in[1249];
     assign  data_out[6961] = data_in[494];
     assign  data_out[6962] = data_in[870];
     assign  data_out[6963] = data_in[16];
     assign  data_out[6964] = data_in[1535];
     assign  data_out[6965] = data_in[1639];
     assign  data_out[6966] = data_in[883];
     assign  data_out[6967] = data_in[1012];
     assign  data_out[6968] = data_in[1029];
     assign  data_out[6969] = data_in[1401];
     assign  data_out[6970] = data_in[173];
     assign  data_out[6971] = data_in[1571];
     assign  data_out[6972] = data_in[854];
     assign  data_out[6973] = data_in[132];
     assign  data_out[6974] = data_in[1214];
     assign  data_out[6975] = data_in[104];
     assign  data_out[6976] = data_in[1244];
     assign  data_out[6977] = data_in[1240];
     assign  data_out[6978] = data_in[1312];
     assign  data_out[6979] = data_in[220];
     assign  data_out[6980] = data_in[451];
     assign  data_out[6981] = data_in[868];
     assign  data_out[6982] = data_in[480];
     assign  data_out[6983] = data_in[1153];
     assign  data_out[6984] = data_in[364];
     assign  data_out[6985] = data_in[619];
     assign  data_out[6986] = data_in[605];
     assign  data_out[6987] = data_in[475];
     assign  data_out[6988] = data_in[1182];
     assign  data_out[6989] = data_in[1291];
     assign  data_out[6990] = data_in[1147];
     assign  data_out[6991] = data_in[288];
     assign  data_out[6992] = data_in[1184];
     assign  data_out[6993] = data_in[333];
     assign  data_out[6994] = data_in[937];
     assign  data_out[6995] = data_in[333];
     assign  data_out[6996] = data_in[1212];
     assign  data_out[6997] = data_in[1076];
     assign  data_out[6998] = data_in[932];
     assign  data_out[6999] = data_in[307];
     assign  data_out[7000] = data_in[525];
     assign  data_out[7001] = data_in[1183];
     assign  data_out[7002] = data_in[210];
     assign  data_out[7003] = data_in[1722];
     assign  data_out[7004] = data_in[943];
     assign  data_out[7005] = data_in[1186];
     assign  data_out[7006] = data_in[810];
     assign  data_out[7007] = data_in[510];
     assign  data_out[7008] = data_in[736];
     assign  data_out[7009] = data_in[554];
     assign  data_out[7010] = data_in[1607];
     assign  data_out[7011] = data_in[443];
     assign  data_out[7012] = data_in[369];
     assign  data_out[7013] = data_in[1428];
     assign  data_out[7014] = data_in[264];
     assign  data_out[7015] = data_in[565];
     assign  data_out[7016] = data_in[1552];
     assign  data_out[7017] = data_in[1301];
     assign  data_out[7018] = data_in[750];
     assign  data_out[7019] = data_in[513];
     assign  data_out[7020] = data_in[977];
     assign  data_out[7021] = data_in[1670];
     assign  data_out[7022] = data_in[532];
     assign  data_out[7023] = data_in[1135];
     assign  data_out[7024] = data_in[1663];
     assign  data_out[7025] = data_in[125];
     assign  data_out[7026] = data_in[1580];
     assign  data_out[7027] = data_in[1073];
     assign  data_out[7028] = data_in[80];
     assign  data_out[7029] = data_in[1552];
     assign  data_out[7030] = data_in[296];
     assign  data_out[7031] = data_in[1269];
     assign  data_out[7032] = data_in[1368];
     assign  data_out[7033] = data_in[344];
     assign  data_out[7034] = data_in[492];
     assign  data_out[7035] = data_in[802];
     assign  data_out[7036] = data_in[62];
     assign  data_out[7037] = data_in[413];
     assign  data_out[7038] = data_in[1088];
     assign  data_out[7039] = data_in[1185];
     assign  data_out[7040] = data_in[1126];
     assign  data_out[7041] = data_in[701];
     assign  data_out[7042] = data_in[916];
     assign  data_out[7043] = data_in[805];
     assign  data_out[7044] = data_in[1415];
     assign  data_out[7045] = data_in[888];
     assign  data_out[7046] = data_in[1679];
     assign  data_out[7047] = data_in[92];
     assign  data_out[7048] = data_in[1181];
     assign  data_out[7049] = data_in[1656];
     assign  data_out[7050] = data_in[1341];
     assign  data_out[7051] = data_in[821];
     assign  data_out[7052] = data_in[315];
     assign  data_out[7053] = data_in[625];
     assign  data_out[7054] = data_in[465];
     assign  data_out[7055] = data_in[1139];
     assign  data_out[7056] = data_in[545];
     assign  data_out[7057] = data_in[1536];
     assign  data_out[7058] = data_in[1689];
     assign  data_out[7059] = data_in[816];
     assign  data_out[7060] = data_in[1110];
     assign  data_out[7061] = data_in[1501];
     assign  data_out[7062] = data_in[653];
     assign  data_out[7063] = data_in[1025];
     assign  data_out[7064] = data_in[514];
     assign  data_out[7065] = data_in[1536];
     assign  data_out[7066] = data_in[410];
     assign  data_out[7067] = data_in[1074];
     assign  data_out[7068] = data_in[495];
     assign  data_out[7069] = data_in[38];
     assign  data_out[7070] = data_in[984];
     assign  data_out[7071] = data_in[564];
     assign  data_out[7072] = data_in[625];
     assign  data_out[7073] = data_in[566];
     assign  data_out[7074] = data_in[1290];
     assign  data_out[7075] = data_in[774];
     assign  data_out[7076] = data_in[430];
     assign  data_out[7077] = data_in[515];
     assign  data_out[7078] = data_in[1356];
     assign  data_out[7079] = data_in[1640];
     assign  data_out[7080] = data_in[878];
     assign  data_out[7081] = data_in[689];
     assign  data_out[7082] = data_in[607];
     assign  data_out[7083] = data_in[233];
     assign  data_out[7084] = data_in[1399];
     assign  data_out[7085] = data_in[627];
     assign  data_out[7086] = data_in[882];
     assign  data_out[7087] = data_in[922];
     assign  data_out[7088] = data_in[1577];
     assign  data_out[7089] = data_in[671];
     assign  data_out[7090] = data_in[1287];
     assign  data_out[7091] = data_in[1647];
     assign  data_out[7092] = data_in[198];
     assign  data_out[7093] = data_in[1568];
     assign  data_out[7094] = data_in[494];
     assign  data_out[7095] = data_in[1076];
     assign  data_out[7096] = data_in[804];
     assign  data_out[7097] = data_in[120];
     assign  data_out[7098] = data_in[486];
     assign  data_out[7099] = data_in[1400];
     assign  data_out[7100] = data_in[904];
     assign  data_out[7101] = data_in[1046];
     assign  data_out[7102] = data_in[1434];
     assign  data_out[7103] = data_in[1459];
     assign  data_out[7104] = data_in[1603];
     assign  data_out[7105] = data_in[386];
     assign  data_out[7106] = data_in[726];
     assign  data_out[7107] = data_in[1600];
     assign  data_out[7108] = data_in[1008];
     assign  data_out[7109] = data_in[334];
     assign  data_out[7110] = data_in[1376];
     assign  data_out[7111] = data_in[1122];
     assign  data_out[7112] = data_in[1244];
     assign  data_out[7113] = data_in[486];
     assign  data_out[7114] = data_in[1367];
     assign  data_out[7115] = data_in[1094];
     assign  data_out[7116] = data_in[1083];
     assign  data_out[7117] = data_in[1173];
     assign  data_out[7118] = data_in[261];
     assign  data_out[7119] = data_in[297];
     assign  data_out[7120] = data_in[569];
     assign  data_out[7121] = data_in[167];
     assign  data_out[7122] = data_in[1532];
     assign  data_out[7123] = data_in[526];
     assign  data_out[7124] = data_in[1718];
     assign  data_out[7125] = data_in[1159];
     assign  data_out[7126] = data_in[309];
     assign  data_out[7127] = data_in[384];
     assign  data_out[7128] = data_in[600];
     assign  data_out[7129] = data_in[1448];
     assign  data_out[7130] = data_in[650];
     assign  data_out[7131] = data_in[696];
     assign  data_out[7132] = data_in[1520];
     assign  data_out[7133] = data_in[1451];
     assign  data_out[7134] = data_in[186];
     assign  data_out[7135] = data_in[686];
     assign  data_out[7136] = data_in[220];
     assign  data_out[7137] = data_in[15];
     assign  data_out[7138] = data_in[86];
     assign  data_out[7139] = data_in[1133];
     assign  data_out[7140] = data_in[1392];
     assign  data_out[7141] = data_in[858];
     assign  data_out[7142] = data_in[636];
     assign  data_out[7143] = data_in[550];
     assign  data_out[7144] = data_in[126];
     assign  data_out[7145] = data_in[1024];
     assign  data_out[7146] = data_in[662];
     assign  data_out[7147] = data_in[618];
     assign  data_out[7148] = data_in[1244];
     assign  data_out[7149] = data_in[521];
     assign  data_out[7150] = data_in[808];
     assign  data_out[7151] = data_in[1723];
     assign  data_out[7152] = data_in[943];
     assign  data_out[7153] = data_in[556];
     assign  data_out[7154] = data_in[1261];
     assign  data_out[7155] = data_in[1377];
     assign  data_out[7156] = data_in[1243];
     assign  data_out[7157] = data_in[165];
     assign  data_out[7158] = data_in[858];
     assign  data_out[7159] = data_in[557];
     assign  data_out[7160] = data_in[690];
     assign  data_out[7161] = data_in[125];
     assign  data_out[7162] = data_in[238];
     assign  data_out[7163] = data_in[1386];
     assign  data_out[7164] = data_in[682];
     assign  data_out[7165] = data_in[1480];
     assign  data_out[7166] = data_in[445];
     assign  data_out[7167] = data_in[1161];
     assign  data_out[7168] = data_in[250];
     assign  data_out[7169] = data_in[663];
     assign  data_out[7170] = data_in[1364];
     assign  data_out[7171] = data_in[731];
     assign  data_out[7172] = data_in[1394];
     assign  data_out[7173] = data_in[1356];
     assign  data_out[7174] = data_in[32];
     assign  data_out[7175] = data_in[1128];
     assign  data_out[7176] = data_in[1258];
     assign  data_out[7177] = data_in[177];
     assign  data_out[7178] = data_in[121];
     assign  data_out[7179] = data_in[1258];
     assign  data_out[7180] = data_in[141];
     assign  data_out[7181] = data_in[870];
     assign  data_out[7182] = data_in[1539];
     assign  data_out[7183] = data_in[1667];
     assign  data_out[7184] = data_in[1639];
     assign  data_out[7185] = data_in[264];
     assign  data_out[7186] = data_in[444];
     assign  data_out[7187] = data_in[1264];
     assign  data_out[7188] = data_in[1095];
     assign  data_out[7189] = data_in[689];
     assign  data_out[7190] = data_in[1443];
     assign  data_out[7191] = data_in[667];
     assign  data_out[7192] = data_in[841];
     assign  data_out[7193] = data_in[747];
     assign  data_out[7194] = data_in[1447];
     assign  data_out[7195] = data_in[766];
     assign  data_out[7196] = data_in[25];
     assign  data_out[7197] = data_in[121];
     assign  data_out[7198] = data_in[500];
     assign  data_out[7199] = data_in[1538];
     assign  data_out[7200] = data_in[983];
     assign  data_out[7201] = data_in[1428];
     assign  data_out[7202] = data_in[779];
     assign  data_out[7203] = data_in[79];
     assign  data_out[7204] = data_in[664];
     assign  data_out[7205] = data_in[1583];
     assign  data_out[7206] = data_in[727];
     assign  data_out[7207] = data_in[1522];
     assign  data_out[7208] = data_in[435];
     assign  data_out[7209] = data_in[622];
     assign  data_out[7210] = data_in[781];
     assign  data_out[7211] = data_in[336];
     assign  data_out[7212] = data_in[1054];
     assign  data_out[7213] = data_in[1451];
     assign  data_out[7214] = data_in[16];
     assign  data_out[7215] = data_in[966];
     assign  data_out[7216] = data_in[572];
     assign  data_out[7217] = data_in[796];
     assign  data_out[7218] = data_in[184];
     assign  data_out[7219] = data_in[764];
     assign  data_out[7220] = data_in[1707];
     assign  data_out[7221] = data_in[140];
     assign  data_out[7222] = data_in[1636];
     assign  data_out[7223] = data_in[702];
     assign  data_out[7224] = data_in[1516];
     assign  data_out[7225] = data_in[618];
     assign  data_out[7226] = data_in[697];
     assign  data_out[7227] = data_in[1369];
     assign  data_out[7228] = data_in[1020];
     assign  data_out[7229] = data_in[302];
     assign  data_out[7230] = data_in[637];
     assign  data_out[7231] = data_in[1386];
     assign  data_out[7232] = data_in[687];
     assign  data_out[7233] = data_in[1035];
     assign  data_out[7234] = data_in[864];
     assign  data_out[7235] = data_in[645];
     assign  data_out[7236] = data_in[417];
     assign  data_out[7237] = data_in[54];
     assign  data_out[7238] = data_in[702];
     assign  data_out[7239] = data_in[1316];
     assign  data_out[7240] = data_in[1066];
     assign  data_out[7241] = data_in[1204];
     assign  data_out[7242] = data_in[1357];
     assign  data_out[7243] = data_in[412];
     assign  data_out[7244] = data_in[191];
     assign  data_out[7245] = data_in[249];
     assign  data_out[7246] = data_in[981];
     assign  data_out[7247] = data_in[1377];
     assign  data_out[7248] = data_in[1543];
     assign  data_out[7249] = data_in[1549];
     assign  data_out[7250] = data_in[992];
     assign  data_out[7251] = data_in[507];
     assign  data_out[7252] = data_in[1621];
     assign  data_out[7253] = data_in[1593];
     assign  data_out[7254] = data_in[1278];
     assign  data_out[7255] = data_in[1568];
     assign  data_out[7256] = data_in[430];
     assign  data_out[7257] = data_in[124];
     assign  data_out[7258] = data_in[726];
     assign  data_out[7259] = data_in[599];
     assign  data_out[7260] = data_in[1522];
     assign  data_out[7261] = data_in[252];
     assign  data_out[7262] = data_in[1414];
     assign  data_out[7263] = data_in[1194];
     assign  data_out[7264] = data_in[55];
     assign  data_out[7265] = data_in[1285];
     assign  data_out[7266] = data_in[106];
     assign  data_out[7267] = data_in[492];
     assign  data_out[7268] = data_in[1707];
     assign  data_out[7269] = data_in[952];
     assign  data_out[7270] = data_in[1660];
     assign  data_out[7271] = data_in[1011];
     assign  data_out[7272] = data_in[350];
     assign  data_out[7273] = data_in[390];
     assign  data_out[7274] = data_in[1698];
     assign  data_out[7275] = data_in[644];
     assign  data_out[7276] = data_in[509];
     assign  data_out[7277] = data_in[922];
     assign  data_out[7278] = data_in[805];
     assign  data_out[7279] = data_in[393];
     assign  data_out[7280] = data_in[415];
     assign  data_out[7281] = data_in[1543];
     assign  data_out[7282] = data_in[1056];
     assign  data_out[7283] = data_in[1176];
     assign  data_out[7284] = data_in[945];
     assign  data_out[7285] = data_in[1700];
     assign  data_out[7286] = data_in[482];
     assign  data_out[7287] = data_in[1634];
     assign  data_out[7288] = data_in[1179];
     assign  data_out[7289] = data_in[996];
     assign  data_out[7290] = data_in[221];
     assign  data_out[7291] = data_in[1097];
     assign  data_out[7292] = data_in[950];
     assign  data_out[7293] = data_in[416];
     assign  data_out[7294] = data_in[202];
     assign  data_out[7295] = data_in[640];
     assign  data_out[7296] = data_in[487];
     assign  data_out[7297] = data_in[144];
     assign  data_out[7298] = data_in[1578];
     assign  data_out[7299] = data_in[1196];
     assign  data_out[7300] = data_in[241];
     assign  data_out[7301] = data_in[307];
     assign  data_out[7302] = data_in[392];
     assign  data_out[7303] = data_in[299];
     assign  data_out[7304] = data_in[1372];
     assign  data_out[7305] = data_in[1452];
     assign  data_out[7306] = data_in[1058];
     assign  data_out[7307] = data_in[245];
     assign  data_out[7308] = data_in[1346];
     assign  data_out[7309] = data_in[702];
     assign  data_out[7310] = data_in[1316];
     assign  data_out[7311] = data_in[1606];
     assign  data_out[7312] = data_in[664];
     assign  data_out[7313] = data_in[1149];
     assign  data_out[7314] = data_in[1425];
     assign  data_out[7315] = data_in[55];
     assign  data_out[7316] = data_in[1354];
     assign  data_out[7317] = data_in[1053];
     assign  data_out[7318] = data_in[1356];
     assign  data_out[7319] = data_in[187];
     assign  data_out[7320] = data_in[1153];
     assign  data_out[7321] = data_in[1136];
     assign  data_out[7322] = data_in[731];
     assign  data_out[7323] = data_in[375];
     assign  data_out[7324] = data_in[291];
     assign  data_out[7325] = data_in[1725];
     assign  data_out[7326] = data_in[1555];
     assign  data_out[7327] = data_in[320];
     assign  data_out[7328] = data_in[626];
     assign  data_out[7329] = data_in[386];
     assign  data_out[7330] = data_in[851];
     assign  data_out[7331] = data_in[930];
     assign  data_out[7332] = data_in[204];
     assign  data_out[7333] = data_in[1547];
     assign  data_out[7334] = data_in[872];
     assign  data_out[7335] = data_in[1517];
     assign  data_out[7336] = data_in[1007];
     assign  data_out[7337] = data_in[373];
     assign  data_out[7338] = data_in[1553];
     assign  data_out[7339] = data_in[210];
     assign  data_out[7340] = data_in[151];
     assign  data_out[7341] = data_in[761];
     assign  data_out[7342] = data_in[1153];
     assign  data_out[7343] = data_in[887];
     assign  data_out[7344] = data_in[1285];
     assign  data_out[7345] = data_in[357];
     assign  data_out[7346] = data_in[828];
     assign  data_out[7347] = data_in[1389];
     assign  data_out[7348] = data_in[905];
     assign  data_out[7349] = data_in[730];
     assign  data_out[7350] = data_in[1097];
     assign  data_out[7351] = data_in[888];
     assign  data_out[7352] = data_in[169];
     assign  data_out[7353] = data_in[1519];
     assign  data_out[7354] = data_in[1484];
     assign  data_out[7355] = data_in[1181];
     assign  data_out[7356] = data_in[367];
     assign  data_out[7357] = data_in[410];
     assign  data_out[7358] = data_in[1656];
     assign  data_out[7359] = data_in[19];
     assign  data_out[7360] = data_in[1546];
     assign  data_out[7361] = data_in[949];
     assign  data_out[7362] = data_in[1538];
     assign  data_out[7363] = data_in[1376];
     assign  data_out[7364] = data_in[436];
     assign  data_out[7365] = data_in[1674];
     assign  data_out[7366] = data_in[429];
     assign  data_out[7367] = data_in[1009];
     assign  data_out[7368] = data_in[289];
     assign  data_out[7369] = data_in[1397];
     assign  data_out[7370] = data_in[1250];
     assign  data_out[7371] = data_in[1587];
     assign  data_out[7372] = data_in[1124];
     assign  data_out[7373] = data_in[1032];
     assign  data_out[7374] = data_in[956];
     assign  data_out[7375] = data_in[209];
     assign  data_out[7376] = data_in[247];
     assign  data_out[7377] = data_in[511];
     assign  data_out[7378] = data_in[856];
     assign  data_out[7379] = data_in[841];
     assign  data_out[7380] = data_in[947];
     assign  data_out[7381] = data_in[569];
     assign  data_out[7382] = data_in[627];
     assign  data_out[7383] = data_in[1403];
     assign  data_out[7384] = data_in[475];
     assign  data_out[7385] = data_in[1018];
     assign  data_out[7386] = data_in[1113];
     assign  data_out[7387] = data_in[1135];
     assign  data_out[7388] = data_in[114];
     assign  data_out[7389] = data_in[102];
     assign  data_out[7390] = data_in[415];
     assign  data_out[7391] = data_in[443];
     assign  data_out[7392] = data_in[1565];
     assign  data_out[7393] = data_in[394];
     assign  data_out[7394] = data_in[1478];
     assign  data_out[7395] = data_in[816];
     assign  data_out[7396] = data_in[1342];
     assign  data_out[7397] = data_in[1631];
     assign  data_out[7398] = data_in[121];
     assign  data_out[7399] = data_in[1220];
     assign  data_out[7400] = data_in[953];
     assign  data_out[7401] = data_in[1478];
     assign  data_out[7402] = data_in[1078];
     assign  data_out[7403] = data_in[293];
     assign  data_out[7404] = data_in[1389];
     assign  data_out[7405] = data_in[202];
     assign  data_out[7406] = data_in[1631];
     assign  data_out[7407] = data_in[736];
     assign  data_out[7408] = data_in[1404];
     assign  data_out[7409] = data_in[846];
     assign  data_out[7410] = data_in[775];
     assign  data_out[7411] = data_in[1040];
     assign  data_out[7412] = data_in[942];
     assign  data_out[7413] = data_in[893];
     assign  data_out[7414] = data_in[1138];
     assign  data_out[7415] = data_in[316];
     assign  data_out[7416] = data_in[1565];
     assign  data_out[7417] = data_in[1582];
     assign  data_out[7418] = data_in[1115];
     assign  data_out[7419] = data_in[1367];
     assign  data_out[7420] = data_in[30];
     assign  data_out[7421] = data_in[1460];
     assign  data_out[7422] = data_in[1466];
     assign  data_out[7423] = data_in[1485];
     assign  data_out[7424] = data_in[1434];
     assign  data_out[7425] = data_in[361];
     assign  data_out[7426] = data_in[1369];
     assign  data_out[7427] = data_in[1040];
     assign  data_out[7428] = data_in[1438];
     assign  data_out[7429] = data_in[1119];
     assign  data_out[7430] = data_in[1275];
     assign  data_out[7431] = data_in[331];
     assign  data_out[7432] = data_in[252];
     assign  data_out[7433] = data_in[650];
     assign  data_out[7434] = data_in[1371];
     assign  data_out[7435] = data_in[942];
     assign  data_out[7436] = data_in[1366];
     assign  data_out[7437] = data_in[903];
     assign  data_out[7438] = data_in[902];
     assign  data_out[7439] = data_in[1092];
     assign  data_out[7440] = data_in[672];
     assign  data_out[7441] = data_in[220];
     assign  data_out[7442] = data_in[988];
     assign  data_out[7443] = data_in[1211];
     assign  data_out[7444] = data_in[187];
     assign  data_out[7445] = data_in[782];
     assign  data_out[7446] = data_in[634];
     assign  data_out[7447] = data_in[586];
     assign  data_out[7448] = data_in[181];
     assign  data_out[7449] = data_in[1327];
     assign  data_out[7450] = data_in[663];
     assign  data_out[7451] = data_in[1331];
     assign  data_out[7452] = data_in[455];
     assign  data_out[7453] = data_in[448];
     assign  data_out[7454] = data_in[75];
     assign  data_out[7455] = data_in[501];
     assign  data_out[7456] = data_in[877];
     assign  data_out[7457] = data_in[382];
     assign  data_out[7458] = data_in[1316];
     assign  data_out[7459] = data_in[437];
     assign  data_out[7460] = data_in[804];
     assign  data_out[7461] = data_in[327];
     assign  data_out[7462] = data_in[304];
     assign  data_out[7463] = data_in[894];
     assign  data_out[7464] = data_in[1325];
     assign  data_out[7465] = data_in[294];
     assign  data_out[7466] = data_in[142];
     assign  data_out[7467] = data_in[1287];
     assign  data_out[7468] = data_in[1310];
     assign  data_out[7469] = data_in[1069];
     assign  data_out[7470] = data_in[216];
     assign  data_out[7471] = data_in[821];
     assign  data_out[7472] = data_in[1584];
     assign  data_out[7473] = data_in[569];
     assign  data_out[7474] = data_in[1303];
     assign  data_out[7475] = data_in[633];
     assign  data_out[7476] = data_in[1276];
     assign  data_out[7477] = data_in[1530];
     assign  data_out[7478] = data_in[849];
     assign  data_out[7479] = data_in[906];
     assign  data_out[7480] = data_in[675];
     assign  data_out[7481] = data_in[1445];
     assign  data_out[7482] = data_in[63];
     assign  data_out[7483] = data_in[538];
     assign  data_out[7484] = data_in[1563];
     assign  data_out[7485] = data_in[425];
     assign  data_out[7486] = data_in[417];
     assign  data_out[7487] = data_in[949];
     assign  data_out[7488] = data_in[319];
     assign  data_out[7489] = data_in[1340];
     assign  data_out[7490] = data_in[831];
     assign  data_out[7491] = data_in[906];
     assign  data_out[7492] = data_in[1090];
     assign  data_out[7493] = data_in[1657];
     assign  data_out[7494] = data_in[801];
     assign  data_out[7495] = data_in[1198];
     assign  data_out[7496] = data_in[1101];
     assign  data_out[7497] = data_in[1415];
     assign  data_out[7498] = data_in[1721];
     assign  data_out[7499] = data_in[866];
     assign  data_out[7500] = data_in[1318];
     assign  data_out[7501] = data_in[847];
     assign  data_out[7502] = data_in[1293];
     assign  data_out[7503] = data_in[383];
     assign  data_out[7504] = data_in[1458];
     assign  data_out[7505] = data_in[1723];
     assign  data_out[7506] = data_in[934];
     assign  data_out[7507] = data_in[369];
     assign  data_out[7508] = data_in[1453];
     assign  data_out[7509] = data_in[1463];
     assign  data_out[7510] = data_in[327];
     assign  data_out[7511] = data_in[887];
     assign  data_out[7512] = data_in[1193];
     assign  data_out[7513] = data_in[1026];
     assign  data_out[7514] = data_in[759];
     assign  data_out[7515] = data_in[278];
     assign  data_out[7516] = data_in[1641];
     assign  data_out[7517] = data_in[54];
     assign  data_out[7518] = data_in[25];
     assign  data_out[7519] = data_in[294];
     assign  data_out[7520] = data_in[888];
     assign  data_out[7521] = data_in[285];
     assign  data_out[7522] = data_in[558];
     assign  data_out[7523] = data_in[944];
     assign  data_out[7524] = data_in[323];
     assign  data_out[7525] = data_in[1084];
     assign  data_out[7526] = data_in[1448];
     assign  data_out[7527] = data_in[447];
     assign  data_out[7528] = data_in[668];
     assign  data_out[7529] = data_in[1184];
     assign  data_out[7530] = data_in[1205];
     assign  data_out[7531] = data_in[996];
     assign  data_out[7532] = data_in[1321];
     assign  data_out[7533] = data_in[870];
     assign  data_out[7534] = data_in[936];
     assign  data_out[7535] = data_in[1158];
     assign  data_out[7536] = data_in[47];
     assign  data_out[7537] = data_in[1406];
     assign  data_out[7538] = data_in[230];
     assign  data_out[7539] = data_in[1534];
     assign  data_out[7540] = data_in[1261];
     assign  data_out[7541] = data_in[1119];
     assign  data_out[7542] = data_in[1341];
     assign  data_out[7543] = data_in[1057];
     assign  data_out[7544] = data_in[580];
     assign  data_out[7545] = data_in[505];
     assign  data_out[7546] = data_in[141];
     assign  data_out[7547] = data_in[169];
     assign  data_out[7548] = data_in[540];
     assign  data_out[7549] = data_in[211];
     assign  data_out[7550] = data_in[159];
     assign  data_out[7551] = data_in[374];
     assign  data_out[7552] = data_in[957];
     assign  data_out[7553] = data_in[799];
     assign  data_out[7554] = data_in[548];
     assign  data_out[7555] = data_in[830];
     assign  data_out[7556] = data_in[1555];
     assign  data_out[7557] = data_in[253];
     assign  data_out[7558] = data_in[1197];
     assign  data_out[7559] = data_in[494];
     assign  data_out[7560] = data_in[86];
     assign  data_out[7561] = data_in[1576];
     assign  data_out[7562] = data_in[8];
     assign  data_out[7563] = data_in[1322];
     assign  data_out[7564] = data_in[1091];
     assign  data_out[7565] = data_in[529];
     assign  data_out[7566] = data_in[1404];
     assign  data_out[7567] = data_in[259];
     assign  data_out[7568] = data_in[1258];
     assign  data_out[7569] = data_in[420];
     assign  data_out[7570] = data_in[671];
     assign  data_out[7571] = data_in[115];
     assign  data_out[7572] = data_in[1077];
     assign  data_out[7573] = data_in[1523];
     assign  data_out[7574] = data_in[1249];
     assign  data_out[7575] = data_in[1134];
     assign  data_out[7576] = data_in[112];
     assign  data_out[7577] = data_in[1671];
     assign  data_out[7578] = data_in[190];
     assign  data_out[7579] = data_in[1611];
     assign  data_out[7580] = data_in[1408];
     assign  data_out[7581] = data_in[529];
     assign  data_out[7582] = data_in[620];
     assign  data_out[7583] = data_in[489];
     assign  data_out[7584] = data_in[1331];
     assign  data_out[7585] = data_in[904];
     assign  data_out[7586] = data_in[259];
     assign  data_out[7587] = data_in[896];
     assign  data_out[7588] = data_in[765];
     assign  data_out[7589] = data_in[1298];
     assign  data_out[7590] = data_in[994];
     assign  data_out[7591] = data_in[653];
     assign  data_out[7592] = data_in[119];
     assign  data_out[7593] = data_in[736];
     assign  data_out[7594] = data_in[679];
     assign  data_out[7595] = data_in[1543];
     assign  data_out[7596] = data_in[237];
     assign  data_out[7597] = data_in[1430];
     assign  data_out[7598] = data_in[40];
     assign  data_out[7599] = data_in[902];
     assign  data_out[7600] = data_in[1062];
     assign  data_out[7601] = data_in[918];
     assign  data_out[7602] = data_in[1419];
     assign  data_out[7603] = data_in[791];
     assign  data_out[7604] = data_in[1117];
     assign  data_out[7605] = data_in[730];
     assign  data_out[7606] = data_in[1134];
     assign  data_out[7607] = data_in[27];
     assign  data_out[7608] = data_in[40];
     assign  data_out[7609] = data_in[748];
     assign  data_out[7610] = data_in[567];
     assign  data_out[7611] = data_in[872];
     assign  data_out[7612] = data_in[314];
     assign  data_out[7613] = data_in[1131];
     assign  data_out[7614] = data_in[1480];
     assign  data_out[7615] = data_in[856];
     assign  data_out[7616] = data_in[58];
     assign  data_out[7617] = data_in[1698];
     assign  data_out[7618] = data_in[281];
     assign  data_out[7619] = data_in[1529];
     assign  data_out[7620] = data_in[678];
     assign  data_out[7621] = data_in[1650];
     assign  data_out[7622] = data_in[332];
     assign  data_out[7623] = data_in[1154];
     assign  data_out[7624] = data_in[504];
     assign  data_out[7625] = data_in[1610];
     assign  data_out[7626] = data_in[1717];
     assign  data_out[7627] = data_in[1409];
     assign  data_out[7628] = data_in[1662];
     assign  data_out[7629] = data_in[479];
     assign  data_out[7630] = data_in[1372];
     assign  data_out[7631] = data_in[306];
     assign  data_out[7632] = data_in[1316];
     assign  data_out[7633] = data_in[1216];
     assign  data_out[7634] = data_in[1039];
     assign  data_out[7635] = data_in[1385];
     assign  data_out[7636] = data_in[1437];
     assign  data_out[7637] = data_in[736];
     assign  data_out[7638] = data_in[621];
     assign  data_out[7639] = data_in[1020];
     assign  data_out[7640] = data_in[1316];
     assign  data_out[7641] = data_in[497];
     assign  data_out[7642] = data_in[337];
     assign  data_out[7643] = data_in[1188];
     assign  data_out[7644] = data_in[83];
     assign  data_out[7645] = data_in[892];
     assign  data_out[7646] = data_in[1351];
     assign  data_out[7647] = data_in[884];
     assign  data_out[7648] = data_in[1075];
     assign  data_out[7649] = data_in[446];
     assign  data_out[7650] = data_in[612];
     assign  data_out[7651] = data_in[1443];
     assign  data_out[7652] = data_in[405];
     assign  data_out[7653] = data_in[959];
     assign  data_out[7654] = data_in[700];
     assign  data_out[7655] = data_in[1420];
     assign  data_out[7656] = data_in[1680];
     assign  data_out[7657] = data_in[1585];
     assign  data_out[7658] = data_in[1025];
     assign  data_out[7659] = data_in[729];
     assign  data_out[7660] = data_in[1195];
     assign  data_out[7661] = data_in[254];
     assign  data_out[7662] = data_in[1556];
     assign  data_out[7663] = data_in[67];
     assign  data_out[7664] = data_in[1123];
     assign  data_out[7665] = data_in[984];
     assign  data_out[7666] = data_in[959];
     assign  data_out[7667] = data_in[1499];
     assign  data_out[7668] = data_in[200];
     assign  data_out[7669] = data_in[569];
     assign  data_out[7670] = data_in[1336];
     assign  data_out[7671] = data_in[1399];
     assign  data_out[7672] = data_in[410];
     assign  data_out[7673] = data_in[1572];
     assign  data_out[7674] = data_in[1428];
     assign  data_out[7675] = data_in[664];
     assign  data_out[7676] = data_in[1644];
     assign  data_out[7677] = data_in[907];
     assign  data_out[7678] = data_in[845];
     assign  data_out[7679] = data_in[899];
     assign  data_out[7680] = data_in[379];
     assign  data_out[7681] = data_in[947];
     assign  data_out[7682] = data_in[655];
     assign  data_out[7683] = data_in[1132];
     assign  data_out[7684] = data_in[621];
     assign  data_out[7685] = data_in[1085];
     assign  data_out[7686] = data_in[399];
     assign  data_out[7687] = data_in[61];
     assign  data_out[7688] = data_in[1332];
     assign  data_out[7689] = data_in[1127];
     assign  data_out[7690] = data_in[1099];
     assign  data_out[7691] = data_in[1090];
     assign  data_out[7692] = data_in[1414];
     assign  data_out[7693] = data_in[363];
     assign  data_out[7694] = data_in[473];
     assign  data_out[7695] = data_in[971];
     assign  data_out[7696] = data_in[287];
     assign  data_out[7697] = data_in[1238];
     assign  data_out[7698] = data_in[286];
     assign  data_out[7699] = data_in[792];
     assign  data_out[7700] = data_in[594];
     assign  data_out[7701] = data_in[1468];
     assign  data_out[7702] = data_in[1715];
     assign  data_out[7703] = data_in[1101];
     assign  data_out[7704] = data_in[1406];
     assign  data_out[7705] = data_in[790];
     assign  data_out[7706] = data_in[1717];
     assign  data_out[7707] = data_in[916];
     assign  data_out[7708] = data_in[585];
     assign  data_out[7709] = data_in[1024];
     assign  data_out[7710] = data_in[844];
     assign  data_out[7711] = data_in[418];
     assign  data_out[7712] = data_in[1582];
     assign  data_out[7713] = data_in[1439];
     assign  data_out[7714] = data_in[946];
     assign  data_out[7715] = data_in[1145];
     assign  data_out[7716] = data_in[112];
     assign  data_out[7717] = data_in[921];
     assign  data_out[7718] = data_in[1459];
     assign  data_out[7719] = data_in[65];
     assign  data_out[7720] = data_in[1304];
     assign  data_out[7721] = data_in[321];
     assign  data_out[7722] = data_in[384];
     assign  data_out[7723] = data_in[678];
     assign  data_out[7724] = data_in[1280];
     assign  data_out[7725] = data_in[897];
     assign  data_out[7726] = data_in[4];
     assign  data_out[7727] = data_in[1265];
     assign  data_out[7728] = data_in[1043];
     assign  data_out[7729] = data_in[891];
     assign  data_out[7730] = data_in[987];
     assign  data_out[7731] = data_in[703];
     assign  data_out[7732] = data_in[457];
     assign  data_out[7733] = data_in[1705];
     assign  data_out[7734] = data_in[466];
     assign  data_out[7735] = data_in[978];
     assign  data_out[7736] = data_in[450];
     assign  data_out[7737] = data_in[1507];
     assign  data_out[7738] = data_in[215];
     assign  data_out[7739] = data_in[158];
     assign  data_out[7740] = data_in[969];
     assign  data_out[7741] = data_in[1581];
     assign  data_out[7742] = data_in[770];
     assign  data_out[7743] = data_in[1601];
     assign  data_out[7744] = data_in[357];
     assign  data_out[7745] = data_in[1507];
     assign  data_out[7746] = data_in[1428];
     assign  data_out[7747] = data_in[357];
     assign  data_out[7748] = data_in[956];
     assign  data_out[7749] = data_in[1573];
     assign  data_out[7750] = data_in[994];
     assign  data_out[7751] = data_in[149];
     assign  data_out[7752] = data_in[685];
     assign  data_out[7753] = data_in[604];
     assign  data_out[7754] = data_in[184];
     assign  data_out[7755] = data_in[1191];
     assign  data_out[7756] = data_in[1321];
     assign  data_out[7757] = data_in[710];
     assign  data_out[7758] = data_in[572];
     assign  data_out[7759] = data_in[113];
     assign  data_out[7760] = data_in[1144];
     assign  data_out[7761] = data_in[206];
     assign  data_out[7762] = data_in[981];
     assign  data_out[7763] = data_in[999];
     assign  data_out[7764] = data_in[926];
     assign  data_out[7765] = data_in[37];
     assign  data_out[7766] = data_in[24];
     assign  data_out[7767] = data_in[1072];
     assign  data_out[7768] = data_in[1303];
     assign  data_out[7769] = data_in[1513];
     assign  data_out[7770] = data_in[524];
     assign  data_out[7771] = data_in[111];
     assign  data_out[7772] = data_in[1514];
     assign  data_out[7773] = data_in[1672];
     assign  data_out[7774] = data_in[316];
     assign  data_out[7775] = data_in[618];

endmodule