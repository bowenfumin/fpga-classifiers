
module lut_4level_tree3(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [7775:0] data_in,
                       input       data_valid,
                       output  reg data_out     
                       );

wire    [7775:0] to_level4;
(*S="TRUE"*)reg     [7775:0] level4_in;
wire    [1295:0] to_level3;
(*S="TRUE"*)reg     [1295:0] level3_in;
wire    [215:0] to_level2;
(*S="TRUE"*)reg     [215:0] level2_in;
wire    [35:0] to_level1;
(*S="TRUE"*)reg     [35:0] level1_in;
wire    [5:0] to_level0;
(*S="TRUE"*)reg     [5:0] level0_in;
wire          data_out_temp;


assign  to_level4 = data_in;

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level4_in <= 7776'b0;
  else
    level4_in <= to_level4;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level3_in <= 1296'b0;
  else
    level3_in <= to_level3;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level2_in <= 216'b0;
  else
    level2_in <= to_level2;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level1_in <= 36'b0;
  else
    level1_in <= to_level1;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level0_in <= 6'b0;
  else
    level0_in <= to_level0;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    data_out <= 1'b0;
  else
    if(data_valid == 1'b1)
      data_out <= data_out_temp;
    else;
end
////////////// level 4 starts below:/n
LUT6 #(
   .INIT(64'h8254551282545512)  
) LUT6_inst7776 (
   .O(to_level3[0]),
   .I0(level4_in[0]),
   .I1(level4_in[1]),
   .I2(level4_in[2]),
   .I3(level4_in[3]),
   .I4(level4_in[4]),
   .I5(level4_in[5])
);

LUT6 #(
   .INIT(64'he4f4250be4f4250b)  
) LUT6_inst7777 (
   .O(to_level3[1]),
   .I0(level4_in[6]),
   .I1(level4_in[7]),
   .I2(level4_in[8]),
   .I3(level4_in[9]),
   .I4(level4_in[10]),
   .I5(level4_in[11])
);

LUT6 #(
   .INIT(64'h833f52e3833f52e3)  
) LUT6_inst7778 (
   .O(to_level3[2]),
   .I0(level4_in[12]),
   .I1(level4_in[13]),
   .I2(level4_in[14]),
   .I3(level4_in[15]),
   .I4(level4_in[16]),
   .I5(level4_in[17])
);

LUT6 #(
   .INIT(64'h8e6091e78e6091e7)  
) LUT6_inst7779 (
   .O(to_level3[3]),
   .I0(level4_in[18]),
   .I1(level4_in[19]),
   .I2(level4_in[20]),
   .I3(level4_in[21]),
   .I4(level4_in[22]),
   .I5(level4_in[23])
);

LUT6 #(
   .INIT(64'ha01b2e8ca01b2e8c)  
) LUT6_inst7780 (
   .O(to_level3[4]),
   .I0(level4_in[24]),
   .I1(level4_in[25]),
   .I2(level4_in[26]),
   .I3(level4_in[27]),
   .I4(level4_in[28]),
   .I5(level4_in[29])
);

LUT6 #(
   .INIT(64'h7a4d7fff7a4d7fff)  
) LUT6_inst7781 (
   .O(to_level3[5]),
   .I0(level4_in[30]),
   .I1(level4_in[31]),
   .I2(level4_in[32]),
   .I3(level4_in[33]),
   .I4(level4_in[34]),
   .I5(level4_in[35])
);

LUT6 #(
   .INIT(64'h0ace32280ace3228)  
) LUT6_inst7782 (
   .O(to_level3[6]),
   .I0(level4_in[36]),
   .I1(level4_in[37]),
   .I2(level4_in[38]),
   .I3(level4_in[39]),
   .I4(level4_in[40]),
   .I5(level4_in[41])
);

LUT6 #(
   .INIT(64'hb0e64c1eb0e64c1e)  
) LUT6_inst7783 (
   .O(to_level3[7]),
   .I0(level4_in[42]),
   .I1(level4_in[43]),
   .I2(level4_in[44]),
   .I3(level4_in[45]),
   .I4(level4_in[46]),
   .I5(level4_in[47])
);

LUT6 #(
   .INIT(64'hfec1c46efec1c46e)  
) LUT6_inst7784 (
   .O(to_level3[8]),
   .I0(level4_in[48]),
   .I1(level4_in[49]),
   .I2(level4_in[50]),
   .I3(level4_in[51]),
   .I4(level4_in[52]),
   .I5(level4_in[53])
);

LUT6 #(
   .INIT(64'h3157b4a63157b4a6)  
) LUT6_inst7785 (
   .O(to_level3[9]),
   .I0(level4_in[54]),
   .I1(level4_in[55]),
   .I2(level4_in[56]),
   .I3(level4_in[57]),
   .I4(level4_in[58]),
   .I5(level4_in[59])
);

LUT6 #(
   .INIT(64'h1626e46c1626e46c)  
) LUT6_inst7786 (
   .O(to_level3[10]),
   .I0(level4_in[60]),
   .I1(level4_in[61]),
   .I2(level4_in[62]),
   .I3(level4_in[63]),
   .I4(level4_in[64]),
   .I5(level4_in[65])
);

LUT6 #(
   .INIT(64'h8561f29e8561f29e)  
) LUT6_inst7787 (
   .O(to_level3[11]),
   .I0(level4_in[66]),
   .I1(level4_in[67]),
   .I2(level4_in[68]),
   .I3(level4_in[69]),
   .I4(level4_in[70]),
   .I5(level4_in[71])
);

LUT6 #(
   .INIT(64'h5a1791fe5a1791fe)  
) LUT6_inst7788 (
   .O(to_level3[12]),
   .I0(level4_in[72]),
   .I1(level4_in[73]),
   .I2(level4_in[74]),
   .I3(level4_in[75]),
   .I4(level4_in[76]),
   .I5(level4_in[77])
);

LUT6 #(
   .INIT(64'h550a96a8550a96a8)  
) LUT6_inst7789 (
   .O(to_level3[13]),
   .I0(level4_in[78]),
   .I1(level4_in[79]),
   .I2(level4_in[80]),
   .I3(level4_in[81]),
   .I4(level4_in[82]),
   .I5(level4_in[83])
);

LUT6 #(
   .INIT(64'h579cd8bd579cd8bd)  
) LUT6_inst7790 (
   .O(to_level3[14]),
   .I0(level4_in[84]),
   .I1(level4_in[85]),
   .I2(level4_in[86]),
   .I3(level4_in[87]),
   .I4(level4_in[88]),
   .I5(level4_in[89])
);

LUT6 #(
   .INIT(64'h74f5034f74f5034f)  
) LUT6_inst7791 (
   .O(to_level3[15]),
   .I0(level4_in[90]),
   .I1(level4_in[91]),
   .I2(level4_in[92]),
   .I3(level4_in[93]),
   .I4(level4_in[94]),
   .I5(level4_in[95])
);

LUT6 #(
   .INIT(64'h57f7fb2357f7fb23)  
) LUT6_inst7792 (
   .O(to_level3[16]),
   .I0(level4_in[96]),
   .I1(level4_in[97]),
   .I2(level4_in[98]),
   .I3(level4_in[99]),
   .I4(level4_in[100]),
   .I5(level4_in[101])
);

LUT6 #(
   .INIT(64'he869352ee869352e)  
) LUT6_inst7793 (
   .O(to_level3[17]),
   .I0(level4_in[102]),
   .I1(level4_in[103]),
   .I2(level4_in[104]),
   .I3(level4_in[105]),
   .I4(level4_in[106]),
   .I5(level4_in[107])
);

LUT6 #(
   .INIT(64'h709dbdea709dbdea)  
) LUT6_inst7794 (
   .O(to_level3[18]),
   .I0(level4_in[108]),
   .I1(level4_in[109]),
   .I2(level4_in[110]),
   .I3(level4_in[111]),
   .I4(level4_in[112]),
   .I5(level4_in[113])
);

LUT6 #(
   .INIT(64'h07bf3fca07bf3fca)  
) LUT6_inst7795 (
   .O(to_level3[19]),
   .I0(level4_in[114]),
   .I1(level4_in[115]),
   .I2(level4_in[116]),
   .I3(level4_in[117]),
   .I4(level4_in[118]),
   .I5(level4_in[119])
);

LUT6 #(
   .INIT(64'hba6127a3ba6127a3)  
) LUT6_inst7796 (
   .O(to_level3[20]),
   .I0(level4_in[120]),
   .I1(level4_in[121]),
   .I2(level4_in[122]),
   .I3(level4_in[123]),
   .I4(level4_in[124]),
   .I5(level4_in[125])
);

LUT6 #(
   .INIT(64'hdfcbff00dfcbff00)  
) LUT6_inst7797 (
   .O(to_level3[21]),
   .I0(level4_in[126]),
   .I1(level4_in[127]),
   .I2(level4_in[128]),
   .I3(level4_in[129]),
   .I4(level4_in[130]),
   .I5(level4_in[131])
);

LUT6 #(
   .INIT(64'h1bcdeb621bcdeb62)  
) LUT6_inst7798 (
   .O(to_level3[22]),
   .I0(level4_in[132]),
   .I1(level4_in[133]),
   .I2(level4_in[134]),
   .I3(level4_in[135]),
   .I4(level4_in[136]),
   .I5(level4_in[137])
);

LUT6 #(
   .INIT(64'hcfe4b039cfe4b039)  
) LUT6_inst7799 (
   .O(to_level3[23]),
   .I0(level4_in[138]),
   .I1(level4_in[139]),
   .I2(level4_in[140]),
   .I3(level4_in[141]),
   .I4(level4_in[142]),
   .I5(level4_in[143])
);

LUT6 #(
   .INIT(64'hefbe65a6efbe65a6)  
) LUT6_inst7800 (
   .O(to_level3[24]),
   .I0(level4_in[144]),
   .I1(level4_in[145]),
   .I2(level4_in[146]),
   .I3(level4_in[147]),
   .I4(level4_in[148]),
   .I5(level4_in[149])
);

LUT6 #(
   .INIT(64'h1362ecf81362ecf8)  
) LUT6_inst7801 (
   .O(to_level3[25]),
   .I0(level4_in[150]),
   .I1(level4_in[151]),
   .I2(level4_in[152]),
   .I3(level4_in[153]),
   .I4(level4_in[154]),
   .I5(level4_in[155])
);

LUT6 #(
   .INIT(64'ha5fbd945a5fbd945)  
) LUT6_inst7802 (
   .O(to_level3[26]),
   .I0(level4_in[156]),
   .I1(level4_in[157]),
   .I2(level4_in[158]),
   .I3(level4_in[159]),
   .I4(level4_in[160]),
   .I5(level4_in[161])
);

LUT6 #(
   .INIT(64'hef143d84ef143d84)  
) LUT6_inst7803 (
   .O(to_level3[27]),
   .I0(level4_in[162]),
   .I1(level4_in[163]),
   .I2(level4_in[164]),
   .I3(level4_in[165]),
   .I4(level4_in[166]),
   .I5(level4_in[167])
);

LUT6 #(
   .INIT(64'h55328f1355328f13)  
) LUT6_inst7804 (
   .O(to_level3[28]),
   .I0(level4_in[168]),
   .I1(level4_in[169]),
   .I2(level4_in[170]),
   .I3(level4_in[171]),
   .I4(level4_in[172]),
   .I5(level4_in[173])
);

LUT6 #(
   .INIT(64'h54da210054da2100)  
) LUT6_inst7805 (
   .O(to_level3[29]),
   .I0(level4_in[174]),
   .I1(level4_in[175]),
   .I2(level4_in[176]),
   .I3(level4_in[177]),
   .I4(level4_in[178]),
   .I5(level4_in[179])
);

LUT6 #(
   .INIT(64'h9e1eba529e1eba52)  
) LUT6_inst7806 (
   .O(to_level3[30]),
   .I0(level4_in[180]),
   .I1(level4_in[181]),
   .I2(level4_in[182]),
   .I3(level4_in[183]),
   .I4(level4_in[184]),
   .I5(level4_in[185])
);

LUT6 #(
   .INIT(64'hb0b4aa47b0b4aa47)  
) LUT6_inst7807 (
   .O(to_level3[31]),
   .I0(level4_in[186]),
   .I1(level4_in[187]),
   .I2(level4_in[188]),
   .I3(level4_in[189]),
   .I4(level4_in[190]),
   .I5(level4_in[191])
);

LUT6 #(
   .INIT(64'h7f67e1837f67e183)  
) LUT6_inst7808 (
   .O(to_level3[32]),
   .I0(level4_in[192]),
   .I1(level4_in[193]),
   .I2(level4_in[194]),
   .I3(level4_in[195]),
   .I4(level4_in[196]),
   .I5(level4_in[197])
);

LUT6 #(
   .INIT(64'h64d5812364d58123)  
) LUT6_inst7809 (
   .O(to_level3[33]),
   .I0(level4_in[198]),
   .I1(level4_in[199]),
   .I2(level4_in[200]),
   .I3(level4_in[201]),
   .I4(level4_in[202]),
   .I5(level4_in[203])
);

LUT6 #(
   .INIT(64'h1e35ecfa1e35ecfa)  
) LUT6_inst7810 (
   .O(to_level3[34]),
   .I0(level4_in[204]),
   .I1(level4_in[205]),
   .I2(level4_in[206]),
   .I3(level4_in[207]),
   .I4(level4_in[208]),
   .I5(level4_in[209])
);

LUT6 #(
   .INIT(64'h40b378ac40b378ac)  
) LUT6_inst7811 (
   .O(to_level3[35]),
   .I0(level4_in[210]),
   .I1(level4_in[211]),
   .I2(level4_in[212]),
   .I3(level4_in[213]),
   .I4(level4_in[214]),
   .I5(level4_in[215])
);

LUT6 #(
   .INIT(64'h66001e4f66001e4f)  
) LUT6_inst7812 (
   .O(to_level3[36]),
   .I0(level4_in[216]),
   .I1(level4_in[217]),
   .I2(level4_in[218]),
   .I3(level4_in[219]),
   .I4(level4_in[220]),
   .I5(level4_in[221])
);

LUT6 #(
   .INIT(64'hcb3e2bebcb3e2beb)  
) LUT6_inst7813 (
   .O(to_level3[37]),
   .I0(level4_in[222]),
   .I1(level4_in[223]),
   .I2(level4_in[224]),
   .I3(level4_in[225]),
   .I4(level4_in[226]),
   .I5(level4_in[227])
);

LUT6 #(
   .INIT(64'h6fa74c3e6fa74c3e)  
) LUT6_inst7814 (
   .O(to_level3[38]),
   .I0(level4_in[228]),
   .I1(level4_in[229]),
   .I2(level4_in[230]),
   .I3(level4_in[231]),
   .I4(level4_in[232]),
   .I5(level4_in[233])
);

LUT6 #(
   .INIT(64'hc0ea637dc0ea637d)  
) LUT6_inst7815 (
   .O(to_level3[39]),
   .I0(level4_in[234]),
   .I1(level4_in[235]),
   .I2(level4_in[236]),
   .I3(level4_in[237]),
   .I4(level4_in[238]),
   .I5(level4_in[239])
);

LUT6 #(
   .INIT(64'h58d9192f58d9192f)  
) LUT6_inst7816 (
   .O(to_level3[40]),
   .I0(level4_in[240]),
   .I1(level4_in[241]),
   .I2(level4_in[242]),
   .I3(level4_in[243]),
   .I4(level4_in[244]),
   .I5(level4_in[245])
);

LUT6 #(
   .INIT(64'hf50a7954f50a7954)  
) LUT6_inst7817 (
   .O(to_level3[41]),
   .I0(level4_in[246]),
   .I1(level4_in[247]),
   .I2(level4_in[248]),
   .I3(level4_in[249]),
   .I4(level4_in[250]),
   .I5(level4_in[251])
);

LUT6 #(
   .INIT(64'hb0d4f1d0b0d4f1d0)  
) LUT6_inst7818 (
   .O(to_level3[42]),
   .I0(level4_in[252]),
   .I1(level4_in[253]),
   .I2(level4_in[254]),
   .I3(level4_in[255]),
   .I4(level4_in[256]),
   .I5(level4_in[257])
);

LUT6 #(
   .INIT(64'h0779c4380779c438)  
) LUT6_inst7819 (
   .O(to_level3[43]),
   .I0(level4_in[258]),
   .I1(level4_in[259]),
   .I2(level4_in[260]),
   .I3(level4_in[261]),
   .I4(level4_in[262]),
   .I5(level4_in[263])
);

LUT6 #(
   .INIT(64'h54e761bf54e761bf)  
) LUT6_inst7820 (
   .O(to_level3[44]),
   .I0(level4_in[264]),
   .I1(level4_in[265]),
   .I2(level4_in[266]),
   .I3(level4_in[267]),
   .I4(level4_in[268]),
   .I5(level4_in[269])
);

LUT6 #(
   .INIT(64'h6345726a6345726a)  
) LUT6_inst7821 (
   .O(to_level3[45]),
   .I0(level4_in[270]),
   .I1(level4_in[271]),
   .I2(level4_in[272]),
   .I3(level4_in[273]),
   .I4(level4_in[274]),
   .I5(level4_in[275])
);

LUT6 #(
   .INIT(64'he544c112e544c112)  
) LUT6_inst7822 (
   .O(to_level3[46]),
   .I0(level4_in[276]),
   .I1(level4_in[277]),
   .I2(level4_in[278]),
   .I3(level4_in[279]),
   .I4(level4_in[280]),
   .I5(level4_in[281])
);

LUT6 #(
   .INIT(64'hef883217ef883217)  
) LUT6_inst7823 (
   .O(to_level3[47]),
   .I0(level4_in[282]),
   .I1(level4_in[283]),
   .I2(level4_in[284]),
   .I3(level4_in[285]),
   .I4(level4_in[286]),
   .I5(level4_in[287])
);

LUT6 #(
   .INIT(64'h6256d0276256d027)  
) LUT6_inst7824 (
   .O(to_level3[48]),
   .I0(level4_in[288]),
   .I1(level4_in[289]),
   .I2(level4_in[290]),
   .I3(level4_in[291]),
   .I4(level4_in[292]),
   .I5(level4_in[293])
);

LUT6 #(
   .INIT(64'h78637c8978637c89)  
) LUT6_inst7825 (
   .O(to_level3[49]),
   .I0(level4_in[294]),
   .I1(level4_in[295]),
   .I2(level4_in[296]),
   .I3(level4_in[297]),
   .I4(level4_in[298]),
   .I5(level4_in[299])
);

LUT6 #(
   .INIT(64'he5c9ac17e5c9ac17)  
) LUT6_inst7826 (
   .O(to_level3[50]),
   .I0(level4_in[300]),
   .I1(level4_in[301]),
   .I2(level4_in[302]),
   .I3(level4_in[303]),
   .I4(level4_in[304]),
   .I5(level4_in[305])
);

LUT6 #(
   .INIT(64'h4887afe84887afe8)  
) LUT6_inst7827 (
   .O(to_level3[51]),
   .I0(level4_in[306]),
   .I1(level4_in[307]),
   .I2(level4_in[308]),
   .I3(level4_in[309]),
   .I4(level4_in[310]),
   .I5(level4_in[311])
);

LUT6 #(
   .INIT(64'h5b8bbd535b8bbd53)  
) LUT6_inst7828 (
   .O(to_level3[52]),
   .I0(level4_in[312]),
   .I1(level4_in[313]),
   .I2(level4_in[314]),
   .I3(level4_in[315]),
   .I4(level4_in[316]),
   .I5(level4_in[317])
);

LUT6 #(
   .INIT(64'h4fe226df4fe226df)  
) LUT6_inst7829 (
   .O(to_level3[53]),
   .I0(level4_in[318]),
   .I1(level4_in[319]),
   .I2(level4_in[320]),
   .I3(level4_in[321]),
   .I4(level4_in[322]),
   .I5(level4_in[323])
);

LUT6 #(
   .INIT(64'h9e1d10919e1d1091)  
) LUT6_inst7830 (
   .O(to_level3[54]),
   .I0(level4_in[324]),
   .I1(level4_in[325]),
   .I2(level4_in[326]),
   .I3(level4_in[327]),
   .I4(level4_in[328]),
   .I5(level4_in[329])
);

LUT6 #(
   .INIT(64'hc4029928c4029928)  
) LUT6_inst7831 (
   .O(to_level3[55]),
   .I0(level4_in[330]),
   .I1(level4_in[331]),
   .I2(level4_in[332]),
   .I3(level4_in[333]),
   .I4(level4_in[334]),
   .I5(level4_in[335])
);

LUT6 #(
   .INIT(64'hefc4addfefc4addf)  
) LUT6_inst7832 (
   .O(to_level3[56]),
   .I0(level4_in[336]),
   .I1(level4_in[337]),
   .I2(level4_in[338]),
   .I3(level4_in[339]),
   .I4(level4_in[340]),
   .I5(level4_in[341])
);

LUT6 #(
   .INIT(64'hf748ce38f748ce38)  
) LUT6_inst7833 (
   .O(to_level3[57]),
   .I0(level4_in[342]),
   .I1(level4_in[343]),
   .I2(level4_in[344]),
   .I3(level4_in[345]),
   .I4(level4_in[346]),
   .I5(level4_in[347])
);

LUT6 #(
   .INIT(64'hb06007c4b06007c4)  
) LUT6_inst7834 (
   .O(to_level3[58]),
   .I0(level4_in[348]),
   .I1(level4_in[349]),
   .I2(level4_in[350]),
   .I3(level4_in[351]),
   .I4(level4_in[352]),
   .I5(level4_in[353])
);

LUT6 #(
   .INIT(64'hedbaebf5edbaebf5)  
) LUT6_inst7835 (
   .O(to_level3[59]),
   .I0(level4_in[354]),
   .I1(level4_in[355]),
   .I2(level4_in[356]),
   .I3(level4_in[357]),
   .I4(level4_in[358]),
   .I5(level4_in[359])
);

LUT6 #(
   .INIT(64'hd0d8c0b6d0d8c0b6)  
) LUT6_inst7836 (
   .O(to_level3[60]),
   .I0(level4_in[360]),
   .I1(level4_in[361]),
   .I2(level4_in[362]),
   .I3(level4_in[363]),
   .I4(level4_in[364]),
   .I5(level4_in[365])
);

LUT6 #(
   .INIT(64'h9063cd129063cd12)  
) LUT6_inst7837 (
   .O(to_level3[61]),
   .I0(level4_in[366]),
   .I1(level4_in[367]),
   .I2(level4_in[368]),
   .I3(level4_in[369]),
   .I4(level4_in[370]),
   .I5(level4_in[371])
);

LUT6 #(
   .INIT(64'hc2dfa8c4c2dfa8c4)  
) LUT6_inst7838 (
   .O(to_level3[62]),
   .I0(level4_in[372]),
   .I1(level4_in[373]),
   .I2(level4_in[374]),
   .I3(level4_in[375]),
   .I4(level4_in[376]),
   .I5(level4_in[377])
);

LUT6 #(
   .INIT(64'h307adf1c307adf1c)  
) LUT6_inst7839 (
   .O(to_level3[63]),
   .I0(level4_in[378]),
   .I1(level4_in[379]),
   .I2(level4_in[380]),
   .I3(level4_in[381]),
   .I4(level4_in[382]),
   .I5(level4_in[383])
);

LUT6 #(
   .INIT(64'hb77483e4b77483e4)  
) LUT6_inst7840 (
   .O(to_level3[64]),
   .I0(level4_in[384]),
   .I1(level4_in[385]),
   .I2(level4_in[386]),
   .I3(level4_in[387]),
   .I4(level4_in[388]),
   .I5(level4_in[389])
);

LUT6 #(
   .INIT(64'h133b398d133b398d)  
) LUT6_inst7841 (
   .O(to_level3[65]),
   .I0(level4_in[390]),
   .I1(level4_in[391]),
   .I2(level4_in[392]),
   .I3(level4_in[393]),
   .I4(level4_in[394]),
   .I5(level4_in[395])
);

LUT6 #(
   .INIT(64'h7ccbb7277ccbb727)  
) LUT6_inst7842 (
   .O(to_level3[66]),
   .I0(level4_in[396]),
   .I1(level4_in[397]),
   .I2(level4_in[398]),
   .I3(level4_in[399]),
   .I4(level4_in[400]),
   .I5(level4_in[401])
);

LUT6 #(
   .INIT(64'h0d5407fd0d5407fd)  
) LUT6_inst7843 (
   .O(to_level3[67]),
   .I0(level4_in[402]),
   .I1(level4_in[403]),
   .I2(level4_in[404]),
   .I3(level4_in[405]),
   .I4(level4_in[406]),
   .I5(level4_in[407])
);

LUT6 #(
   .INIT(64'hf082d0c7f082d0c7)  
) LUT6_inst7844 (
   .O(to_level3[68]),
   .I0(level4_in[408]),
   .I1(level4_in[409]),
   .I2(level4_in[410]),
   .I3(level4_in[411]),
   .I4(level4_in[412]),
   .I5(level4_in[413])
);

LUT6 #(
   .INIT(64'h5ade64575ade6457)  
) LUT6_inst7845 (
   .O(to_level3[69]),
   .I0(level4_in[414]),
   .I1(level4_in[415]),
   .I2(level4_in[416]),
   .I3(level4_in[417]),
   .I4(level4_in[418]),
   .I5(level4_in[419])
);

LUT6 #(
   .INIT(64'h2fc032402fc03240)  
) LUT6_inst7846 (
   .O(to_level3[70]),
   .I0(level4_in[420]),
   .I1(level4_in[421]),
   .I2(level4_in[422]),
   .I3(level4_in[423]),
   .I4(level4_in[424]),
   .I5(level4_in[425])
);

LUT6 #(
   .INIT(64'hca6585c6ca6585c6)  
) LUT6_inst7847 (
   .O(to_level3[71]),
   .I0(level4_in[426]),
   .I1(level4_in[427]),
   .I2(level4_in[428]),
   .I3(level4_in[429]),
   .I4(level4_in[430]),
   .I5(level4_in[431])
);

LUT6 #(
   .INIT(64'h0c3ffc9b0c3ffc9b)  
) LUT6_inst7848 (
   .O(to_level3[72]),
   .I0(level4_in[432]),
   .I1(level4_in[433]),
   .I2(level4_in[434]),
   .I3(level4_in[435]),
   .I4(level4_in[436]),
   .I5(level4_in[437])
);

LUT6 #(
   .INIT(64'h06641eff06641eff)  
) LUT6_inst7849 (
   .O(to_level3[73]),
   .I0(level4_in[438]),
   .I1(level4_in[439]),
   .I2(level4_in[440]),
   .I3(level4_in[441]),
   .I4(level4_in[442]),
   .I5(level4_in[443])
);

LUT6 #(
   .INIT(64'h2c53c6152c53c615)  
) LUT6_inst7850 (
   .O(to_level3[74]),
   .I0(level4_in[444]),
   .I1(level4_in[445]),
   .I2(level4_in[446]),
   .I3(level4_in[447]),
   .I4(level4_in[448]),
   .I5(level4_in[449])
);

LUT6 #(
   .INIT(64'h8100e5388100e538)  
) LUT6_inst7851 (
   .O(to_level3[75]),
   .I0(level4_in[450]),
   .I1(level4_in[451]),
   .I2(level4_in[452]),
   .I3(level4_in[453]),
   .I4(level4_in[454]),
   .I5(level4_in[455])
);

LUT6 #(
   .INIT(64'h40a5990e40a5990e)  
) LUT6_inst7852 (
   .O(to_level3[76]),
   .I0(level4_in[456]),
   .I1(level4_in[457]),
   .I2(level4_in[458]),
   .I3(level4_in[459]),
   .I4(level4_in[460]),
   .I5(level4_in[461])
);

LUT6 #(
   .INIT(64'hdc7f7376dc7f7376)  
) LUT6_inst7853 (
   .O(to_level3[77]),
   .I0(level4_in[462]),
   .I1(level4_in[463]),
   .I2(level4_in[464]),
   .I3(level4_in[465]),
   .I4(level4_in[466]),
   .I5(level4_in[467])
);

LUT6 #(
   .INIT(64'hcc7f3b4dcc7f3b4d)  
) LUT6_inst7854 (
   .O(to_level3[78]),
   .I0(level4_in[468]),
   .I1(level4_in[469]),
   .I2(level4_in[470]),
   .I3(level4_in[471]),
   .I4(level4_in[472]),
   .I5(level4_in[473])
);

LUT6 #(
   .INIT(64'h72c3e3a372c3e3a3)  
) LUT6_inst7855 (
   .O(to_level3[79]),
   .I0(level4_in[474]),
   .I1(level4_in[475]),
   .I2(level4_in[476]),
   .I3(level4_in[477]),
   .I4(level4_in[478]),
   .I5(level4_in[479])
);

LUT6 #(
   .INIT(64'hd554d79fd554d79f)  
) LUT6_inst7856 (
   .O(to_level3[80]),
   .I0(level4_in[480]),
   .I1(level4_in[481]),
   .I2(level4_in[482]),
   .I3(level4_in[483]),
   .I4(level4_in[484]),
   .I5(level4_in[485])
);

LUT6 #(
   .INIT(64'h53761a9c53761a9c)  
) LUT6_inst7857 (
   .O(to_level3[81]),
   .I0(level4_in[486]),
   .I1(level4_in[487]),
   .I2(level4_in[488]),
   .I3(level4_in[489]),
   .I4(level4_in[490]),
   .I5(level4_in[491])
);

LUT6 #(
   .INIT(64'h3a0bd80f3a0bd80f)  
) LUT6_inst7858 (
   .O(to_level3[82]),
   .I0(level4_in[492]),
   .I1(level4_in[493]),
   .I2(level4_in[494]),
   .I3(level4_in[495]),
   .I4(level4_in[496]),
   .I5(level4_in[497])
);

LUT6 #(
   .INIT(64'h9f32d3379f32d337)  
) LUT6_inst7859 (
   .O(to_level3[83]),
   .I0(level4_in[498]),
   .I1(level4_in[499]),
   .I2(level4_in[500]),
   .I3(level4_in[501]),
   .I4(level4_in[502]),
   .I5(level4_in[503])
);

LUT6 #(
   .INIT(64'hdcc6327ddcc6327d)  
) LUT6_inst7860 (
   .O(to_level3[84]),
   .I0(level4_in[504]),
   .I1(level4_in[505]),
   .I2(level4_in[506]),
   .I3(level4_in[507]),
   .I4(level4_in[508]),
   .I5(level4_in[509])
);

LUT6 #(
   .INIT(64'hfb2b08c1fb2b08c1)  
) LUT6_inst7861 (
   .O(to_level3[85]),
   .I0(level4_in[510]),
   .I1(level4_in[511]),
   .I2(level4_in[512]),
   .I3(level4_in[513]),
   .I4(level4_in[514]),
   .I5(level4_in[515])
);

LUT6 #(
   .INIT(64'h88326d4088326d40)  
) LUT6_inst7862 (
   .O(to_level3[86]),
   .I0(level4_in[516]),
   .I1(level4_in[517]),
   .I2(level4_in[518]),
   .I3(level4_in[519]),
   .I4(level4_in[520]),
   .I5(level4_in[521])
);

LUT6 #(
   .INIT(64'hd02b8aa6d02b8aa6)  
) LUT6_inst7863 (
   .O(to_level3[87]),
   .I0(level4_in[522]),
   .I1(level4_in[523]),
   .I2(level4_in[524]),
   .I3(level4_in[525]),
   .I4(level4_in[526]),
   .I5(level4_in[527])
);

LUT6 #(
   .INIT(64'h55aca04755aca047)  
) LUT6_inst7864 (
   .O(to_level3[88]),
   .I0(level4_in[528]),
   .I1(level4_in[529]),
   .I2(level4_in[530]),
   .I3(level4_in[531]),
   .I4(level4_in[532]),
   .I5(level4_in[533])
);

LUT6 #(
   .INIT(64'h24799ef824799ef8)  
) LUT6_inst7865 (
   .O(to_level3[89]),
   .I0(level4_in[534]),
   .I1(level4_in[535]),
   .I2(level4_in[536]),
   .I3(level4_in[537]),
   .I4(level4_in[538]),
   .I5(level4_in[539])
);

LUT6 #(
   .INIT(64'haa4cf9b9aa4cf9b9)  
) LUT6_inst7866 (
   .O(to_level3[90]),
   .I0(level4_in[540]),
   .I1(level4_in[541]),
   .I2(level4_in[542]),
   .I3(level4_in[543]),
   .I4(level4_in[544]),
   .I5(level4_in[545])
);

LUT6 #(
   .INIT(64'hf185e551f185e551)  
) LUT6_inst7867 (
   .O(to_level3[91]),
   .I0(level4_in[546]),
   .I1(level4_in[547]),
   .I2(level4_in[548]),
   .I3(level4_in[549]),
   .I4(level4_in[550]),
   .I5(level4_in[551])
);

LUT6 #(
   .INIT(64'h3af1778d3af1778d)  
) LUT6_inst7868 (
   .O(to_level3[92]),
   .I0(level4_in[552]),
   .I1(level4_in[553]),
   .I2(level4_in[554]),
   .I3(level4_in[555]),
   .I4(level4_in[556]),
   .I5(level4_in[557])
);

LUT6 #(
   .INIT(64'h2571a9f32571a9f3)  
) LUT6_inst7869 (
   .O(to_level3[93]),
   .I0(level4_in[558]),
   .I1(level4_in[559]),
   .I2(level4_in[560]),
   .I3(level4_in[561]),
   .I4(level4_in[562]),
   .I5(level4_in[563])
);

LUT6 #(
   .INIT(64'h7bb726727bb72672)  
) LUT6_inst7870 (
   .O(to_level3[94]),
   .I0(level4_in[564]),
   .I1(level4_in[565]),
   .I2(level4_in[566]),
   .I3(level4_in[567]),
   .I4(level4_in[568]),
   .I5(level4_in[569])
);

LUT6 #(
   .INIT(64'hc48d923ac48d923a)  
) LUT6_inst7871 (
   .O(to_level3[95]),
   .I0(level4_in[570]),
   .I1(level4_in[571]),
   .I2(level4_in[572]),
   .I3(level4_in[573]),
   .I4(level4_in[574]),
   .I5(level4_in[575])
);

LUT6 #(
   .INIT(64'h5497673e5497673e)  
) LUT6_inst7872 (
   .O(to_level3[96]),
   .I0(level4_in[576]),
   .I1(level4_in[577]),
   .I2(level4_in[578]),
   .I3(level4_in[579]),
   .I4(level4_in[580]),
   .I5(level4_in[581])
);

LUT6 #(
   .INIT(64'h293e5423293e5423)  
) LUT6_inst7873 (
   .O(to_level3[97]),
   .I0(level4_in[582]),
   .I1(level4_in[583]),
   .I2(level4_in[584]),
   .I3(level4_in[585]),
   .I4(level4_in[586]),
   .I5(level4_in[587])
);

LUT6 #(
   .INIT(64'hc70adb84c70adb84)  
) LUT6_inst7874 (
   .O(to_level3[98]),
   .I0(level4_in[588]),
   .I1(level4_in[589]),
   .I2(level4_in[590]),
   .I3(level4_in[591]),
   .I4(level4_in[592]),
   .I5(level4_in[593])
);

LUT6 #(
   .INIT(64'hfd5b6814fd5b6814)  
) LUT6_inst7875 (
   .O(to_level3[99]),
   .I0(level4_in[594]),
   .I1(level4_in[595]),
   .I2(level4_in[596]),
   .I3(level4_in[597]),
   .I4(level4_in[598]),
   .I5(level4_in[599])
);

LUT6 #(
   .INIT(64'h76d99e3d76d99e3d)  
) LUT6_inst7876 (
   .O(to_level3[100]),
   .I0(level4_in[600]),
   .I1(level4_in[601]),
   .I2(level4_in[602]),
   .I3(level4_in[603]),
   .I4(level4_in[604]),
   .I5(level4_in[605])
);

LUT6 #(
   .INIT(64'h4014557b4014557b)  
) LUT6_inst7877 (
   .O(to_level3[101]),
   .I0(level4_in[606]),
   .I1(level4_in[607]),
   .I2(level4_in[608]),
   .I3(level4_in[609]),
   .I4(level4_in[610]),
   .I5(level4_in[611])
);

LUT6 #(
   .INIT(64'h42245d7742245d77)  
) LUT6_inst7878 (
   .O(to_level3[102]),
   .I0(level4_in[612]),
   .I1(level4_in[613]),
   .I2(level4_in[614]),
   .I3(level4_in[615]),
   .I4(level4_in[616]),
   .I5(level4_in[617])
);

LUT6 #(
   .INIT(64'he66fcc33e66fcc33)  
) LUT6_inst7879 (
   .O(to_level3[103]),
   .I0(level4_in[618]),
   .I1(level4_in[619]),
   .I2(level4_in[620]),
   .I3(level4_in[621]),
   .I4(level4_in[622]),
   .I5(level4_in[623])
);

LUT6 #(
   .INIT(64'h33ec85ca33ec85ca)  
) LUT6_inst7880 (
   .O(to_level3[104]),
   .I0(level4_in[624]),
   .I1(level4_in[625]),
   .I2(level4_in[626]),
   .I3(level4_in[627]),
   .I4(level4_in[628]),
   .I5(level4_in[629])
);

LUT6 #(
   .INIT(64'h7ebfafa07ebfafa0)  
) LUT6_inst7881 (
   .O(to_level3[105]),
   .I0(level4_in[630]),
   .I1(level4_in[631]),
   .I2(level4_in[632]),
   .I3(level4_in[633]),
   .I4(level4_in[634]),
   .I5(level4_in[635])
);

LUT6 #(
   .INIT(64'h93de6b6593de6b65)  
) LUT6_inst7882 (
   .O(to_level3[106]),
   .I0(level4_in[636]),
   .I1(level4_in[637]),
   .I2(level4_in[638]),
   .I3(level4_in[639]),
   .I4(level4_in[640]),
   .I5(level4_in[641])
);

LUT6 #(
   .INIT(64'h3d515fba3d515fba)  
) LUT6_inst7883 (
   .O(to_level3[107]),
   .I0(level4_in[642]),
   .I1(level4_in[643]),
   .I2(level4_in[644]),
   .I3(level4_in[645]),
   .I4(level4_in[646]),
   .I5(level4_in[647])
);

LUT6 #(
   .INIT(64'h266c3407266c3407)  
) LUT6_inst7884 (
   .O(to_level3[108]),
   .I0(level4_in[648]),
   .I1(level4_in[649]),
   .I2(level4_in[650]),
   .I3(level4_in[651]),
   .I4(level4_in[652]),
   .I5(level4_in[653])
);

LUT6 #(
   .INIT(64'hab93a205ab93a205)  
) LUT6_inst7885 (
   .O(to_level3[109]),
   .I0(level4_in[654]),
   .I1(level4_in[655]),
   .I2(level4_in[656]),
   .I3(level4_in[657]),
   .I4(level4_in[658]),
   .I5(level4_in[659])
);

LUT6 #(
   .INIT(64'h3638424836384248)  
) LUT6_inst7886 (
   .O(to_level3[110]),
   .I0(level4_in[660]),
   .I1(level4_in[661]),
   .I2(level4_in[662]),
   .I3(level4_in[663]),
   .I4(level4_in[664]),
   .I5(level4_in[665])
);

LUT6 #(
   .INIT(64'h36d13f2d36d13f2d)  
) LUT6_inst7887 (
   .O(to_level3[111]),
   .I0(level4_in[666]),
   .I1(level4_in[667]),
   .I2(level4_in[668]),
   .I3(level4_in[669]),
   .I4(level4_in[670]),
   .I5(level4_in[671])
);

LUT6 #(
   .INIT(64'hcbfd0da6cbfd0da6)  
) LUT6_inst7888 (
   .O(to_level3[112]),
   .I0(level4_in[672]),
   .I1(level4_in[673]),
   .I2(level4_in[674]),
   .I3(level4_in[675]),
   .I4(level4_in[676]),
   .I5(level4_in[677])
);

LUT6 #(
   .INIT(64'ha49d4a9fa49d4a9f)  
) LUT6_inst7889 (
   .O(to_level3[113]),
   .I0(level4_in[678]),
   .I1(level4_in[679]),
   .I2(level4_in[680]),
   .I3(level4_in[681]),
   .I4(level4_in[682]),
   .I5(level4_in[683])
);

LUT6 #(
   .INIT(64'h8a8b6bab8a8b6bab)  
) LUT6_inst7890 (
   .O(to_level3[114]),
   .I0(level4_in[684]),
   .I1(level4_in[685]),
   .I2(level4_in[686]),
   .I3(level4_in[687]),
   .I4(level4_in[688]),
   .I5(level4_in[689])
);

LUT6 #(
   .INIT(64'h17d9f7e217d9f7e2)  
) LUT6_inst7891 (
   .O(to_level3[115]),
   .I0(level4_in[690]),
   .I1(level4_in[691]),
   .I2(level4_in[692]),
   .I3(level4_in[693]),
   .I4(level4_in[694]),
   .I5(level4_in[695])
);

LUT6 #(
   .INIT(64'h565dbffb565dbffb)  
) LUT6_inst7892 (
   .O(to_level3[116]),
   .I0(level4_in[696]),
   .I1(level4_in[697]),
   .I2(level4_in[698]),
   .I3(level4_in[699]),
   .I4(level4_in[700]),
   .I5(level4_in[701])
);

LUT6 #(
   .INIT(64'h2ac2aee22ac2aee2)  
) LUT6_inst7893 (
   .O(to_level3[117]),
   .I0(level4_in[702]),
   .I1(level4_in[703]),
   .I2(level4_in[704]),
   .I3(level4_in[705]),
   .I4(level4_in[706]),
   .I5(level4_in[707])
);

LUT6 #(
   .INIT(64'hf428dda9f428dda9)  
) LUT6_inst7894 (
   .O(to_level3[118]),
   .I0(level4_in[708]),
   .I1(level4_in[709]),
   .I2(level4_in[710]),
   .I3(level4_in[711]),
   .I4(level4_in[712]),
   .I5(level4_in[713])
);

LUT6 #(
   .INIT(64'h1c5a9ddc1c5a9ddc)  
) LUT6_inst7895 (
   .O(to_level3[119]),
   .I0(level4_in[714]),
   .I1(level4_in[715]),
   .I2(level4_in[716]),
   .I3(level4_in[717]),
   .I4(level4_in[718]),
   .I5(level4_in[719])
);

LUT6 #(
   .INIT(64'h4d8167184d816718)  
) LUT6_inst7896 (
   .O(to_level3[120]),
   .I0(level4_in[720]),
   .I1(level4_in[721]),
   .I2(level4_in[722]),
   .I3(level4_in[723]),
   .I4(level4_in[724]),
   .I5(level4_in[725])
);

LUT6 #(
   .INIT(64'hd4107664d4107664)  
) LUT6_inst7897 (
   .O(to_level3[121]),
   .I0(level4_in[726]),
   .I1(level4_in[727]),
   .I2(level4_in[728]),
   .I3(level4_in[729]),
   .I4(level4_in[730]),
   .I5(level4_in[731])
);

LUT6 #(
   .INIT(64'h9daad82e9daad82e)  
) LUT6_inst7898 (
   .O(to_level3[122]),
   .I0(level4_in[732]),
   .I1(level4_in[733]),
   .I2(level4_in[734]),
   .I3(level4_in[735]),
   .I4(level4_in[736]),
   .I5(level4_in[737])
);

LUT6 #(
   .INIT(64'h459e55c2459e55c2)  
) LUT6_inst7899 (
   .O(to_level3[123]),
   .I0(level4_in[738]),
   .I1(level4_in[739]),
   .I2(level4_in[740]),
   .I3(level4_in[741]),
   .I4(level4_in[742]),
   .I5(level4_in[743])
);

LUT6 #(
   .INIT(64'haba8ac81aba8ac81)  
) LUT6_inst7900 (
   .O(to_level3[124]),
   .I0(level4_in[744]),
   .I1(level4_in[745]),
   .I2(level4_in[746]),
   .I3(level4_in[747]),
   .I4(level4_in[748]),
   .I5(level4_in[749])
);

LUT6 #(
   .INIT(64'h3d0ec1fb3d0ec1fb)  
) LUT6_inst7901 (
   .O(to_level3[125]),
   .I0(level4_in[750]),
   .I1(level4_in[751]),
   .I2(level4_in[752]),
   .I3(level4_in[753]),
   .I4(level4_in[754]),
   .I5(level4_in[755])
);

LUT6 #(
   .INIT(64'ha4a25ca4a4a25ca4)  
) LUT6_inst7902 (
   .O(to_level3[126]),
   .I0(level4_in[756]),
   .I1(level4_in[757]),
   .I2(level4_in[758]),
   .I3(level4_in[759]),
   .I4(level4_in[760]),
   .I5(level4_in[761])
);

LUT6 #(
   .INIT(64'ha7e80edba7e80edb)  
) LUT6_inst7903 (
   .O(to_level3[127]),
   .I0(level4_in[762]),
   .I1(level4_in[763]),
   .I2(level4_in[764]),
   .I3(level4_in[765]),
   .I4(level4_in[766]),
   .I5(level4_in[767])
);

LUT6 #(
   .INIT(64'h91f885bc91f885bc)  
) LUT6_inst7904 (
   .O(to_level3[128]),
   .I0(level4_in[768]),
   .I1(level4_in[769]),
   .I2(level4_in[770]),
   .I3(level4_in[771]),
   .I4(level4_in[772]),
   .I5(level4_in[773])
);

LUT6 #(
   .INIT(64'hc2da1e3ec2da1e3e)  
) LUT6_inst7905 (
   .O(to_level3[129]),
   .I0(level4_in[774]),
   .I1(level4_in[775]),
   .I2(level4_in[776]),
   .I3(level4_in[777]),
   .I4(level4_in[778]),
   .I5(level4_in[779])
);

LUT6 #(
   .INIT(64'h291d643a291d643a)  
) LUT6_inst7906 (
   .O(to_level3[130]),
   .I0(level4_in[780]),
   .I1(level4_in[781]),
   .I2(level4_in[782]),
   .I3(level4_in[783]),
   .I4(level4_in[784]),
   .I5(level4_in[785])
);

LUT6 #(
   .INIT(64'h1bd3c50c1bd3c50c)  
) LUT6_inst7907 (
   .O(to_level3[131]),
   .I0(level4_in[786]),
   .I1(level4_in[787]),
   .I2(level4_in[788]),
   .I3(level4_in[789]),
   .I4(level4_in[790]),
   .I5(level4_in[791])
);

LUT6 #(
   .INIT(64'h03f161ac03f161ac)  
) LUT6_inst7908 (
   .O(to_level3[132]),
   .I0(level4_in[792]),
   .I1(level4_in[793]),
   .I2(level4_in[794]),
   .I3(level4_in[795]),
   .I4(level4_in[796]),
   .I5(level4_in[797])
);

LUT6 #(
   .INIT(64'hb83d2773b83d2773)  
) LUT6_inst7909 (
   .O(to_level3[133]),
   .I0(level4_in[798]),
   .I1(level4_in[799]),
   .I2(level4_in[800]),
   .I3(level4_in[801]),
   .I4(level4_in[802]),
   .I5(level4_in[803])
);

LUT6 #(
   .INIT(64'h04fea7dd04fea7dd)  
) LUT6_inst7910 (
   .O(to_level3[134]),
   .I0(level4_in[804]),
   .I1(level4_in[805]),
   .I2(level4_in[806]),
   .I3(level4_in[807]),
   .I4(level4_in[808]),
   .I5(level4_in[809])
);

LUT6 #(
   .INIT(64'h500432fd500432fd)  
) LUT6_inst7911 (
   .O(to_level3[135]),
   .I0(level4_in[810]),
   .I1(level4_in[811]),
   .I2(level4_in[812]),
   .I3(level4_in[813]),
   .I4(level4_in[814]),
   .I5(level4_in[815])
);

LUT6 #(
   .INIT(64'hf92bf0f7f92bf0f7)  
) LUT6_inst7912 (
   .O(to_level3[136]),
   .I0(level4_in[816]),
   .I1(level4_in[817]),
   .I2(level4_in[818]),
   .I3(level4_in[819]),
   .I4(level4_in[820]),
   .I5(level4_in[821])
);

LUT6 #(
   .INIT(64'h66f5559166f55591)  
) LUT6_inst7913 (
   .O(to_level3[137]),
   .I0(level4_in[822]),
   .I1(level4_in[823]),
   .I2(level4_in[824]),
   .I3(level4_in[825]),
   .I4(level4_in[826]),
   .I5(level4_in[827])
);

LUT6 #(
   .INIT(64'h20601bd920601bd9)  
) LUT6_inst7914 (
   .O(to_level3[138]),
   .I0(level4_in[828]),
   .I1(level4_in[829]),
   .I2(level4_in[830]),
   .I3(level4_in[831]),
   .I4(level4_in[832]),
   .I5(level4_in[833])
);

LUT6 #(
   .INIT(64'h36654bd736654bd7)  
) LUT6_inst7915 (
   .O(to_level3[139]),
   .I0(level4_in[834]),
   .I1(level4_in[835]),
   .I2(level4_in[836]),
   .I3(level4_in[837]),
   .I4(level4_in[838]),
   .I5(level4_in[839])
);

LUT6 #(
   .INIT(64'h22568bd222568bd2)  
) LUT6_inst7916 (
   .O(to_level3[140]),
   .I0(level4_in[840]),
   .I1(level4_in[841]),
   .I2(level4_in[842]),
   .I3(level4_in[843]),
   .I4(level4_in[844]),
   .I5(level4_in[845])
);

LUT6 #(
   .INIT(64'h0adb49220adb4922)  
) LUT6_inst7917 (
   .O(to_level3[141]),
   .I0(level4_in[846]),
   .I1(level4_in[847]),
   .I2(level4_in[848]),
   .I3(level4_in[849]),
   .I4(level4_in[850]),
   .I5(level4_in[851])
);

LUT6 #(
   .INIT(64'h3cb81f5d3cb81f5d)  
) LUT6_inst7918 (
   .O(to_level3[142]),
   .I0(level4_in[852]),
   .I1(level4_in[853]),
   .I2(level4_in[854]),
   .I3(level4_in[855]),
   .I4(level4_in[856]),
   .I5(level4_in[857])
);

LUT6 #(
   .INIT(64'h36dc42a036dc42a0)  
) LUT6_inst7919 (
   .O(to_level3[143]),
   .I0(level4_in[858]),
   .I1(level4_in[859]),
   .I2(level4_in[860]),
   .I3(level4_in[861]),
   .I4(level4_in[862]),
   .I5(level4_in[863])
);

LUT6 #(
   .INIT(64'h4e5aaa654e5aaa65)  
) LUT6_inst7920 (
   .O(to_level3[144]),
   .I0(level4_in[864]),
   .I1(level4_in[865]),
   .I2(level4_in[866]),
   .I3(level4_in[867]),
   .I4(level4_in[868]),
   .I5(level4_in[869])
);

LUT6 #(
   .INIT(64'h8301048d8301048d)  
) LUT6_inst7921 (
   .O(to_level3[145]),
   .I0(level4_in[870]),
   .I1(level4_in[871]),
   .I2(level4_in[872]),
   .I3(level4_in[873]),
   .I4(level4_in[874]),
   .I5(level4_in[875])
);

LUT6 #(
   .INIT(64'h0d6380370d638037)  
) LUT6_inst7922 (
   .O(to_level3[146]),
   .I0(level4_in[876]),
   .I1(level4_in[877]),
   .I2(level4_in[878]),
   .I3(level4_in[879]),
   .I4(level4_in[880]),
   .I5(level4_in[881])
);

LUT6 #(
   .INIT(64'hea8514f1ea8514f1)  
) LUT6_inst7923 (
   .O(to_level3[147]),
   .I0(level4_in[882]),
   .I1(level4_in[883]),
   .I2(level4_in[884]),
   .I3(level4_in[885]),
   .I4(level4_in[886]),
   .I5(level4_in[887])
);

LUT6 #(
   .INIT(64'h04595f2604595f26)  
) LUT6_inst7924 (
   .O(to_level3[148]),
   .I0(level4_in[888]),
   .I1(level4_in[889]),
   .I2(level4_in[890]),
   .I3(level4_in[891]),
   .I4(level4_in[892]),
   .I5(level4_in[893])
);

LUT6 #(
   .INIT(64'hf8bf237bf8bf237b)  
) LUT6_inst7925 (
   .O(to_level3[149]),
   .I0(level4_in[894]),
   .I1(level4_in[895]),
   .I2(level4_in[896]),
   .I3(level4_in[897]),
   .I4(level4_in[898]),
   .I5(level4_in[899])
);

LUT6 #(
   .INIT(64'h0b2789d70b2789d7)  
) LUT6_inst7926 (
   .O(to_level3[150]),
   .I0(level4_in[900]),
   .I1(level4_in[901]),
   .I2(level4_in[902]),
   .I3(level4_in[903]),
   .I4(level4_in[904]),
   .I5(level4_in[905])
);

LUT6 #(
   .INIT(64'hb1b7ede5b1b7ede5)  
) LUT6_inst7927 (
   .O(to_level3[151]),
   .I0(level4_in[906]),
   .I1(level4_in[907]),
   .I2(level4_in[908]),
   .I3(level4_in[909]),
   .I4(level4_in[910]),
   .I5(level4_in[911])
);

LUT6 #(
   .INIT(64'hd07c1c5bd07c1c5b)  
) LUT6_inst7928 (
   .O(to_level3[152]),
   .I0(level4_in[912]),
   .I1(level4_in[913]),
   .I2(level4_in[914]),
   .I3(level4_in[915]),
   .I4(level4_in[916]),
   .I5(level4_in[917])
);

LUT6 #(
   .INIT(64'h23477f9523477f95)  
) LUT6_inst7929 (
   .O(to_level3[153]),
   .I0(level4_in[918]),
   .I1(level4_in[919]),
   .I2(level4_in[920]),
   .I3(level4_in[921]),
   .I4(level4_in[922]),
   .I5(level4_in[923])
);

LUT6 #(
   .INIT(64'hb3a2cf4cb3a2cf4c)  
) LUT6_inst7930 (
   .O(to_level3[154]),
   .I0(level4_in[924]),
   .I1(level4_in[925]),
   .I2(level4_in[926]),
   .I3(level4_in[927]),
   .I4(level4_in[928]),
   .I5(level4_in[929])
);

LUT6 #(
   .INIT(64'hf1ff5464f1ff5464)  
) LUT6_inst7931 (
   .O(to_level3[155]),
   .I0(level4_in[930]),
   .I1(level4_in[931]),
   .I2(level4_in[932]),
   .I3(level4_in[933]),
   .I4(level4_in[934]),
   .I5(level4_in[935])
);

LUT6 #(
   .INIT(64'h3f179bee3f179bee)  
) LUT6_inst7932 (
   .O(to_level3[156]),
   .I0(level4_in[936]),
   .I1(level4_in[937]),
   .I2(level4_in[938]),
   .I3(level4_in[939]),
   .I4(level4_in[940]),
   .I5(level4_in[941])
);

LUT6 #(
   .INIT(64'he1445e16e1445e16)  
) LUT6_inst7933 (
   .O(to_level3[157]),
   .I0(level4_in[942]),
   .I1(level4_in[943]),
   .I2(level4_in[944]),
   .I3(level4_in[945]),
   .I4(level4_in[946]),
   .I5(level4_in[947])
);

LUT6 #(
   .INIT(64'h86fa555686fa5556)  
) LUT6_inst7934 (
   .O(to_level3[158]),
   .I0(level4_in[948]),
   .I1(level4_in[949]),
   .I2(level4_in[950]),
   .I3(level4_in[951]),
   .I4(level4_in[952]),
   .I5(level4_in[953])
);

LUT6 #(
   .INIT(64'he2c54d09e2c54d09)  
) LUT6_inst7935 (
   .O(to_level3[159]),
   .I0(level4_in[954]),
   .I1(level4_in[955]),
   .I2(level4_in[956]),
   .I3(level4_in[957]),
   .I4(level4_in[958]),
   .I5(level4_in[959])
);

LUT6 #(
   .INIT(64'h78b3278778b32787)  
) LUT6_inst7936 (
   .O(to_level3[160]),
   .I0(level4_in[960]),
   .I1(level4_in[961]),
   .I2(level4_in[962]),
   .I3(level4_in[963]),
   .I4(level4_in[964]),
   .I5(level4_in[965])
);

LUT6 #(
   .INIT(64'hf75970d9f75970d9)  
) LUT6_inst7937 (
   .O(to_level3[161]),
   .I0(level4_in[966]),
   .I1(level4_in[967]),
   .I2(level4_in[968]),
   .I3(level4_in[969]),
   .I4(level4_in[970]),
   .I5(level4_in[971])
);

LUT6 #(
   .INIT(64'hbc1e8b65bc1e8b65)  
) LUT6_inst7938 (
   .O(to_level3[162]),
   .I0(level4_in[972]),
   .I1(level4_in[973]),
   .I2(level4_in[974]),
   .I3(level4_in[975]),
   .I4(level4_in[976]),
   .I5(level4_in[977])
);

LUT6 #(
   .INIT(64'h910738fe910738fe)  
) LUT6_inst7939 (
   .O(to_level3[163]),
   .I0(level4_in[978]),
   .I1(level4_in[979]),
   .I2(level4_in[980]),
   .I3(level4_in[981]),
   .I4(level4_in[982]),
   .I5(level4_in[983])
);

LUT6 #(
   .INIT(64'hc114644dc114644d)  
) LUT6_inst7940 (
   .O(to_level3[164]),
   .I0(level4_in[984]),
   .I1(level4_in[985]),
   .I2(level4_in[986]),
   .I3(level4_in[987]),
   .I4(level4_in[988]),
   .I5(level4_in[989])
);

LUT6 #(
   .INIT(64'hdb50e657db50e657)  
) LUT6_inst7941 (
   .O(to_level3[165]),
   .I0(level4_in[990]),
   .I1(level4_in[991]),
   .I2(level4_in[992]),
   .I3(level4_in[993]),
   .I4(level4_in[994]),
   .I5(level4_in[995])
);

LUT6 #(
   .INIT(64'h7f564b8c7f564b8c)  
) LUT6_inst7942 (
   .O(to_level3[166]),
   .I0(level4_in[996]),
   .I1(level4_in[997]),
   .I2(level4_in[998]),
   .I3(level4_in[999]),
   .I4(level4_in[1000]),
   .I5(level4_in[1001])
);

LUT6 #(
   .INIT(64'h308c021f308c021f)  
) LUT6_inst7943 (
   .O(to_level3[167]),
   .I0(level4_in[1002]),
   .I1(level4_in[1003]),
   .I2(level4_in[1004]),
   .I3(level4_in[1005]),
   .I4(level4_in[1006]),
   .I5(level4_in[1007])
);

LUT6 #(
   .INIT(64'h6705652b6705652b)  
) LUT6_inst7944 (
   .O(to_level3[168]),
   .I0(level4_in[1008]),
   .I1(level4_in[1009]),
   .I2(level4_in[1010]),
   .I3(level4_in[1011]),
   .I4(level4_in[1012]),
   .I5(level4_in[1013])
);

LUT6 #(
   .INIT(64'h095f39cd095f39cd)  
) LUT6_inst7945 (
   .O(to_level3[169]),
   .I0(level4_in[1014]),
   .I1(level4_in[1015]),
   .I2(level4_in[1016]),
   .I3(level4_in[1017]),
   .I4(level4_in[1018]),
   .I5(level4_in[1019])
);

LUT6 #(
   .INIT(64'hdc21df7bdc21df7b)  
) LUT6_inst7946 (
   .O(to_level3[170]),
   .I0(level4_in[1020]),
   .I1(level4_in[1021]),
   .I2(level4_in[1022]),
   .I3(level4_in[1023]),
   .I4(level4_in[1024]),
   .I5(level4_in[1025])
);

LUT6 #(
   .INIT(64'h9566c4c89566c4c8)  
) LUT6_inst7947 (
   .O(to_level3[171]),
   .I0(level4_in[1026]),
   .I1(level4_in[1027]),
   .I2(level4_in[1028]),
   .I3(level4_in[1029]),
   .I4(level4_in[1030]),
   .I5(level4_in[1031])
);

LUT6 #(
   .INIT(64'h5c8c98ab5c8c98ab)  
) LUT6_inst7948 (
   .O(to_level3[172]),
   .I0(level4_in[1032]),
   .I1(level4_in[1033]),
   .I2(level4_in[1034]),
   .I3(level4_in[1035]),
   .I4(level4_in[1036]),
   .I5(level4_in[1037])
);

LUT6 #(
   .INIT(64'h0361520603615206)  
) LUT6_inst7949 (
   .O(to_level3[173]),
   .I0(level4_in[1038]),
   .I1(level4_in[1039]),
   .I2(level4_in[1040]),
   .I3(level4_in[1041]),
   .I4(level4_in[1042]),
   .I5(level4_in[1043])
);

LUT6 #(
   .INIT(64'hfa09cb85fa09cb85)  
) LUT6_inst7950 (
   .O(to_level3[174]),
   .I0(level4_in[1044]),
   .I1(level4_in[1045]),
   .I2(level4_in[1046]),
   .I3(level4_in[1047]),
   .I4(level4_in[1048]),
   .I5(level4_in[1049])
);

LUT6 #(
   .INIT(64'habed4454abed4454)  
) LUT6_inst7951 (
   .O(to_level3[175]),
   .I0(level4_in[1050]),
   .I1(level4_in[1051]),
   .I2(level4_in[1052]),
   .I3(level4_in[1053]),
   .I4(level4_in[1054]),
   .I5(level4_in[1055])
);

LUT6 #(
   .INIT(64'h97b4c8f697b4c8f6)  
) LUT6_inst7952 (
   .O(to_level3[176]),
   .I0(level4_in[1056]),
   .I1(level4_in[1057]),
   .I2(level4_in[1058]),
   .I3(level4_in[1059]),
   .I4(level4_in[1060]),
   .I5(level4_in[1061])
);

LUT6 #(
   .INIT(64'h1cdc959f1cdc959f)  
) LUT6_inst7953 (
   .O(to_level3[177]),
   .I0(level4_in[1062]),
   .I1(level4_in[1063]),
   .I2(level4_in[1064]),
   .I3(level4_in[1065]),
   .I4(level4_in[1066]),
   .I5(level4_in[1067])
);

LUT6 #(
   .INIT(64'hbece30cbbece30cb)  
) LUT6_inst7954 (
   .O(to_level3[178]),
   .I0(level4_in[1068]),
   .I1(level4_in[1069]),
   .I2(level4_in[1070]),
   .I3(level4_in[1071]),
   .I4(level4_in[1072]),
   .I5(level4_in[1073])
);

LUT6 #(
   .INIT(64'h2161649021616490)  
) LUT6_inst7955 (
   .O(to_level3[179]),
   .I0(level4_in[1074]),
   .I1(level4_in[1075]),
   .I2(level4_in[1076]),
   .I3(level4_in[1077]),
   .I4(level4_in[1078]),
   .I5(level4_in[1079])
);

LUT6 #(
   .INIT(64'he0e44cf8e0e44cf8)  
) LUT6_inst7956 (
   .O(to_level3[180]),
   .I0(level4_in[1080]),
   .I1(level4_in[1081]),
   .I2(level4_in[1082]),
   .I3(level4_in[1083]),
   .I4(level4_in[1084]),
   .I5(level4_in[1085])
);

LUT6 #(
   .INIT(64'h6f3cb1756f3cb175)  
) LUT6_inst7957 (
   .O(to_level3[181]),
   .I0(level4_in[1086]),
   .I1(level4_in[1087]),
   .I2(level4_in[1088]),
   .I3(level4_in[1089]),
   .I4(level4_in[1090]),
   .I5(level4_in[1091])
);

LUT6 #(
   .INIT(64'hd73aabe2d73aabe2)  
) LUT6_inst7958 (
   .O(to_level3[182]),
   .I0(level4_in[1092]),
   .I1(level4_in[1093]),
   .I2(level4_in[1094]),
   .I3(level4_in[1095]),
   .I4(level4_in[1096]),
   .I5(level4_in[1097])
);

LUT6 #(
   .INIT(64'hcb8db3dacb8db3da)  
) LUT6_inst7959 (
   .O(to_level3[183]),
   .I0(level4_in[1098]),
   .I1(level4_in[1099]),
   .I2(level4_in[1100]),
   .I3(level4_in[1101]),
   .I4(level4_in[1102]),
   .I5(level4_in[1103])
);

LUT6 #(
   .INIT(64'h3788c93c3788c93c)  
) LUT6_inst7960 (
   .O(to_level3[184]),
   .I0(level4_in[1104]),
   .I1(level4_in[1105]),
   .I2(level4_in[1106]),
   .I3(level4_in[1107]),
   .I4(level4_in[1108]),
   .I5(level4_in[1109])
);

LUT6 #(
   .INIT(64'h2927d5a52927d5a5)  
) LUT6_inst7961 (
   .O(to_level3[185]),
   .I0(level4_in[1110]),
   .I1(level4_in[1111]),
   .I2(level4_in[1112]),
   .I3(level4_in[1113]),
   .I4(level4_in[1114]),
   .I5(level4_in[1115])
);

LUT6 #(
   .INIT(64'h157fe83d157fe83d)  
) LUT6_inst7962 (
   .O(to_level3[186]),
   .I0(level4_in[1116]),
   .I1(level4_in[1117]),
   .I2(level4_in[1118]),
   .I3(level4_in[1119]),
   .I4(level4_in[1120]),
   .I5(level4_in[1121])
);

LUT6 #(
   .INIT(64'h11d3fd6f11d3fd6f)  
) LUT6_inst7963 (
   .O(to_level3[187]),
   .I0(level4_in[1122]),
   .I1(level4_in[1123]),
   .I2(level4_in[1124]),
   .I3(level4_in[1125]),
   .I4(level4_in[1126]),
   .I5(level4_in[1127])
);

LUT6 #(
   .INIT(64'h10574ddd10574ddd)  
) LUT6_inst7964 (
   .O(to_level3[188]),
   .I0(level4_in[1128]),
   .I1(level4_in[1129]),
   .I2(level4_in[1130]),
   .I3(level4_in[1131]),
   .I4(level4_in[1132]),
   .I5(level4_in[1133])
);

LUT6 #(
   .INIT(64'h5d5d8a7e5d5d8a7e)  
) LUT6_inst7965 (
   .O(to_level3[189]),
   .I0(level4_in[1134]),
   .I1(level4_in[1135]),
   .I2(level4_in[1136]),
   .I3(level4_in[1137]),
   .I4(level4_in[1138]),
   .I5(level4_in[1139])
);

LUT6 #(
   .INIT(64'h2d974bcf2d974bcf)  
) LUT6_inst7966 (
   .O(to_level3[190]),
   .I0(level4_in[1140]),
   .I1(level4_in[1141]),
   .I2(level4_in[1142]),
   .I3(level4_in[1143]),
   .I4(level4_in[1144]),
   .I5(level4_in[1145])
);

LUT6 #(
   .INIT(64'h905d790e905d790e)  
) LUT6_inst7967 (
   .O(to_level3[191]),
   .I0(level4_in[1146]),
   .I1(level4_in[1147]),
   .I2(level4_in[1148]),
   .I3(level4_in[1149]),
   .I4(level4_in[1150]),
   .I5(level4_in[1151])
);

LUT6 #(
   .INIT(64'h21f058a921f058a9)  
) LUT6_inst7968 (
   .O(to_level3[192]),
   .I0(level4_in[1152]),
   .I1(level4_in[1153]),
   .I2(level4_in[1154]),
   .I3(level4_in[1155]),
   .I4(level4_in[1156]),
   .I5(level4_in[1157])
);

LUT6 #(
   .INIT(64'he2c3b51de2c3b51d)  
) LUT6_inst7969 (
   .O(to_level3[193]),
   .I0(level4_in[1158]),
   .I1(level4_in[1159]),
   .I2(level4_in[1160]),
   .I3(level4_in[1161]),
   .I4(level4_in[1162]),
   .I5(level4_in[1163])
);

LUT6 #(
   .INIT(64'h8a166a2e8a166a2e)  
) LUT6_inst7970 (
   .O(to_level3[194]),
   .I0(level4_in[1164]),
   .I1(level4_in[1165]),
   .I2(level4_in[1166]),
   .I3(level4_in[1167]),
   .I4(level4_in[1168]),
   .I5(level4_in[1169])
);

LUT6 #(
   .INIT(64'ha9ffeb05a9ffeb05)  
) LUT6_inst7971 (
   .O(to_level3[195]),
   .I0(level4_in[1170]),
   .I1(level4_in[1171]),
   .I2(level4_in[1172]),
   .I3(level4_in[1173]),
   .I4(level4_in[1174]),
   .I5(level4_in[1175])
);

LUT6 #(
   .INIT(64'he95ac22be95ac22b)  
) LUT6_inst7972 (
   .O(to_level3[196]),
   .I0(level4_in[1176]),
   .I1(level4_in[1177]),
   .I2(level4_in[1178]),
   .I3(level4_in[1179]),
   .I4(level4_in[1180]),
   .I5(level4_in[1181])
);

LUT6 #(
   .INIT(64'ha48ac942a48ac942)  
) LUT6_inst7973 (
   .O(to_level3[197]),
   .I0(level4_in[1182]),
   .I1(level4_in[1183]),
   .I2(level4_in[1184]),
   .I3(level4_in[1185]),
   .I4(level4_in[1186]),
   .I5(level4_in[1187])
);

LUT6 #(
   .INIT(64'hbb6663cfbb6663cf)  
) LUT6_inst7974 (
   .O(to_level3[198]),
   .I0(level4_in[1188]),
   .I1(level4_in[1189]),
   .I2(level4_in[1190]),
   .I3(level4_in[1191]),
   .I4(level4_in[1192]),
   .I5(level4_in[1193])
);

LUT6 #(
   .INIT(64'h82e345b382e345b3)  
) LUT6_inst7975 (
   .O(to_level3[199]),
   .I0(level4_in[1194]),
   .I1(level4_in[1195]),
   .I2(level4_in[1196]),
   .I3(level4_in[1197]),
   .I4(level4_in[1198]),
   .I5(level4_in[1199])
);

LUT6 #(
   .INIT(64'hb7a5e072b7a5e072)  
) LUT6_inst7976 (
   .O(to_level3[200]),
   .I0(level4_in[1200]),
   .I1(level4_in[1201]),
   .I2(level4_in[1202]),
   .I3(level4_in[1203]),
   .I4(level4_in[1204]),
   .I5(level4_in[1205])
);

LUT6 #(
   .INIT(64'h71e8868c71e8868c)  
) LUT6_inst7977 (
   .O(to_level3[201]),
   .I0(level4_in[1206]),
   .I1(level4_in[1207]),
   .I2(level4_in[1208]),
   .I3(level4_in[1209]),
   .I4(level4_in[1210]),
   .I5(level4_in[1211])
);

LUT6 #(
   .INIT(64'hf23dc376f23dc376)  
) LUT6_inst7978 (
   .O(to_level3[202]),
   .I0(level4_in[1212]),
   .I1(level4_in[1213]),
   .I2(level4_in[1214]),
   .I3(level4_in[1215]),
   .I4(level4_in[1216]),
   .I5(level4_in[1217])
);

LUT6 #(
   .INIT(64'h857f13a8857f13a8)  
) LUT6_inst7979 (
   .O(to_level3[203]),
   .I0(level4_in[1218]),
   .I1(level4_in[1219]),
   .I2(level4_in[1220]),
   .I3(level4_in[1221]),
   .I4(level4_in[1222]),
   .I5(level4_in[1223])
);

LUT6 #(
   .INIT(64'he019767be019767b)  
) LUT6_inst7980 (
   .O(to_level3[204]),
   .I0(level4_in[1224]),
   .I1(level4_in[1225]),
   .I2(level4_in[1226]),
   .I3(level4_in[1227]),
   .I4(level4_in[1228]),
   .I5(level4_in[1229])
);

LUT6 #(
   .INIT(64'hd04017cbd04017cb)  
) LUT6_inst7981 (
   .O(to_level3[205]),
   .I0(level4_in[1230]),
   .I1(level4_in[1231]),
   .I2(level4_in[1232]),
   .I3(level4_in[1233]),
   .I4(level4_in[1234]),
   .I5(level4_in[1235])
);

LUT6 #(
   .INIT(64'h985672fb985672fb)  
) LUT6_inst7982 (
   .O(to_level3[206]),
   .I0(level4_in[1236]),
   .I1(level4_in[1237]),
   .I2(level4_in[1238]),
   .I3(level4_in[1239]),
   .I4(level4_in[1240]),
   .I5(level4_in[1241])
);

LUT6 #(
   .INIT(64'ha02f3054a02f3054)  
) LUT6_inst7983 (
   .O(to_level3[207]),
   .I0(level4_in[1242]),
   .I1(level4_in[1243]),
   .I2(level4_in[1244]),
   .I3(level4_in[1245]),
   .I4(level4_in[1246]),
   .I5(level4_in[1247])
);

LUT6 #(
   .INIT(64'hb0178274b0178274)  
) LUT6_inst7984 (
   .O(to_level3[208]),
   .I0(level4_in[1248]),
   .I1(level4_in[1249]),
   .I2(level4_in[1250]),
   .I3(level4_in[1251]),
   .I4(level4_in[1252]),
   .I5(level4_in[1253])
);

LUT6 #(
   .INIT(64'h683804d0683804d0)  
) LUT6_inst7985 (
   .O(to_level3[209]),
   .I0(level4_in[1254]),
   .I1(level4_in[1255]),
   .I2(level4_in[1256]),
   .I3(level4_in[1257]),
   .I4(level4_in[1258]),
   .I5(level4_in[1259])
);

LUT6 #(
   .INIT(64'hc8b6b573c8b6b573)  
) LUT6_inst7986 (
   .O(to_level3[210]),
   .I0(level4_in[1260]),
   .I1(level4_in[1261]),
   .I2(level4_in[1262]),
   .I3(level4_in[1263]),
   .I4(level4_in[1264]),
   .I5(level4_in[1265])
);

LUT6 #(
   .INIT(64'hf8a8f1d9f8a8f1d9)  
) LUT6_inst7987 (
   .O(to_level3[211]),
   .I0(level4_in[1266]),
   .I1(level4_in[1267]),
   .I2(level4_in[1268]),
   .I3(level4_in[1269]),
   .I4(level4_in[1270]),
   .I5(level4_in[1271])
);

LUT6 #(
   .INIT(64'h3328a0ac3328a0ac)  
) LUT6_inst7988 (
   .O(to_level3[212]),
   .I0(level4_in[1272]),
   .I1(level4_in[1273]),
   .I2(level4_in[1274]),
   .I3(level4_in[1275]),
   .I4(level4_in[1276]),
   .I5(level4_in[1277])
);

LUT6 #(
   .INIT(64'ha864622ba864622b)  
) LUT6_inst7989 (
   .O(to_level3[213]),
   .I0(level4_in[1278]),
   .I1(level4_in[1279]),
   .I2(level4_in[1280]),
   .I3(level4_in[1281]),
   .I4(level4_in[1282]),
   .I5(level4_in[1283])
);

LUT6 #(
   .INIT(64'h829b4e06829b4e06)  
) LUT6_inst7990 (
   .O(to_level3[214]),
   .I0(level4_in[1284]),
   .I1(level4_in[1285]),
   .I2(level4_in[1286]),
   .I3(level4_in[1287]),
   .I4(level4_in[1288]),
   .I5(level4_in[1289])
);

LUT6 #(
   .INIT(64'h73c7fae673c7fae6)  
) LUT6_inst7991 (
   .O(to_level3[215]),
   .I0(level4_in[1290]),
   .I1(level4_in[1291]),
   .I2(level4_in[1292]),
   .I3(level4_in[1293]),
   .I4(level4_in[1294]),
   .I5(level4_in[1295])
);

LUT6 #(
   .INIT(64'h7dfea8d37dfea8d3)  
) LUT6_inst7992 (
   .O(to_level3[216]),
   .I0(level4_in[1296]),
   .I1(level4_in[1297]),
   .I2(level4_in[1298]),
   .I3(level4_in[1299]),
   .I4(level4_in[1300]),
   .I5(level4_in[1301])
);

LUT6 #(
   .INIT(64'hf1cc91bff1cc91bf)  
) LUT6_inst7993 (
   .O(to_level3[217]),
   .I0(level4_in[1302]),
   .I1(level4_in[1303]),
   .I2(level4_in[1304]),
   .I3(level4_in[1305]),
   .I4(level4_in[1306]),
   .I5(level4_in[1307])
);

LUT6 #(
   .INIT(64'hed1b4c1ced1b4c1c)  
) LUT6_inst7994 (
   .O(to_level3[218]),
   .I0(level4_in[1308]),
   .I1(level4_in[1309]),
   .I2(level4_in[1310]),
   .I3(level4_in[1311]),
   .I4(level4_in[1312]),
   .I5(level4_in[1313])
);

LUT6 #(
   .INIT(64'hdf5369eedf5369ee)  
) LUT6_inst7995 (
   .O(to_level3[219]),
   .I0(level4_in[1314]),
   .I1(level4_in[1315]),
   .I2(level4_in[1316]),
   .I3(level4_in[1317]),
   .I4(level4_in[1318]),
   .I5(level4_in[1319])
);

LUT6 #(
   .INIT(64'h5683ed595683ed59)  
) LUT6_inst7996 (
   .O(to_level3[220]),
   .I0(level4_in[1320]),
   .I1(level4_in[1321]),
   .I2(level4_in[1322]),
   .I3(level4_in[1323]),
   .I4(level4_in[1324]),
   .I5(level4_in[1325])
);

LUT6 #(
   .INIT(64'h9a535f4c9a535f4c)  
) LUT6_inst7997 (
   .O(to_level3[221]),
   .I0(level4_in[1326]),
   .I1(level4_in[1327]),
   .I2(level4_in[1328]),
   .I3(level4_in[1329]),
   .I4(level4_in[1330]),
   .I5(level4_in[1331])
);

LUT6 #(
   .INIT(64'hc2d539fcc2d539fc)  
) LUT6_inst7998 (
   .O(to_level3[222]),
   .I0(level4_in[1332]),
   .I1(level4_in[1333]),
   .I2(level4_in[1334]),
   .I3(level4_in[1335]),
   .I4(level4_in[1336]),
   .I5(level4_in[1337])
);

LUT6 #(
   .INIT(64'heb9bbcc4eb9bbcc4)  
) LUT6_inst7999 (
   .O(to_level3[223]),
   .I0(level4_in[1338]),
   .I1(level4_in[1339]),
   .I2(level4_in[1340]),
   .I3(level4_in[1341]),
   .I4(level4_in[1342]),
   .I5(level4_in[1343])
);

LUT6 #(
   .INIT(64'hc9ca325dc9ca325d)  
) LUT6_inst8000 (
   .O(to_level3[224]),
   .I0(level4_in[1344]),
   .I1(level4_in[1345]),
   .I2(level4_in[1346]),
   .I3(level4_in[1347]),
   .I4(level4_in[1348]),
   .I5(level4_in[1349])
);

LUT6 #(
   .INIT(64'hbe44e635be44e635)  
) LUT6_inst8001 (
   .O(to_level3[225]),
   .I0(level4_in[1350]),
   .I1(level4_in[1351]),
   .I2(level4_in[1352]),
   .I3(level4_in[1353]),
   .I4(level4_in[1354]),
   .I5(level4_in[1355])
);

LUT6 #(
   .INIT(64'hde4f1bafde4f1baf)  
) LUT6_inst8002 (
   .O(to_level3[226]),
   .I0(level4_in[1356]),
   .I1(level4_in[1357]),
   .I2(level4_in[1358]),
   .I3(level4_in[1359]),
   .I4(level4_in[1360]),
   .I5(level4_in[1361])
);

LUT6 #(
   .INIT(64'h4dc6d9594dc6d959)  
) LUT6_inst8003 (
   .O(to_level3[227]),
   .I0(level4_in[1362]),
   .I1(level4_in[1363]),
   .I2(level4_in[1364]),
   .I3(level4_in[1365]),
   .I4(level4_in[1366]),
   .I5(level4_in[1367])
);

LUT6 #(
   .INIT(64'h66df937066df9370)  
) LUT6_inst8004 (
   .O(to_level3[228]),
   .I0(level4_in[1368]),
   .I1(level4_in[1369]),
   .I2(level4_in[1370]),
   .I3(level4_in[1371]),
   .I4(level4_in[1372]),
   .I5(level4_in[1373])
);

LUT6 #(
   .INIT(64'h6cf3dd7e6cf3dd7e)  
) LUT6_inst8005 (
   .O(to_level3[229]),
   .I0(level4_in[1374]),
   .I1(level4_in[1375]),
   .I2(level4_in[1376]),
   .I3(level4_in[1377]),
   .I4(level4_in[1378]),
   .I5(level4_in[1379])
);

LUT6 #(
   .INIT(64'he45a288ee45a288e)  
) LUT6_inst8006 (
   .O(to_level3[230]),
   .I0(level4_in[1380]),
   .I1(level4_in[1381]),
   .I2(level4_in[1382]),
   .I3(level4_in[1383]),
   .I4(level4_in[1384]),
   .I5(level4_in[1385])
);

LUT6 #(
   .INIT(64'h8f4225f28f4225f2)  
) LUT6_inst8007 (
   .O(to_level3[231]),
   .I0(level4_in[1386]),
   .I1(level4_in[1387]),
   .I2(level4_in[1388]),
   .I3(level4_in[1389]),
   .I4(level4_in[1390]),
   .I5(level4_in[1391])
);

LUT6 #(
   .INIT(64'hf234aa25f234aa25)  
) LUT6_inst8008 (
   .O(to_level3[232]),
   .I0(level4_in[1392]),
   .I1(level4_in[1393]),
   .I2(level4_in[1394]),
   .I3(level4_in[1395]),
   .I4(level4_in[1396]),
   .I5(level4_in[1397])
);

LUT6 #(
   .INIT(64'hb8da47cab8da47ca)  
) LUT6_inst8009 (
   .O(to_level3[233]),
   .I0(level4_in[1398]),
   .I1(level4_in[1399]),
   .I2(level4_in[1400]),
   .I3(level4_in[1401]),
   .I4(level4_in[1402]),
   .I5(level4_in[1403])
);

LUT6 #(
   .INIT(64'h8ccc2ff48ccc2ff4)  
) LUT6_inst8010 (
   .O(to_level3[234]),
   .I0(level4_in[1404]),
   .I1(level4_in[1405]),
   .I2(level4_in[1406]),
   .I3(level4_in[1407]),
   .I4(level4_in[1408]),
   .I5(level4_in[1409])
);

LUT6 #(
   .INIT(64'h1fb933811fb93381)  
) LUT6_inst8011 (
   .O(to_level3[235]),
   .I0(level4_in[1410]),
   .I1(level4_in[1411]),
   .I2(level4_in[1412]),
   .I3(level4_in[1413]),
   .I4(level4_in[1414]),
   .I5(level4_in[1415])
);

LUT6 #(
   .INIT(64'hf8376e7cf8376e7c)  
) LUT6_inst8012 (
   .O(to_level3[236]),
   .I0(level4_in[1416]),
   .I1(level4_in[1417]),
   .I2(level4_in[1418]),
   .I3(level4_in[1419]),
   .I4(level4_in[1420]),
   .I5(level4_in[1421])
);

LUT6 #(
   .INIT(64'h9ba0837c9ba0837c)  
) LUT6_inst8013 (
   .O(to_level3[237]),
   .I0(level4_in[1422]),
   .I1(level4_in[1423]),
   .I2(level4_in[1424]),
   .I3(level4_in[1425]),
   .I4(level4_in[1426]),
   .I5(level4_in[1427])
);

LUT6 #(
   .INIT(64'h31b74cc831b74cc8)  
) LUT6_inst8014 (
   .O(to_level3[238]),
   .I0(level4_in[1428]),
   .I1(level4_in[1429]),
   .I2(level4_in[1430]),
   .I3(level4_in[1431]),
   .I4(level4_in[1432]),
   .I5(level4_in[1433])
);

LUT6 #(
   .INIT(64'h5fcb4fcb5fcb4fcb)  
) LUT6_inst8015 (
   .O(to_level3[239]),
   .I0(level4_in[1434]),
   .I1(level4_in[1435]),
   .I2(level4_in[1436]),
   .I3(level4_in[1437]),
   .I4(level4_in[1438]),
   .I5(level4_in[1439])
);

LUT6 #(
   .INIT(64'hd39b0218d39b0218)  
) LUT6_inst8016 (
   .O(to_level3[240]),
   .I0(level4_in[1440]),
   .I1(level4_in[1441]),
   .I2(level4_in[1442]),
   .I3(level4_in[1443]),
   .I4(level4_in[1444]),
   .I5(level4_in[1445])
);

LUT6 #(
   .INIT(64'hb2207d8ab2207d8a)  
) LUT6_inst8017 (
   .O(to_level3[241]),
   .I0(level4_in[1446]),
   .I1(level4_in[1447]),
   .I2(level4_in[1448]),
   .I3(level4_in[1449]),
   .I4(level4_in[1450]),
   .I5(level4_in[1451])
);

LUT6 #(
   .INIT(64'h5374297853742978)  
) LUT6_inst8018 (
   .O(to_level3[242]),
   .I0(level4_in[1452]),
   .I1(level4_in[1453]),
   .I2(level4_in[1454]),
   .I3(level4_in[1455]),
   .I4(level4_in[1456]),
   .I5(level4_in[1457])
);

LUT6 #(
   .INIT(64'h8862e5f48862e5f4)  
) LUT6_inst8019 (
   .O(to_level3[243]),
   .I0(level4_in[1458]),
   .I1(level4_in[1459]),
   .I2(level4_in[1460]),
   .I3(level4_in[1461]),
   .I4(level4_in[1462]),
   .I5(level4_in[1463])
);

LUT6 #(
   .INIT(64'h0830755c0830755c)  
) LUT6_inst8020 (
   .O(to_level3[244]),
   .I0(level4_in[1464]),
   .I1(level4_in[1465]),
   .I2(level4_in[1466]),
   .I3(level4_in[1467]),
   .I4(level4_in[1468]),
   .I5(level4_in[1469])
);

LUT6 #(
   .INIT(64'hee506f98ee506f98)  
) LUT6_inst8021 (
   .O(to_level3[245]),
   .I0(level4_in[1470]),
   .I1(level4_in[1471]),
   .I2(level4_in[1472]),
   .I3(level4_in[1473]),
   .I4(level4_in[1474]),
   .I5(level4_in[1475])
);

LUT6 #(
   .INIT(64'h47449c4c47449c4c)  
) LUT6_inst8022 (
   .O(to_level3[246]),
   .I0(level4_in[1476]),
   .I1(level4_in[1477]),
   .I2(level4_in[1478]),
   .I3(level4_in[1479]),
   .I4(level4_in[1480]),
   .I5(level4_in[1481])
);

LUT6 #(
   .INIT(64'hc49efb23c49efb23)  
) LUT6_inst8023 (
   .O(to_level3[247]),
   .I0(level4_in[1482]),
   .I1(level4_in[1483]),
   .I2(level4_in[1484]),
   .I3(level4_in[1485]),
   .I4(level4_in[1486]),
   .I5(level4_in[1487])
);

LUT6 #(
   .INIT(64'hbde9c34cbde9c34c)  
) LUT6_inst8024 (
   .O(to_level3[248]),
   .I0(level4_in[1488]),
   .I1(level4_in[1489]),
   .I2(level4_in[1490]),
   .I3(level4_in[1491]),
   .I4(level4_in[1492]),
   .I5(level4_in[1493])
);

LUT6 #(
   .INIT(64'hc55edcfbc55edcfb)  
) LUT6_inst8025 (
   .O(to_level3[249]),
   .I0(level4_in[1494]),
   .I1(level4_in[1495]),
   .I2(level4_in[1496]),
   .I3(level4_in[1497]),
   .I4(level4_in[1498]),
   .I5(level4_in[1499])
);

LUT6 #(
   .INIT(64'h46d1160246d11602)  
) LUT6_inst8026 (
   .O(to_level3[250]),
   .I0(level4_in[1500]),
   .I1(level4_in[1501]),
   .I2(level4_in[1502]),
   .I3(level4_in[1503]),
   .I4(level4_in[1504]),
   .I5(level4_in[1505])
);

LUT6 #(
   .INIT(64'h449ac3eb449ac3eb)  
) LUT6_inst8027 (
   .O(to_level3[251]),
   .I0(level4_in[1506]),
   .I1(level4_in[1507]),
   .I2(level4_in[1508]),
   .I3(level4_in[1509]),
   .I4(level4_in[1510]),
   .I5(level4_in[1511])
);

LUT6 #(
   .INIT(64'h2dd5949a2dd5949a)  
) LUT6_inst8028 (
   .O(to_level3[252]),
   .I0(level4_in[1512]),
   .I1(level4_in[1513]),
   .I2(level4_in[1514]),
   .I3(level4_in[1515]),
   .I4(level4_in[1516]),
   .I5(level4_in[1517])
);

LUT6 #(
   .INIT(64'hd260f7aad260f7aa)  
) LUT6_inst8029 (
   .O(to_level3[253]),
   .I0(level4_in[1518]),
   .I1(level4_in[1519]),
   .I2(level4_in[1520]),
   .I3(level4_in[1521]),
   .I4(level4_in[1522]),
   .I5(level4_in[1523])
);

LUT6 #(
   .INIT(64'h6ebd67256ebd6725)  
) LUT6_inst8030 (
   .O(to_level3[254]),
   .I0(level4_in[1524]),
   .I1(level4_in[1525]),
   .I2(level4_in[1526]),
   .I3(level4_in[1527]),
   .I4(level4_in[1528]),
   .I5(level4_in[1529])
);

LUT6 #(
   .INIT(64'hfcc93f95fcc93f95)  
) LUT6_inst8031 (
   .O(to_level3[255]),
   .I0(level4_in[1530]),
   .I1(level4_in[1531]),
   .I2(level4_in[1532]),
   .I3(level4_in[1533]),
   .I4(level4_in[1534]),
   .I5(level4_in[1535])
);

LUT6 #(
   .INIT(64'h774cee9c774cee9c)  
) LUT6_inst8032 (
   .O(to_level3[256]),
   .I0(level4_in[1536]),
   .I1(level4_in[1537]),
   .I2(level4_in[1538]),
   .I3(level4_in[1539]),
   .I4(level4_in[1540]),
   .I5(level4_in[1541])
);

LUT6 #(
   .INIT(64'h84052d3b84052d3b)  
) LUT6_inst8033 (
   .O(to_level3[257]),
   .I0(level4_in[1542]),
   .I1(level4_in[1543]),
   .I2(level4_in[1544]),
   .I3(level4_in[1545]),
   .I4(level4_in[1546]),
   .I5(level4_in[1547])
);

LUT6 #(
   .INIT(64'hb0d5b9e2b0d5b9e2)  
) LUT6_inst8034 (
   .O(to_level3[258]),
   .I0(level4_in[1548]),
   .I1(level4_in[1549]),
   .I2(level4_in[1550]),
   .I3(level4_in[1551]),
   .I4(level4_in[1552]),
   .I5(level4_in[1553])
);

LUT6 #(
   .INIT(64'ha7a55a06a7a55a06)  
) LUT6_inst8035 (
   .O(to_level3[259]),
   .I0(level4_in[1554]),
   .I1(level4_in[1555]),
   .I2(level4_in[1556]),
   .I3(level4_in[1557]),
   .I4(level4_in[1558]),
   .I5(level4_in[1559])
);

LUT6 #(
   .INIT(64'h81bc024681bc0246)  
) LUT6_inst8036 (
   .O(to_level3[260]),
   .I0(level4_in[1560]),
   .I1(level4_in[1561]),
   .I2(level4_in[1562]),
   .I3(level4_in[1563]),
   .I4(level4_in[1564]),
   .I5(level4_in[1565])
);

LUT6 #(
   .INIT(64'h2db54ae52db54ae5)  
) LUT6_inst8037 (
   .O(to_level3[261]),
   .I0(level4_in[1566]),
   .I1(level4_in[1567]),
   .I2(level4_in[1568]),
   .I3(level4_in[1569]),
   .I4(level4_in[1570]),
   .I5(level4_in[1571])
);

LUT6 #(
   .INIT(64'h332a8516332a8516)  
) LUT6_inst8038 (
   .O(to_level3[262]),
   .I0(level4_in[1572]),
   .I1(level4_in[1573]),
   .I2(level4_in[1574]),
   .I3(level4_in[1575]),
   .I4(level4_in[1576]),
   .I5(level4_in[1577])
);

LUT6 #(
   .INIT(64'h41d3bdf641d3bdf6)  
) LUT6_inst8039 (
   .O(to_level3[263]),
   .I0(level4_in[1578]),
   .I1(level4_in[1579]),
   .I2(level4_in[1580]),
   .I3(level4_in[1581]),
   .I4(level4_in[1582]),
   .I5(level4_in[1583])
);

LUT6 #(
   .INIT(64'h44bdcd3d44bdcd3d)  
) LUT6_inst8040 (
   .O(to_level3[264]),
   .I0(level4_in[1584]),
   .I1(level4_in[1585]),
   .I2(level4_in[1586]),
   .I3(level4_in[1587]),
   .I4(level4_in[1588]),
   .I5(level4_in[1589])
);

LUT6 #(
   .INIT(64'h075f94b0075f94b0)  
) LUT6_inst8041 (
   .O(to_level3[265]),
   .I0(level4_in[1590]),
   .I1(level4_in[1591]),
   .I2(level4_in[1592]),
   .I3(level4_in[1593]),
   .I4(level4_in[1594]),
   .I5(level4_in[1595])
);

LUT6 #(
   .INIT(64'ha3eafd1da3eafd1d)  
) LUT6_inst8042 (
   .O(to_level3[266]),
   .I0(level4_in[1596]),
   .I1(level4_in[1597]),
   .I2(level4_in[1598]),
   .I3(level4_in[1599]),
   .I4(level4_in[1600]),
   .I5(level4_in[1601])
);

LUT6 #(
   .INIT(64'h7d3f5d8c7d3f5d8c)  
) LUT6_inst8043 (
   .O(to_level3[267]),
   .I0(level4_in[1602]),
   .I1(level4_in[1603]),
   .I2(level4_in[1604]),
   .I3(level4_in[1605]),
   .I4(level4_in[1606]),
   .I5(level4_in[1607])
);

LUT6 #(
   .INIT(64'h9cff6bc89cff6bc8)  
) LUT6_inst8044 (
   .O(to_level3[268]),
   .I0(level4_in[1608]),
   .I1(level4_in[1609]),
   .I2(level4_in[1610]),
   .I3(level4_in[1611]),
   .I4(level4_in[1612]),
   .I5(level4_in[1613])
);

LUT6 #(
   .INIT(64'h5ebcde335ebcde33)  
) LUT6_inst8045 (
   .O(to_level3[269]),
   .I0(level4_in[1614]),
   .I1(level4_in[1615]),
   .I2(level4_in[1616]),
   .I3(level4_in[1617]),
   .I4(level4_in[1618]),
   .I5(level4_in[1619])
);

LUT6 #(
   .INIT(64'hef596418ef596418)  
) LUT6_inst8046 (
   .O(to_level3[270]),
   .I0(level4_in[1620]),
   .I1(level4_in[1621]),
   .I2(level4_in[1622]),
   .I3(level4_in[1623]),
   .I4(level4_in[1624]),
   .I5(level4_in[1625])
);

LUT6 #(
   .INIT(64'hc2cdadb1c2cdadb1)  
) LUT6_inst8047 (
   .O(to_level3[271]),
   .I0(level4_in[1626]),
   .I1(level4_in[1627]),
   .I2(level4_in[1628]),
   .I3(level4_in[1629]),
   .I4(level4_in[1630]),
   .I5(level4_in[1631])
);

LUT6 #(
   .INIT(64'h1c7c71dd1c7c71dd)  
) LUT6_inst8048 (
   .O(to_level3[272]),
   .I0(level4_in[1632]),
   .I1(level4_in[1633]),
   .I2(level4_in[1634]),
   .I3(level4_in[1635]),
   .I4(level4_in[1636]),
   .I5(level4_in[1637])
);

LUT6 #(
   .INIT(64'h12ed1aa612ed1aa6)  
) LUT6_inst8049 (
   .O(to_level3[273]),
   .I0(level4_in[1638]),
   .I1(level4_in[1639]),
   .I2(level4_in[1640]),
   .I3(level4_in[1641]),
   .I4(level4_in[1642]),
   .I5(level4_in[1643])
);

LUT6 #(
   .INIT(64'h8b0387d38b0387d3)  
) LUT6_inst8050 (
   .O(to_level3[274]),
   .I0(level4_in[1644]),
   .I1(level4_in[1645]),
   .I2(level4_in[1646]),
   .I3(level4_in[1647]),
   .I4(level4_in[1648]),
   .I5(level4_in[1649])
);

LUT6 #(
   .INIT(64'hdaaa5a0ddaaa5a0d)  
) LUT6_inst8051 (
   .O(to_level3[275]),
   .I0(level4_in[1650]),
   .I1(level4_in[1651]),
   .I2(level4_in[1652]),
   .I3(level4_in[1653]),
   .I4(level4_in[1654]),
   .I5(level4_in[1655])
);

LUT6 #(
   .INIT(64'h7924f4127924f412)  
) LUT6_inst8052 (
   .O(to_level3[276]),
   .I0(level4_in[1656]),
   .I1(level4_in[1657]),
   .I2(level4_in[1658]),
   .I3(level4_in[1659]),
   .I4(level4_in[1660]),
   .I5(level4_in[1661])
);

LUT6 #(
   .INIT(64'h3a3bc2e43a3bc2e4)  
) LUT6_inst8053 (
   .O(to_level3[277]),
   .I0(level4_in[1662]),
   .I1(level4_in[1663]),
   .I2(level4_in[1664]),
   .I3(level4_in[1665]),
   .I4(level4_in[1666]),
   .I5(level4_in[1667])
);

LUT6 #(
   .INIT(64'h2f8ebedf2f8ebedf)  
) LUT6_inst8054 (
   .O(to_level3[278]),
   .I0(level4_in[1668]),
   .I1(level4_in[1669]),
   .I2(level4_in[1670]),
   .I3(level4_in[1671]),
   .I4(level4_in[1672]),
   .I5(level4_in[1673])
);

LUT6 #(
   .INIT(64'hf62cb0baf62cb0ba)  
) LUT6_inst8055 (
   .O(to_level3[279]),
   .I0(level4_in[1674]),
   .I1(level4_in[1675]),
   .I2(level4_in[1676]),
   .I3(level4_in[1677]),
   .I4(level4_in[1678]),
   .I5(level4_in[1679])
);

LUT6 #(
   .INIT(64'h2f5264cf2f5264cf)  
) LUT6_inst8056 (
   .O(to_level3[280]),
   .I0(level4_in[1680]),
   .I1(level4_in[1681]),
   .I2(level4_in[1682]),
   .I3(level4_in[1683]),
   .I4(level4_in[1684]),
   .I5(level4_in[1685])
);

LUT6 #(
   .INIT(64'haff8d175aff8d175)  
) LUT6_inst8057 (
   .O(to_level3[281]),
   .I0(level4_in[1686]),
   .I1(level4_in[1687]),
   .I2(level4_in[1688]),
   .I3(level4_in[1689]),
   .I4(level4_in[1690]),
   .I5(level4_in[1691])
);

LUT6 #(
   .INIT(64'h3aa9701a3aa9701a)  
) LUT6_inst8058 (
   .O(to_level3[282]),
   .I0(level4_in[1692]),
   .I1(level4_in[1693]),
   .I2(level4_in[1694]),
   .I3(level4_in[1695]),
   .I4(level4_in[1696]),
   .I5(level4_in[1697])
);

LUT6 #(
   .INIT(64'h9ab135b09ab135b0)  
) LUT6_inst8059 (
   .O(to_level3[283]),
   .I0(level4_in[1698]),
   .I1(level4_in[1699]),
   .I2(level4_in[1700]),
   .I3(level4_in[1701]),
   .I4(level4_in[1702]),
   .I5(level4_in[1703])
);

LUT6 #(
   .INIT(64'had577dcbad577dcb)  
) LUT6_inst8060 (
   .O(to_level3[284]),
   .I0(level4_in[1704]),
   .I1(level4_in[1705]),
   .I2(level4_in[1706]),
   .I3(level4_in[1707]),
   .I4(level4_in[1708]),
   .I5(level4_in[1709])
);

LUT6 #(
   .INIT(64'h2fae8ca32fae8ca3)  
) LUT6_inst8061 (
   .O(to_level3[285]),
   .I0(level4_in[1710]),
   .I1(level4_in[1711]),
   .I2(level4_in[1712]),
   .I3(level4_in[1713]),
   .I4(level4_in[1714]),
   .I5(level4_in[1715])
);

LUT6 #(
   .INIT(64'h3c5ae0653c5ae065)  
) LUT6_inst8062 (
   .O(to_level3[286]),
   .I0(level4_in[1716]),
   .I1(level4_in[1717]),
   .I2(level4_in[1718]),
   .I3(level4_in[1719]),
   .I4(level4_in[1720]),
   .I5(level4_in[1721])
);

LUT6 #(
   .INIT(64'hdef0fd7bdef0fd7b)  
) LUT6_inst8063 (
   .O(to_level3[287]),
   .I0(level4_in[1722]),
   .I1(level4_in[1723]),
   .I2(level4_in[1724]),
   .I3(level4_in[1725]),
   .I4(level4_in[1726]),
   .I5(level4_in[1727])
);

LUT6 #(
   .INIT(64'h47be87a047be87a0)  
) LUT6_inst8064 (
   .O(to_level3[288]),
   .I0(level4_in[1728]),
   .I1(level4_in[1729]),
   .I2(level4_in[1730]),
   .I3(level4_in[1731]),
   .I4(level4_in[1732]),
   .I5(level4_in[1733])
);

LUT6 #(
   .INIT(64'h6e0195496e019549)  
) LUT6_inst8065 (
   .O(to_level3[289]),
   .I0(level4_in[1734]),
   .I1(level4_in[1735]),
   .I2(level4_in[1736]),
   .I3(level4_in[1737]),
   .I4(level4_in[1738]),
   .I5(level4_in[1739])
);

LUT6 #(
   .INIT(64'h4bb06d214bb06d21)  
) LUT6_inst8066 (
   .O(to_level3[290]),
   .I0(level4_in[1740]),
   .I1(level4_in[1741]),
   .I2(level4_in[1742]),
   .I3(level4_in[1743]),
   .I4(level4_in[1744]),
   .I5(level4_in[1745])
);

LUT6 #(
   .INIT(64'hf0a85936f0a85936)  
) LUT6_inst8067 (
   .O(to_level3[291]),
   .I0(level4_in[1746]),
   .I1(level4_in[1747]),
   .I2(level4_in[1748]),
   .I3(level4_in[1749]),
   .I4(level4_in[1750]),
   .I5(level4_in[1751])
);

LUT6 #(
   .INIT(64'h461b28b6461b28b6)  
) LUT6_inst8068 (
   .O(to_level3[292]),
   .I0(level4_in[1752]),
   .I1(level4_in[1753]),
   .I2(level4_in[1754]),
   .I3(level4_in[1755]),
   .I4(level4_in[1756]),
   .I5(level4_in[1757])
);

LUT6 #(
   .INIT(64'h03fb2bd103fb2bd1)  
) LUT6_inst8069 (
   .O(to_level3[293]),
   .I0(level4_in[1758]),
   .I1(level4_in[1759]),
   .I2(level4_in[1760]),
   .I3(level4_in[1761]),
   .I4(level4_in[1762]),
   .I5(level4_in[1763])
);

LUT6 #(
   .INIT(64'ha302d37ea302d37e)  
) LUT6_inst8070 (
   .O(to_level3[294]),
   .I0(level4_in[1764]),
   .I1(level4_in[1765]),
   .I2(level4_in[1766]),
   .I3(level4_in[1767]),
   .I4(level4_in[1768]),
   .I5(level4_in[1769])
);

LUT6 #(
   .INIT(64'he2b126dae2b126da)  
) LUT6_inst8071 (
   .O(to_level3[295]),
   .I0(level4_in[1770]),
   .I1(level4_in[1771]),
   .I2(level4_in[1772]),
   .I3(level4_in[1773]),
   .I4(level4_in[1774]),
   .I5(level4_in[1775])
);

LUT6 #(
   .INIT(64'hd56953d5d56953d5)  
) LUT6_inst8072 (
   .O(to_level3[296]),
   .I0(level4_in[1776]),
   .I1(level4_in[1777]),
   .I2(level4_in[1778]),
   .I3(level4_in[1779]),
   .I4(level4_in[1780]),
   .I5(level4_in[1781])
);

LUT6 #(
   .INIT(64'h8a51b8888a51b888)  
) LUT6_inst8073 (
   .O(to_level3[297]),
   .I0(level4_in[1782]),
   .I1(level4_in[1783]),
   .I2(level4_in[1784]),
   .I3(level4_in[1785]),
   .I4(level4_in[1786]),
   .I5(level4_in[1787])
);

LUT6 #(
   .INIT(64'h82b069fe82b069fe)  
) LUT6_inst8074 (
   .O(to_level3[298]),
   .I0(level4_in[1788]),
   .I1(level4_in[1789]),
   .I2(level4_in[1790]),
   .I3(level4_in[1791]),
   .I4(level4_in[1792]),
   .I5(level4_in[1793])
);

LUT6 #(
   .INIT(64'hba3a9cd5ba3a9cd5)  
) LUT6_inst8075 (
   .O(to_level3[299]),
   .I0(level4_in[1794]),
   .I1(level4_in[1795]),
   .I2(level4_in[1796]),
   .I3(level4_in[1797]),
   .I4(level4_in[1798]),
   .I5(level4_in[1799])
);

LUT6 #(
   .INIT(64'hf88ca589f88ca589)  
) LUT6_inst8076 (
   .O(to_level3[300]),
   .I0(level4_in[1800]),
   .I1(level4_in[1801]),
   .I2(level4_in[1802]),
   .I3(level4_in[1803]),
   .I4(level4_in[1804]),
   .I5(level4_in[1805])
);

LUT6 #(
   .INIT(64'h437e3438437e3438)  
) LUT6_inst8077 (
   .O(to_level3[301]),
   .I0(level4_in[1806]),
   .I1(level4_in[1807]),
   .I2(level4_in[1808]),
   .I3(level4_in[1809]),
   .I4(level4_in[1810]),
   .I5(level4_in[1811])
);

LUT6 #(
   .INIT(64'hdc53d503dc53d503)  
) LUT6_inst8078 (
   .O(to_level3[302]),
   .I0(level4_in[1812]),
   .I1(level4_in[1813]),
   .I2(level4_in[1814]),
   .I3(level4_in[1815]),
   .I4(level4_in[1816]),
   .I5(level4_in[1817])
);

LUT6 #(
   .INIT(64'h226d6241226d6241)  
) LUT6_inst8079 (
   .O(to_level3[303]),
   .I0(level4_in[1818]),
   .I1(level4_in[1819]),
   .I2(level4_in[1820]),
   .I3(level4_in[1821]),
   .I4(level4_in[1822]),
   .I5(level4_in[1823])
);

LUT6 #(
   .INIT(64'h92b2dafb92b2dafb)  
) LUT6_inst8080 (
   .O(to_level3[304]),
   .I0(level4_in[1824]),
   .I1(level4_in[1825]),
   .I2(level4_in[1826]),
   .I3(level4_in[1827]),
   .I4(level4_in[1828]),
   .I5(level4_in[1829])
);

LUT6 #(
   .INIT(64'h9489e4609489e460)  
) LUT6_inst8081 (
   .O(to_level3[305]),
   .I0(level4_in[1830]),
   .I1(level4_in[1831]),
   .I2(level4_in[1832]),
   .I3(level4_in[1833]),
   .I4(level4_in[1834]),
   .I5(level4_in[1835])
);

LUT6 #(
   .INIT(64'h789c17c0789c17c0)  
) LUT6_inst8082 (
   .O(to_level3[306]),
   .I0(level4_in[1836]),
   .I1(level4_in[1837]),
   .I2(level4_in[1838]),
   .I3(level4_in[1839]),
   .I4(level4_in[1840]),
   .I5(level4_in[1841])
);

LUT6 #(
   .INIT(64'h19ba7a1d19ba7a1d)  
) LUT6_inst8083 (
   .O(to_level3[307]),
   .I0(level4_in[1842]),
   .I1(level4_in[1843]),
   .I2(level4_in[1844]),
   .I3(level4_in[1845]),
   .I4(level4_in[1846]),
   .I5(level4_in[1847])
);

LUT6 #(
   .INIT(64'haf304917af304917)  
) LUT6_inst8084 (
   .O(to_level3[308]),
   .I0(level4_in[1848]),
   .I1(level4_in[1849]),
   .I2(level4_in[1850]),
   .I3(level4_in[1851]),
   .I4(level4_in[1852]),
   .I5(level4_in[1853])
);

LUT6 #(
   .INIT(64'hb71ea72ab71ea72a)  
) LUT6_inst8085 (
   .O(to_level3[309]),
   .I0(level4_in[1854]),
   .I1(level4_in[1855]),
   .I2(level4_in[1856]),
   .I3(level4_in[1857]),
   .I4(level4_in[1858]),
   .I5(level4_in[1859])
);

LUT6 #(
   .INIT(64'h4565bec84565bec8)  
) LUT6_inst8086 (
   .O(to_level3[310]),
   .I0(level4_in[1860]),
   .I1(level4_in[1861]),
   .I2(level4_in[1862]),
   .I3(level4_in[1863]),
   .I4(level4_in[1864]),
   .I5(level4_in[1865])
);

LUT6 #(
   .INIT(64'h149b53b5149b53b5)  
) LUT6_inst8087 (
   .O(to_level3[311]),
   .I0(level4_in[1866]),
   .I1(level4_in[1867]),
   .I2(level4_in[1868]),
   .I3(level4_in[1869]),
   .I4(level4_in[1870]),
   .I5(level4_in[1871])
);

LUT6 #(
   .INIT(64'hde838557de838557)  
) LUT6_inst8088 (
   .O(to_level3[312]),
   .I0(level4_in[1872]),
   .I1(level4_in[1873]),
   .I2(level4_in[1874]),
   .I3(level4_in[1875]),
   .I4(level4_in[1876]),
   .I5(level4_in[1877])
);

LUT6 #(
   .INIT(64'hb8b39b56b8b39b56)  
) LUT6_inst8089 (
   .O(to_level3[313]),
   .I0(level4_in[1878]),
   .I1(level4_in[1879]),
   .I2(level4_in[1880]),
   .I3(level4_in[1881]),
   .I4(level4_in[1882]),
   .I5(level4_in[1883])
);

LUT6 #(
   .INIT(64'h02cf848e02cf848e)  
) LUT6_inst8090 (
   .O(to_level3[314]),
   .I0(level4_in[1884]),
   .I1(level4_in[1885]),
   .I2(level4_in[1886]),
   .I3(level4_in[1887]),
   .I4(level4_in[1888]),
   .I5(level4_in[1889])
);

LUT6 #(
   .INIT(64'hdbd3d747dbd3d747)  
) LUT6_inst8091 (
   .O(to_level3[315]),
   .I0(level4_in[1890]),
   .I1(level4_in[1891]),
   .I2(level4_in[1892]),
   .I3(level4_in[1893]),
   .I4(level4_in[1894]),
   .I5(level4_in[1895])
);

LUT6 #(
   .INIT(64'he232a0e7e232a0e7)  
) LUT6_inst8092 (
   .O(to_level3[316]),
   .I0(level4_in[1896]),
   .I1(level4_in[1897]),
   .I2(level4_in[1898]),
   .I3(level4_in[1899]),
   .I4(level4_in[1900]),
   .I5(level4_in[1901])
);

LUT6 #(
   .INIT(64'hbb372960bb372960)  
) LUT6_inst8093 (
   .O(to_level3[317]),
   .I0(level4_in[1902]),
   .I1(level4_in[1903]),
   .I2(level4_in[1904]),
   .I3(level4_in[1905]),
   .I4(level4_in[1906]),
   .I5(level4_in[1907])
);

LUT6 #(
   .INIT(64'h46e5ded646e5ded6)  
) LUT6_inst8094 (
   .O(to_level3[318]),
   .I0(level4_in[1908]),
   .I1(level4_in[1909]),
   .I2(level4_in[1910]),
   .I3(level4_in[1911]),
   .I4(level4_in[1912]),
   .I5(level4_in[1913])
);

LUT6 #(
   .INIT(64'hcb4b2091cb4b2091)  
) LUT6_inst8095 (
   .O(to_level3[319]),
   .I0(level4_in[1914]),
   .I1(level4_in[1915]),
   .I2(level4_in[1916]),
   .I3(level4_in[1917]),
   .I4(level4_in[1918]),
   .I5(level4_in[1919])
);

LUT6 #(
   .INIT(64'h731b36a4731b36a4)  
) LUT6_inst8096 (
   .O(to_level3[320]),
   .I0(level4_in[1920]),
   .I1(level4_in[1921]),
   .I2(level4_in[1922]),
   .I3(level4_in[1923]),
   .I4(level4_in[1924]),
   .I5(level4_in[1925])
);

LUT6 #(
   .INIT(64'h9680687896806878)  
) LUT6_inst8097 (
   .O(to_level3[321]),
   .I0(level4_in[1926]),
   .I1(level4_in[1927]),
   .I2(level4_in[1928]),
   .I3(level4_in[1929]),
   .I4(level4_in[1930]),
   .I5(level4_in[1931])
);

LUT6 #(
   .INIT(64'haa3a5186aa3a5186)  
) LUT6_inst8098 (
   .O(to_level3[322]),
   .I0(level4_in[1932]),
   .I1(level4_in[1933]),
   .I2(level4_in[1934]),
   .I3(level4_in[1935]),
   .I4(level4_in[1936]),
   .I5(level4_in[1937])
);

LUT6 #(
   .INIT(64'h34e8100134e81001)  
) LUT6_inst8099 (
   .O(to_level3[323]),
   .I0(level4_in[1938]),
   .I1(level4_in[1939]),
   .I2(level4_in[1940]),
   .I3(level4_in[1941]),
   .I4(level4_in[1942]),
   .I5(level4_in[1943])
);

LUT6 #(
   .INIT(64'hed1611faed1611fa)  
) LUT6_inst8100 (
   .O(to_level3[324]),
   .I0(level4_in[1944]),
   .I1(level4_in[1945]),
   .I2(level4_in[1946]),
   .I3(level4_in[1947]),
   .I4(level4_in[1948]),
   .I5(level4_in[1949])
);

LUT6 #(
   .INIT(64'h35ce994c35ce994c)  
) LUT6_inst8101 (
   .O(to_level3[325]),
   .I0(level4_in[1950]),
   .I1(level4_in[1951]),
   .I2(level4_in[1952]),
   .I3(level4_in[1953]),
   .I4(level4_in[1954]),
   .I5(level4_in[1955])
);

LUT6 #(
   .INIT(64'h7d2a1cc17d2a1cc1)  
) LUT6_inst8102 (
   .O(to_level3[326]),
   .I0(level4_in[1956]),
   .I1(level4_in[1957]),
   .I2(level4_in[1958]),
   .I3(level4_in[1959]),
   .I4(level4_in[1960]),
   .I5(level4_in[1961])
);

LUT6 #(
   .INIT(64'h9cf48ac89cf48ac8)  
) LUT6_inst8103 (
   .O(to_level3[327]),
   .I0(level4_in[1962]),
   .I1(level4_in[1963]),
   .I2(level4_in[1964]),
   .I3(level4_in[1965]),
   .I4(level4_in[1966]),
   .I5(level4_in[1967])
);

LUT6 #(
   .INIT(64'hb1528617b1528617)  
) LUT6_inst8104 (
   .O(to_level3[328]),
   .I0(level4_in[1968]),
   .I1(level4_in[1969]),
   .I2(level4_in[1970]),
   .I3(level4_in[1971]),
   .I4(level4_in[1972]),
   .I5(level4_in[1973])
);

LUT6 #(
   .INIT(64'h4829ad5c4829ad5c)  
) LUT6_inst8105 (
   .O(to_level3[329]),
   .I0(level4_in[1974]),
   .I1(level4_in[1975]),
   .I2(level4_in[1976]),
   .I3(level4_in[1977]),
   .I4(level4_in[1978]),
   .I5(level4_in[1979])
);

LUT6 #(
   .INIT(64'h32689baf32689baf)  
) LUT6_inst8106 (
   .O(to_level3[330]),
   .I0(level4_in[1980]),
   .I1(level4_in[1981]),
   .I2(level4_in[1982]),
   .I3(level4_in[1983]),
   .I4(level4_in[1984]),
   .I5(level4_in[1985])
);

LUT6 #(
   .INIT(64'h0fb41a840fb41a84)  
) LUT6_inst8107 (
   .O(to_level3[331]),
   .I0(level4_in[1986]),
   .I1(level4_in[1987]),
   .I2(level4_in[1988]),
   .I3(level4_in[1989]),
   .I4(level4_in[1990]),
   .I5(level4_in[1991])
);

LUT6 #(
   .INIT(64'h24f848d924f848d9)  
) LUT6_inst8108 (
   .O(to_level3[332]),
   .I0(level4_in[1992]),
   .I1(level4_in[1993]),
   .I2(level4_in[1994]),
   .I3(level4_in[1995]),
   .I4(level4_in[1996]),
   .I5(level4_in[1997])
);

LUT6 #(
   .INIT(64'h8411ae988411ae98)  
) LUT6_inst8109 (
   .O(to_level3[333]),
   .I0(level4_in[1998]),
   .I1(level4_in[1999]),
   .I2(level4_in[2000]),
   .I3(level4_in[2001]),
   .I4(level4_in[2002]),
   .I5(level4_in[2003])
);

LUT6 #(
   .INIT(64'h11c1c7b411c1c7b4)  
) LUT6_inst8110 (
   .O(to_level3[334]),
   .I0(level4_in[2004]),
   .I1(level4_in[2005]),
   .I2(level4_in[2006]),
   .I3(level4_in[2007]),
   .I4(level4_in[2008]),
   .I5(level4_in[2009])
);

LUT6 #(
   .INIT(64'h99b599b699b599b6)  
) LUT6_inst8111 (
   .O(to_level3[335]),
   .I0(level4_in[2010]),
   .I1(level4_in[2011]),
   .I2(level4_in[2012]),
   .I3(level4_in[2013]),
   .I4(level4_in[2014]),
   .I5(level4_in[2015])
);

LUT6 #(
   .INIT(64'h7189678e7189678e)  
) LUT6_inst8112 (
   .O(to_level3[336]),
   .I0(level4_in[2016]),
   .I1(level4_in[2017]),
   .I2(level4_in[2018]),
   .I3(level4_in[2019]),
   .I4(level4_in[2020]),
   .I5(level4_in[2021])
);

LUT6 #(
   .INIT(64'h613f25ef613f25ef)  
) LUT6_inst8113 (
   .O(to_level3[337]),
   .I0(level4_in[2022]),
   .I1(level4_in[2023]),
   .I2(level4_in[2024]),
   .I3(level4_in[2025]),
   .I4(level4_in[2026]),
   .I5(level4_in[2027])
);

LUT6 #(
   .INIT(64'h464ae557464ae557)  
) LUT6_inst8114 (
   .O(to_level3[338]),
   .I0(level4_in[2028]),
   .I1(level4_in[2029]),
   .I2(level4_in[2030]),
   .I3(level4_in[2031]),
   .I4(level4_in[2032]),
   .I5(level4_in[2033])
);

LUT6 #(
   .INIT(64'h6f8c5f6f6f8c5f6f)  
) LUT6_inst8115 (
   .O(to_level3[339]),
   .I0(level4_in[2034]),
   .I1(level4_in[2035]),
   .I2(level4_in[2036]),
   .I3(level4_in[2037]),
   .I4(level4_in[2038]),
   .I5(level4_in[2039])
);

LUT6 #(
   .INIT(64'hb67d7c65b67d7c65)  
) LUT6_inst8116 (
   .O(to_level3[340]),
   .I0(level4_in[2040]),
   .I1(level4_in[2041]),
   .I2(level4_in[2042]),
   .I3(level4_in[2043]),
   .I4(level4_in[2044]),
   .I5(level4_in[2045])
);

LUT6 #(
   .INIT(64'h8e2436948e243694)  
) LUT6_inst8117 (
   .O(to_level3[341]),
   .I0(level4_in[2046]),
   .I1(level4_in[2047]),
   .I2(level4_in[2048]),
   .I3(level4_in[2049]),
   .I4(level4_in[2050]),
   .I5(level4_in[2051])
);

LUT6 #(
   .INIT(64'hd2f1b750d2f1b750)  
) LUT6_inst8118 (
   .O(to_level3[342]),
   .I0(level4_in[2052]),
   .I1(level4_in[2053]),
   .I2(level4_in[2054]),
   .I3(level4_in[2055]),
   .I4(level4_in[2056]),
   .I5(level4_in[2057])
);

LUT6 #(
   .INIT(64'h59f50e5f59f50e5f)  
) LUT6_inst8119 (
   .O(to_level3[343]),
   .I0(level4_in[2058]),
   .I1(level4_in[2059]),
   .I2(level4_in[2060]),
   .I3(level4_in[2061]),
   .I4(level4_in[2062]),
   .I5(level4_in[2063])
);

LUT6 #(
   .INIT(64'hf477411df477411d)  
) LUT6_inst8120 (
   .O(to_level3[344]),
   .I0(level4_in[2064]),
   .I1(level4_in[2065]),
   .I2(level4_in[2066]),
   .I3(level4_in[2067]),
   .I4(level4_in[2068]),
   .I5(level4_in[2069])
);

LUT6 #(
   .INIT(64'h2bcb32c82bcb32c8)  
) LUT6_inst8121 (
   .O(to_level3[345]),
   .I0(level4_in[2070]),
   .I1(level4_in[2071]),
   .I2(level4_in[2072]),
   .I3(level4_in[2073]),
   .I4(level4_in[2074]),
   .I5(level4_in[2075])
);

LUT6 #(
   .INIT(64'hb94c6b56b94c6b56)  
) LUT6_inst8122 (
   .O(to_level3[346]),
   .I0(level4_in[2076]),
   .I1(level4_in[2077]),
   .I2(level4_in[2078]),
   .I3(level4_in[2079]),
   .I4(level4_in[2080]),
   .I5(level4_in[2081])
);

LUT6 #(
   .INIT(64'h3218b6d93218b6d9)  
) LUT6_inst8123 (
   .O(to_level3[347]),
   .I0(level4_in[2082]),
   .I1(level4_in[2083]),
   .I2(level4_in[2084]),
   .I3(level4_in[2085]),
   .I4(level4_in[2086]),
   .I5(level4_in[2087])
);

LUT6 #(
   .INIT(64'h1581492615814926)  
) LUT6_inst8124 (
   .O(to_level3[348]),
   .I0(level4_in[2088]),
   .I1(level4_in[2089]),
   .I2(level4_in[2090]),
   .I3(level4_in[2091]),
   .I4(level4_in[2092]),
   .I5(level4_in[2093])
);

LUT6 #(
   .INIT(64'haf35f72caf35f72c)  
) LUT6_inst8125 (
   .O(to_level3[349]),
   .I0(level4_in[2094]),
   .I1(level4_in[2095]),
   .I2(level4_in[2096]),
   .I3(level4_in[2097]),
   .I4(level4_in[2098]),
   .I5(level4_in[2099])
);

LUT6 #(
   .INIT(64'hc5885b92c5885b92)  
) LUT6_inst8126 (
   .O(to_level3[350]),
   .I0(level4_in[2100]),
   .I1(level4_in[2101]),
   .I2(level4_in[2102]),
   .I3(level4_in[2103]),
   .I4(level4_in[2104]),
   .I5(level4_in[2105])
);

LUT6 #(
   .INIT(64'hccd4f20fccd4f20f)  
) LUT6_inst8127 (
   .O(to_level3[351]),
   .I0(level4_in[2106]),
   .I1(level4_in[2107]),
   .I2(level4_in[2108]),
   .I3(level4_in[2109]),
   .I4(level4_in[2110]),
   .I5(level4_in[2111])
);

LUT6 #(
   .INIT(64'h049d2691049d2691)  
) LUT6_inst8128 (
   .O(to_level3[352]),
   .I0(level4_in[2112]),
   .I1(level4_in[2113]),
   .I2(level4_in[2114]),
   .I3(level4_in[2115]),
   .I4(level4_in[2116]),
   .I5(level4_in[2117])
);

LUT6 #(
   .INIT(64'h269e9e03269e9e03)  
) LUT6_inst8129 (
   .O(to_level3[353]),
   .I0(level4_in[2118]),
   .I1(level4_in[2119]),
   .I2(level4_in[2120]),
   .I3(level4_in[2121]),
   .I4(level4_in[2122]),
   .I5(level4_in[2123])
);

LUT6 #(
   .INIT(64'he55e9f0ae55e9f0a)  
) LUT6_inst8130 (
   .O(to_level3[354]),
   .I0(level4_in[2124]),
   .I1(level4_in[2125]),
   .I2(level4_in[2126]),
   .I3(level4_in[2127]),
   .I4(level4_in[2128]),
   .I5(level4_in[2129])
);

LUT6 #(
   .INIT(64'hab9eaa93ab9eaa93)  
) LUT6_inst8131 (
   .O(to_level3[355]),
   .I0(level4_in[2130]),
   .I1(level4_in[2131]),
   .I2(level4_in[2132]),
   .I3(level4_in[2133]),
   .I4(level4_in[2134]),
   .I5(level4_in[2135])
);

LUT6 #(
   .INIT(64'h71d7052d71d7052d)  
) LUT6_inst8132 (
   .O(to_level3[356]),
   .I0(level4_in[2136]),
   .I1(level4_in[2137]),
   .I2(level4_in[2138]),
   .I3(level4_in[2139]),
   .I4(level4_in[2140]),
   .I5(level4_in[2141])
);

LUT6 #(
   .INIT(64'hbf59cf70bf59cf70)  
) LUT6_inst8133 (
   .O(to_level3[357]),
   .I0(level4_in[2142]),
   .I1(level4_in[2143]),
   .I2(level4_in[2144]),
   .I3(level4_in[2145]),
   .I4(level4_in[2146]),
   .I5(level4_in[2147])
);

LUT6 #(
   .INIT(64'hcb9d6b3acb9d6b3a)  
) LUT6_inst8134 (
   .O(to_level3[358]),
   .I0(level4_in[2148]),
   .I1(level4_in[2149]),
   .I2(level4_in[2150]),
   .I3(level4_in[2151]),
   .I4(level4_in[2152]),
   .I5(level4_in[2153])
);

LUT6 #(
   .INIT(64'h6ac803c96ac803c9)  
) LUT6_inst8135 (
   .O(to_level3[359]),
   .I0(level4_in[2154]),
   .I1(level4_in[2155]),
   .I2(level4_in[2156]),
   .I3(level4_in[2157]),
   .I4(level4_in[2158]),
   .I5(level4_in[2159])
);

LUT6 #(
   .INIT(64'h00a3703d00a3703d)  
) LUT6_inst8136 (
   .O(to_level3[360]),
   .I0(level4_in[2160]),
   .I1(level4_in[2161]),
   .I2(level4_in[2162]),
   .I3(level4_in[2163]),
   .I4(level4_in[2164]),
   .I5(level4_in[2165])
);

LUT6 #(
   .INIT(64'h6ec29d266ec29d26)  
) LUT6_inst8137 (
   .O(to_level3[361]),
   .I0(level4_in[2166]),
   .I1(level4_in[2167]),
   .I2(level4_in[2168]),
   .I3(level4_in[2169]),
   .I4(level4_in[2170]),
   .I5(level4_in[2171])
);

LUT6 #(
   .INIT(64'hee0cae6aee0cae6a)  
) LUT6_inst8138 (
   .O(to_level3[362]),
   .I0(level4_in[2172]),
   .I1(level4_in[2173]),
   .I2(level4_in[2174]),
   .I3(level4_in[2175]),
   .I4(level4_in[2176]),
   .I5(level4_in[2177])
);

LUT6 #(
   .INIT(64'h76f8f0b476f8f0b4)  
) LUT6_inst8139 (
   .O(to_level3[363]),
   .I0(level4_in[2178]),
   .I1(level4_in[2179]),
   .I2(level4_in[2180]),
   .I3(level4_in[2181]),
   .I4(level4_in[2182]),
   .I5(level4_in[2183])
);

LUT6 #(
   .INIT(64'h5c7d6ed35c7d6ed3)  
) LUT6_inst8140 (
   .O(to_level3[364]),
   .I0(level4_in[2184]),
   .I1(level4_in[2185]),
   .I2(level4_in[2186]),
   .I3(level4_in[2187]),
   .I4(level4_in[2188]),
   .I5(level4_in[2189])
);

LUT6 #(
   .INIT(64'h2bcd566a2bcd566a)  
) LUT6_inst8141 (
   .O(to_level3[365]),
   .I0(level4_in[2190]),
   .I1(level4_in[2191]),
   .I2(level4_in[2192]),
   .I3(level4_in[2193]),
   .I4(level4_in[2194]),
   .I5(level4_in[2195])
);

LUT6 #(
   .INIT(64'he9dc5655e9dc5655)  
) LUT6_inst8142 (
   .O(to_level3[366]),
   .I0(level4_in[2196]),
   .I1(level4_in[2197]),
   .I2(level4_in[2198]),
   .I3(level4_in[2199]),
   .I4(level4_in[2200]),
   .I5(level4_in[2201])
);

LUT6 #(
   .INIT(64'h32d07c0932d07c09)  
) LUT6_inst8143 (
   .O(to_level3[367]),
   .I0(level4_in[2202]),
   .I1(level4_in[2203]),
   .I2(level4_in[2204]),
   .I3(level4_in[2205]),
   .I4(level4_in[2206]),
   .I5(level4_in[2207])
);

LUT6 #(
   .INIT(64'hc3f931a0c3f931a0)  
) LUT6_inst8144 (
   .O(to_level3[368]),
   .I0(level4_in[2208]),
   .I1(level4_in[2209]),
   .I2(level4_in[2210]),
   .I3(level4_in[2211]),
   .I4(level4_in[2212]),
   .I5(level4_in[2213])
);

LUT6 #(
   .INIT(64'hb4f7e830b4f7e830)  
) LUT6_inst8145 (
   .O(to_level3[369]),
   .I0(level4_in[2214]),
   .I1(level4_in[2215]),
   .I2(level4_in[2216]),
   .I3(level4_in[2217]),
   .I4(level4_in[2218]),
   .I5(level4_in[2219])
);

LUT6 #(
   .INIT(64'h1e271aa41e271aa4)  
) LUT6_inst8146 (
   .O(to_level3[370]),
   .I0(level4_in[2220]),
   .I1(level4_in[2221]),
   .I2(level4_in[2222]),
   .I3(level4_in[2223]),
   .I4(level4_in[2224]),
   .I5(level4_in[2225])
);

LUT6 #(
   .INIT(64'hf65923fcf65923fc)  
) LUT6_inst8147 (
   .O(to_level3[371]),
   .I0(level4_in[2226]),
   .I1(level4_in[2227]),
   .I2(level4_in[2228]),
   .I3(level4_in[2229]),
   .I4(level4_in[2230]),
   .I5(level4_in[2231])
);

LUT6 #(
   .INIT(64'hc5f5a828c5f5a828)  
) LUT6_inst8148 (
   .O(to_level3[372]),
   .I0(level4_in[2232]),
   .I1(level4_in[2233]),
   .I2(level4_in[2234]),
   .I3(level4_in[2235]),
   .I4(level4_in[2236]),
   .I5(level4_in[2237])
);

LUT6 #(
   .INIT(64'hc976994cc976994c)  
) LUT6_inst8149 (
   .O(to_level3[373]),
   .I0(level4_in[2238]),
   .I1(level4_in[2239]),
   .I2(level4_in[2240]),
   .I3(level4_in[2241]),
   .I4(level4_in[2242]),
   .I5(level4_in[2243])
);

LUT6 #(
   .INIT(64'hd07de374d07de374)  
) LUT6_inst8150 (
   .O(to_level3[374]),
   .I0(level4_in[2244]),
   .I1(level4_in[2245]),
   .I2(level4_in[2246]),
   .I3(level4_in[2247]),
   .I4(level4_in[2248]),
   .I5(level4_in[2249])
);

LUT6 #(
   .INIT(64'hce75ec92ce75ec92)  
) LUT6_inst8151 (
   .O(to_level3[375]),
   .I0(level4_in[2250]),
   .I1(level4_in[2251]),
   .I2(level4_in[2252]),
   .I3(level4_in[2253]),
   .I4(level4_in[2254]),
   .I5(level4_in[2255])
);

LUT6 #(
   .INIT(64'h8c67d04d8c67d04d)  
) LUT6_inst8152 (
   .O(to_level3[376]),
   .I0(level4_in[2256]),
   .I1(level4_in[2257]),
   .I2(level4_in[2258]),
   .I3(level4_in[2259]),
   .I4(level4_in[2260]),
   .I5(level4_in[2261])
);

LUT6 #(
   .INIT(64'h1248f1d51248f1d5)  
) LUT6_inst8153 (
   .O(to_level3[377]),
   .I0(level4_in[2262]),
   .I1(level4_in[2263]),
   .I2(level4_in[2264]),
   .I3(level4_in[2265]),
   .I4(level4_in[2266]),
   .I5(level4_in[2267])
);

LUT6 #(
   .INIT(64'h684920bf684920bf)  
) LUT6_inst8154 (
   .O(to_level3[378]),
   .I0(level4_in[2268]),
   .I1(level4_in[2269]),
   .I2(level4_in[2270]),
   .I3(level4_in[2271]),
   .I4(level4_in[2272]),
   .I5(level4_in[2273])
);

LUT6 #(
   .INIT(64'hc98d1a81c98d1a81)  
) LUT6_inst8155 (
   .O(to_level3[379]),
   .I0(level4_in[2274]),
   .I1(level4_in[2275]),
   .I2(level4_in[2276]),
   .I3(level4_in[2277]),
   .I4(level4_in[2278]),
   .I5(level4_in[2279])
);

LUT6 #(
   .INIT(64'h517d72a4517d72a4)  
) LUT6_inst8156 (
   .O(to_level3[380]),
   .I0(level4_in[2280]),
   .I1(level4_in[2281]),
   .I2(level4_in[2282]),
   .I3(level4_in[2283]),
   .I4(level4_in[2284]),
   .I5(level4_in[2285])
);

LUT6 #(
   .INIT(64'h07c210d007c210d0)  
) LUT6_inst8157 (
   .O(to_level3[381]),
   .I0(level4_in[2286]),
   .I1(level4_in[2287]),
   .I2(level4_in[2288]),
   .I3(level4_in[2289]),
   .I4(level4_in[2290]),
   .I5(level4_in[2291])
);

LUT6 #(
   .INIT(64'hd54e81c2d54e81c2)  
) LUT6_inst8158 (
   .O(to_level3[382]),
   .I0(level4_in[2292]),
   .I1(level4_in[2293]),
   .I2(level4_in[2294]),
   .I3(level4_in[2295]),
   .I4(level4_in[2296]),
   .I5(level4_in[2297])
);

LUT6 #(
   .INIT(64'h0cc46cf00cc46cf0)  
) LUT6_inst8159 (
   .O(to_level3[383]),
   .I0(level4_in[2298]),
   .I1(level4_in[2299]),
   .I2(level4_in[2300]),
   .I3(level4_in[2301]),
   .I4(level4_in[2302]),
   .I5(level4_in[2303])
);

LUT6 #(
   .INIT(64'h245e51b1245e51b1)  
) LUT6_inst8160 (
   .O(to_level3[384]),
   .I0(level4_in[2304]),
   .I1(level4_in[2305]),
   .I2(level4_in[2306]),
   .I3(level4_in[2307]),
   .I4(level4_in[2308]),
   .I5(level4_in[2309])
);

LUT6 #(
   .INIT(64'h296463f3296463f3)  
) LUT6_inst8161 (
   .O(to_level3[385]),
   .I0(level4_in[2310]),
   .I1(level4_in[2311]),
   .I2(level4_in[2312]),
   .I3(level4_in[2313]),
   .I4(level4_in[2314]),
   .I5(level4_in[2315])
);

LUT6 #(
   .INIT(64'h485642f9485642f9)  
) LUT6_inst8162 (
   .O(to_level3[386]),
   .I0(level4_in[2316]),
   .I1(level4_in[2317]),
   .I2(level4_in[2318]),
   .I3(level4_in[2319]),
   .I4(level4_in[2320]),
   .I5(level4_in[2321])
);

LUT6 #(
   .INIT(64'h50d62ff550d62ff5)  
) LUT6_inst8163 (
   .O(to_level3[387]),
   .I0(level4_in[2322]),
   .I1(level4_in[2323]),
   .I2(level4_in[2324]),
   .I3(level4_in[2325]),
   .I4(level4_in[2326]),
   .I5(level4_in[2327])
);

LUT6 #(
   .INIT(64'h1b7900591b790059)  
) LUT6_inst8164 (
   .O(to_level3[388]),
   .I0(level4_in[2328]),
   .I1(level4_in[2329]),
   .I2(level4_in[2330]),
   .I3(level4_in[2331]),
   .I4(level4_in[2332]),
   .I5(level4_in[2333])
);

LUT6 #(
   .INIT(64'hcbb5d767cbb5d767)  
) LUT6_inst8165 (
   .O(to_level3[389]),
   .I0(level4_in[2334]),
   .I1(level4_in[2335]),
   .I2(level4_in[2336]),
   .I3(level4_in[2337]),
   .I4(level4_in[2338]),
   .I5(level4_in[2339])
);

LUT6 #(
   .INIT(64'h9764f9e29764f9e2)  
) LUT6_inst8166 (
   .O(to_level3[390]),
   .I0(level4_in[2340]),
   .I1(level4_in[2341]),
   .I2(level4_in[2342]),
   .I3(level4_in[2343]),
   .I4(level4_in[2344]),
   .I5(level4_in[2345])
);

LUT6 #(
   .INIT(64'h7445cc187445cc18)  
) LUT6_inst8167 (
   .O(to_level3[391]),
   .I0(level4_in[2346]),
   .I1(level4_in[2347]),
   .I2(level4_in[2348]),
   .I3(level4_in[2349]),
   .I4(level4_in[2350]),
   .I5(level4_in[2351])
);

LUT6 #(
   .INIT(64'hfe753c31fe753c31)  
) LUT6_inst8168 (
   .O(to_level3[392]),
   .I0(level4_in[2352]),
   .I1(level4_in[2353]),
   .I2(level4_in[2354]),
   .I3(level4_in[2355]),
   .I4(level4_in[2356]),
   .I5(level4_in[2357])
);

LUT6 #(
   .INIT(64'h1566923115669231)  
) LUT6_inst8169 (
   .O(to_level3[393]),
   .I0(level4_in[2358]),
   .I1(level4_in[2359]),
   .I2(level4_in[2360]),
   .I3(level4_in[2361]),
   .I4(level4_in[2362]),
   .I5(level4_in[2363])
);

LUT6 #(
   .INIT(64'hafb6ac3aafb6ac3a)  
) LUT6_inst8170 (
   .O(to_level3[394]),
   .I0(level4_in[2364]),
   .I1(level4_in[2365]),
   .I2(level4_in[2366]),
   .I3(level4_in[2367]),
   .I4(level4_in[2368]),
   .I5(level4_in[2369])
);

LUT6 #(
   .INIT(64'h3aff489f3aff489f)  
) LUT6_inst8171 (
   .O(to_level3[395]),
   .I0(level4_in[2370]),
   .I1(level4_in[2371]),
   .I2(level4_in[2372]),
   .I3(level4_in[2373]),
   .I4(level4_in[2374]),
   .I5(level4_in[2375])
);

LUT6 #(
   .INIT(64'h9914209f9914209f)  
) LUT6_inst8172 (
   .O(to_level3[396]),
   .I0(level4_in[2376]),
   .I1(level4_in[2377]),
   .I2(level4_in[2378]),
   .I3(level4_in[2379]),
   .I4(level4_in[2380]),
   .I5(level4_in[2381])
);

LUT6 #(
   .INIT(64'h528d66da528d66da)  
) LUT6_inst8173 (
   .O(to_level3[397]),
   .I0(level4_in[2382]),
   .I1(level4_in[2383]),
   .I2(level4_in[2384]),
   .I3(level4_in[2385]),
   .I4(level4_in[2386]),
   .I5(level4_in[2387])
);

LUT6 #(
   .INIT(64'h4f9faaef4f9faaef)  
) LUT6_inst8174 (
   .O(to_level3[398]),
   .I0(level4_in[2388]),
   .I1(level4_in[2389]),
   .I2(level4_in[2390]),
   .I3(level4_in[2391]),
   .I4(level4_in[2392]),
   .I5(level4_in[2393])
);

LUT6 #(
   .INIT(64'h27e8155327e81553)  
) LUT6_inst8175 (
   .O(to_level3[399]),
   .I0(level4_in[2394]),
   .I1(level4_in[2395]),
   .I2(level4_in[2396]),
   .I3(level4_in[2397]),
   .I4(level4_in[2398]),
   .I5(level4_in[2399])
);

LUT6 #(
   .INIT(64'hb03d628ab03d628a)  
) LUT6_inst8176 (
   .O(to_level3[400]),
   .I0(level4_in[2400]),
   .I1(level4_in[2401]),
   .I2(level4_in[2402]),
   .I3(level4_in[2403]),
   .I4(level4_in[2404]),
   .I5(level4_in[2405])
);

LUT6 #(
   .INIT(64'h860e569b860e569b)  
) LUT6_inst8177 (
   .O(to_level3[401]),
   .I0(level4_in[2406]),
   .I1(level4_in[2407]),
   .I2(level4_in[2408]),
   .I3(level4_in[2409]),
   .I4(level4_in[2410]),
   .I5(level4_in[2411])
);

LUT6 #(
   .INIT(64'h0a7cd1d00a7cd1d0)  
) LUT6_inst8178 (
   .O(to_level3[402]),
   .I0(level4_in[2412]),
   .I1(level4_in[2413]),
   .I2(level4_in[2414]),
   .I3(level4_in[2415]),
   .I4(level4_in[2416]),
   .I5(level4_in[2417])
);

LUT6 #(
   .INIT(64'hc83de1fec83de1fe)  
) LUT6_inst8179 (
   .O(to_level3[403]),
   .I0(level4_in[2418]),
   .I1(level4_in[2419]),
   .I2(level4_in[2420]),
   .I3(level4_in[2421]),
   .I4(level4_in[2422]),
   .I5(level4_in[2423])
);

LUT6 #(
   .INIT(64'hf9f3f787f9f3f787)  
) LUT6_inst8180 (
   .O(to_level3[404]),
   .I0(level4_in[2424]),
   .I1(level4_in[2425]),
   .I2(level4_in[2426]),
   .I3(level4_in[2427]),
   .I4(level4_in[2428]),
   .I5(level4_in[2429])
);

LUT6 #(
   .INIT(64'ha32fdc5ca32fdc5c)  
) LUT6_inst8181 (
   .O(to_level3[405]),
   .I0(level4_in[2430]),
   .I1(level4_in[2431]),
   .I2(level4_in[2432]),
   .I3(level4_in[2433]),
   .I4(level4_in[2434]),
   .I5(level4_in[2435])
);

LUT6 #(
   .INIT(64'h89f36a7b89f36a7b)  
) LUT6_inst8182 (
   .O(to_level3[406]),
   .I0(level4_in[2436]),
   .I1(level4_in[2437]),
   .I2(level4_in[2438]),
   .I3(level4_in[2439]),
   .I4(level4_in[2440]),
   .I5(level4_in[2441])
);

LUT6 #(
   .INIT(64'h8d3306b78d3306b7)  
) LUT6_inst8183 (
   .O(to_level3[407]),
   .I0(level4_in[2442]),
   .I1(level4_in[2443]),
   .I2(level4_in[2444]),
   .I3(level4_in[2445]),
   .I4(level4_in[2446]),
   .I5(level4_in[2447])
);

LUT6 #(
   .INIT(64'hde7e5ee0de7e5ee0)  
) LUT6_inst8184 (
   .O(to_level3[408]),
   .I0(level4_in[2448]),
   .I1(level4_in[2449]),
   .I2(level4_in[2450]),
   .I3(level4_in[2451]),
   .I4(level4_in[2452]),
   .I5(level4_in[2453])
);

LUT6 #(
   .INIT(64'h8655d2a78655d2a7)  
) LUT6_inst8185 (
   .O(to_level3[409]),
   .I0(level4_in[2454]),
   .I1(level4_in[2455]),
   .I2(level4_in[2456]),
   .I3(level4_in[2457]),
   .I4(level4_in[2458]),
   .I5(level4_in[2459])
);

LUT6 #(
   .INIT(64'h4af2fdc14af2fdc1)  
) LUT6_inst8186 (
   .O(to_level3[410]),
   .I0(level4_in[2460]),
   .I1(level4_in[2461]),
   .I2(level4_in[2462]),
   .I3(level4_in[2463]),
   .I4(level4_in[2464]),
   .I5(level4_in[2465])
);

LUT6 #(
   .INIT(64'hb859fd59b859fd59)  
) LUT6_inst8187 (
   .O(to_level3[411]),
   .I0(level4_in[2466]),
   .I1(level4_in[2467]),
   .I2(level4_in[2468]),
   .I3(level4_in[2469]),
   .I4(level4_in[2470]),
   .I5(level4_in[2471])
);

LUT6 #(
   .INIT(64'hbe12438abe12438a)  
) LUT6_inst8188 (
   .O(to_level3[412]),
   .I0(level4_in[2472]),
   .I1(level4_in[2473]),
   .I2(level4_in[2474]),
   .I3(level4_in[2475]),
   .I4(level4_in[2476]),
   .I5(level4_in[2477])
);

LUT6 #(
   .INIT(64'h0c089eb60c089eb6)  
) LUT6_inst8189 (
   .O(to_level3[413]),
   .I0(level4_in[2478]),
   .I1(level4_in[2479]),
   .I2(level4_in[2480]),
   .I3(level4_in[2481]),
   .I4(level4_in[2482]),
   .I5(level4_in[2483])
);

LUT6 #(
   .INIT(64'h9e508a919e508a91)  
) LUT6_inst8190 (
   .O(to_level3[414]),
   .I0(level4_in[2484]),
   .I1(level4_in[2485]),
   .I2(level4_in[2486]),
   .I3(level4_in[2487]),
   .I4(level4_in[2488]),
   .I5(level4_in[2489])
);

LUT6 #(
   .INIT(64'ha446b98fa446b98f)  
) LUT6_inst8191 (
   .O(to_level3[415]),
   .I0(level4_in[2490]),
   .I1(level4_in[2491]),
   .I2(level4_in[2492]),
   .I3(level4_in[2493]),
   .I4(level4_in[2494]),
   .I5(level4_in[2495])
);

LUT6 #(
   .INIT(64'h0e68000f0e68000f)  
) LUT6_inst8192 (
   .O(to_level3[416]),
   .I0(level4_in[2496]),
   .I1(level4_in[2497]),
   .I2(level4_in[2498]),
   .I3(level4_in[2499]),
   .I4(level4_in[2500]),
   .I5(level4_in[2501])
);

LUT6 #(
   .INIT(64'hd80de174d80de174)  
) LUT6_inst8193 (
   .O(to_level3[417]),
   .I0(level4_in[2502]),
   .I1(level4_in[2503]),
   .I2(level4_in[2504]),
   .I3(level4_in[2505]),
   .I4(level4_in[2506]),
   .I5(level4_in[2507])
);

LUT6 #(
   .INIT(64'hdb3b834cdb3b834c)  
) LUT6_inst8194 (
   .O(to_level3[418]),
   .I0(level4_in[2508]),
   .I1(level4_in[2509]),
   .I2(level4_in[2510]),
   .I3(level4_in[2511]),
   .I4(level4_in[2512]),
   .I5(level4_in[2513])
);

LUT6 #(
   .INIT(64'h5ea8cb625ea8cb62)  
) LUT6_inst8195 (
   .O(to_level3[419]),
   .I0(level4_in[2514]),
   .I1(level4_in[2515]),
   .I2(level4_in[2516]),
   .I3(level4_in[2517]),
   .I4(level4_in[2518]),
   .I5(level4_in[2519])
);

LUT6 #(
   .INIT(64'he6154aa8e6154aa8)  
) LUT6_inst8196 (
   .O(to_level3[420]),
   .I0(level4_in[2520]),
   .I1(level4_in[2521]),
   .I2(level4_in[2522]),
   .I3(level4_in[2523]),
   .I4(level4_in[2524]),
   .I5(level4_in[2525])
);

LUT6 #(
   .INIT(64'h720ddb5a720ddb5a)  
) LUT6_inst8197 (
   .O(to_level3[421]),
   .I0(level4_in[2526]),
   .I1(level4_in[2527]),
   .I2(level4_in[2528]),
   .I3(level4_in[2529]),
   .I4(level4_in[2530]),
   .I5(level4_in[2531])
);

LUT6 #(
   .INIT(64'h2cdbe1f32cdbe1f3)  
) LUT6_inst8198 (
   .O(to_level3[422]),
   .I0(level4_in[2532]),
   .I1(level4_in[2533]),
   .I2(level4_in[2534]),
   .I3(level4_in[2535]),
   .I4(level4_in[2536]),
   .I5(level4_in[2537])
);

LUT6 #(
   .INIT(64'hf687decef687dece)  
) LUT6_inst8199 (
   .O(to_level3[423]),
   .I0(level4_in[2538]),
   .I1(level4_in[2539]),
   .I2(level4_in[2540]),
   .I3(level4_in[2541]),
   .I4(level4_in[2542]),
   .I5(level4_in[2543])
);

LUT6 #(
   .INIT(64'h93f3f23d93f3f23d)  
) LUT6_inst8200 (
   .O(to_level3[424]),
   .I0(level4_in[2544]),
   .I1(level4_in[2545]),
   .I2(level4_in[2546]),
   .I3(level4_in[2547]),
   .I4(level4_in[2548]),
   .I5(level4_in[2549])
);

LUT6 #(
   .INIT(64'h762ed596762ed596)  
) LUT6_inst8201 (
   .O(to_level3[425]),
   .I0(level4_in[2550]),
   .I1(level4_in[2551]),
   .I2(level4_in[2552]),
   .I3(level4_in[2553]),
   .I4(level4_in[2554]),
   .I5(level4_in[2555])
);

LUT6 #(
   .INIT(64'ha0a0ce48a0a0ce48)  
) LUT6_inst8202 (
   .O(to_level3[426]),
   .I0(level4_in[2556]),
   .I1(level4_in[2557]),
   .I2(level4_in[2558]),
   .I3(level4_in[2559]),
   .I4(level4_in[2560]),
   .I5(level4_in[2561])
);

LUT6 #(
   .INIT(64'h54e44d3e54e44d3e)  
) LUT6_inst8203 (
   .O(to_level3[427]),
   .I0(level4_in[2562]),
   .I1(level4_in[2563]),
   .I2(level4_in[2564]),
   .I3(level4_in[2565]),
   .I4(level4_in[2566]),
   .I5(level4_in[2567])
);

LUT6 #(
   .INIT(64'h2608a8592608a859)  
) LUT6_inst8204 (
   .O(to_level3[428]),
   .I0(level4_in[2568]),
   .I1(level4_in[2569]),
   .I2(level4_in[2570]),
   .I3(level4_in[2571]),
   .I4(level4_in[2572]),
   .I5(level4_in[2573])
);

LUT6 #(
   .INIT(64'h338cf9f2338cf9f2)  
) LUT6_inst8205 (
   .O(to_level3[429]),
   .I0(level4_in[2574]),
   .I1(level4_in[2575]),
   .I2(level4_in[2576]),
   .I3(level4_in[2577]),
   .I4(level4_in[2578]),
   .I5(level4_in[2579])
);

LUT6 #(
   .INIT(64'h6b32dead6b32dead)  
) LUT6_inst8206 (
   .O(to_level3[430]),
   .I0(level4_in[2580]),
   .I1(level4_in[2581]),
   .I2(level4_in[2582]),
   .I3(level4_in[2583]),
   .I4(level4_in[2584]),
   .I5(level4_in[2585])
);

LUT6 #(
   .INIT(64'h72079de072079de0)  
) LUT6_inst8207 (
   .O(to_level3[431]),
   .I0(level4_in[2586]),
   .I1(level4_in[2587]),
   .I2(level4_in[2588]),
   .I3(level4_in[2589]),
   .I4(level4_in[2590]),
   .I5(level4_in[2591])
);

LUT6 #(
   .INIT(64'h7560163675601636)  
) LUT6_inst8208 (
   .O(to_level3[432]),
   .I0(level4_in[2592]),
   .I1(level4_in[2593]),
   .I2(level4_in[2594]),
   .I3(level4_in[2595]),
   .I4(level4_in[2596]),
   .I5(level4_in[2597])
);

LUT6 #(
   .INIT(64'h007b790b007b790b)  
) LUT6_inst8209 (
   .O(to_level3[433]),
   .I0(level4_in[2598]),
   .I1(level4_in[2599]),
   .I2(level4_in[2600]),
   .I3(level4_in[2601]),
   .I4(level4_in[2602]),
   .I5(level4_in[2603])
);

LUT6 #(
   .INIT(64'h3434321434343214)  
) LUT6_inst8210 (
   .O(to_level3[434]),
   .I0(level4_in[2604]),
   .I1(level4_in[2605]),
   .I2(level4_in[2606]),
   .I3(level4_in[2607]),
   .I4(level4_in[2608]),
   .I5(level4_in[2609])
);

LUT6 #(
   .INIT(64'h0f50e18f0f50e18f)  
) LUT6_inst8211 (
   .O(to_level3[435]),
   .I0(level4_in[2610]),
   .I1(level4_in[2611]),
   .I2(level4_in[2612]),
   .I3(level4_in[2613]),
   .I4(level4_in[2614]),
   .I5(level4_in[2615])
);

LUT6 #(
   .INIT(64'h6a70939f6a70939f)  
) LUT6_inst8212 (
   .O(to_level3[436]),
   .I0(level4_in[2616]),
   .I1(level4_in[2617]),
   .I2(level4_in[2618]),
   .I3(level4_in[2619]),
   .I4(level4_in[2620]),
   .I5(level4_in[2621])
);

LUT6 #(
   .INIT(64'h366917ee366917ee)  
) LUT6_inst8213 (
   .O(to_level3[437]),
   .I0(level4_in[2622]),
   .I1(level4_in[2623]),
   .I2(level4_in[2624]),
   .I3(level4_in[2625]),
   .I4(level4_in[2626]),
   .I5(level4_in[2627])
);

LUT6 #(
   .INIT(64'hf89d4941f89d4941)  
) LUT6_inst8214 (
   .O(to_level3[438]),
   .I0(level4_in[2628]),
   .I1(level4_in[2629]),
   .I2(level4_in[2630]),
   .I3(level4_in[2631]),
   .I4(level4_in[2632]),
   .I5(level4_in[2633])
);

LUT6 #(
   .INIT(64'hb04b97b9b04b97b9)  
) LUT6_inst8215 (
   .O(to_level3[439]),
   .I0(level4_in[2634]),
   .I1(level4_in[2635]),
   .I2(level4_in[2636]),
   .I3(level4_in[2637]),
   .I4(level4_in[2638]),
   .I5(level4_in[2639])
);

LUT6 #(
   .INIT(64'hd5a6d42fd5a6d42f)  
) LUT6_inst8216 (
   .O(to_level3[440]),
   .I0(level4_in[2640]),
   .I1(level4_in[2641]),
   .I2(level4_in[2642]),
   .I3(level4_in[2643]),
   .I4(level4_in[2644]),
   .I5(level4_in[2645])
);

LUT6 #(
   .INIT(64'hc20b0f59c20b0f59)  
) LUT6_inst8217 (
   .O(to_level3[441]),
   .I0(level4_in[2646]),
   .I1(level4_in[2647]),
   .I2(level4_in[2648]),
   .I3(level4_in[2649]),
   .I4(level4_in[2650]),
   .I5(level4_in[2651])
);

LUT6 #(
   .INIT(64'h6960eb966960eb96)  
) LUT6_inst8218 (
   .O(to_level3[442]),
   .I0(level4_in[2652]),
   .I1(level4_in[2653]),
   .I2(level4_in[2654]),
   .I3(level4_in[2655]),
   .I4(level4_in[2656]),
   .I5(level4_in[2657])
);

LUT6 #(
   .INIT(64'h2bb88a8b2bb88a8b)  
) LUT6_inst8219 (
   .O(to_level3[443]),
   .I0(level4_in[2658]),
   .I1(level4_in[2659]),
   .I2(level4_in[2660]),
   .I3(level4_in[2661]),
   .I4(level4_in[2662]),
   .I5(level4_in[2663])
);

LUT6 #(
   .INIT(64'h6888e8e26888e8e2)  
) LUT6_inst8220 (
   .O(to_level3[444]),
   .I0(level4_in[2664]),
   .I1(level4_in[2665]),
   .I2(level4_in[2666]),
   .I3(level4_in[2667]),
   .I4(level4_in[2668]),
   .I5(level4_in[2669])
);

LUT6 #(
   .INIT(64'hc811bbe9c811bbe9)  
) LUT6_inst8221 (
   .O(to_level3[445]),
   .I0(level4_in[2670]),
   .I1(level4_in[2671]),
   .I2(level4_in[2672]),
   .I3(level4_in[2673]),
   .I4(level4_in[2674]),
   .I5(level4_in[2675])
);

LUT6 #(
   .INIT(64'h2bc870092bc87009)  
) LUT6_inst8222 (
   .O(to_level3[446]),
   .I0(level4_in[2676]),
   .I1(level4_in[2677]),
   .I2(level4_in[2678]),
   .I3(level4_in[2679]),
   .I4(level4_in[2680]),
   .I5(level4_in[2681])
);

LUT6 #(
   .INIT(64'hbf53f3c4bf53f3c4)  
) LUT6_inst8223 (
   .O(to_level3[447]),
   .I0(level4_in[2682]),
   .I1(level4_in[2683]),
   .I2(level4_in[2684]),
   .I3(level4_in[2685]),
   .I4(level4_in[2686]),
   .I5(level4_in[2687])
);

LUT6 #(
   .INIT(64'h9bf54ed49bf54ed4)  
) LUT6_inst8224 (
   .O(to_level3[448]),
   .I0(level4_in[2688]),
   .I1(level4_in[2689]),
   .I2(level4_in[2690]),
   .I3(level4_in[2691]),
   .I4(level4_in[2692]),
   .I5(level4_in[2693])
);

LUT6 #(
   .INIT(64'h3e9131ae3e9131ae)  
) LUT6_inst8225 (
   .O(to_level3[449]),
   .I0(level4_in[2694]),
   .I1(level4_in[2695]),
   .I2(level4_in[2696]),
   .I3(level4_in[2697]),
   .I4(level4_in[2698]),
   .I5(level4_in[2699])
);

LUT6 #(
   .INIT(64'haa288c3daa288c3d)  
) LUT6_inst8226 (
   .O(to_level3[450]),
   .I0(level4_in[2700]),
   .I1(level4_in[2701]),
   .I2(level4_in[2702]),
   .I3(level4_in[2703]),
   .I4(level4_in[2704]),
   .I5(level4_in[2705])
);

LUT6 #(
   .INIT(64'hed4f96e3ed4f96e3)  
) LUT6_inst8227 (
   .O(to_level3[451]),
   .I0(level4_in[2706]),
   .I1(level4_in[2707]),
   .I2(level4_in[2708]),
   .I3(level4_in[2709]),
   .I4(level4_in[2710]),
   .I5(level4_in[2711])
);

LUT6 #(
   .INIT(64'h0cc5de430cc5de43)  
) LUT6_inst8228 (
   .O(to_level3[452]),
   .I0(level4_in[2712]),
   .I1(level4_in[2713]),
   .I2(level4_in[2714]),
   .I3(level4_in[2715]),
   .I4(level4_in[2716]),
   .I5(level4_in[2717])
);

LUT6 #(
   .INIT(64'hef7be455ef7be455)  
) LUT6_inst8229 (
   .O(to_level3[453]),
   .I0(level4_in[2718]),
   .I1(level4_in[2719]),
   .I2(level4_in[2720]),
   .I3(level4_in[2721]),
   .I4(level4_in[2722]),
   .I5(level4_in[2723])
);

LUT6 #(
   .INIT(64'h83fa4d6883fa4d68)  
) LUT6_inst8230 (
   .O(to_level3[454]),
   .I0(level4_in[2724]),
   .I1(level4_in[2725]),
   .I2(level4_in[2726]),
   .I3(level4_in[2727]),
   .I4(level4_in[2728]),
   .I5(level4_in[2729])
);

LUT6 #(
   .INIT(64'hf9b763f6f9b763f6)  
) LUT6_inst8231 (
   .O(to_level3[455]),
   .I0(level4_in[2730]),
   .I1(level4_in[2731]),
   .I2(level4_in[2732]),
   .I3(level4_in[2733]),
   .I4(level4_in[2734]),
   .I5(level4_in[2735])
);

LUT6 #(
   .INIT(64'h1a27ce7b1a27ce7b)  
) LUT6_inst8232 (
   .O(to_level3[456]),
   .I0(level4_in[2736]),
   .I1(level4_in[2737]),
   .I2(level4_in[2738]),
   .I3(level4_in[2739]),
   .I4(level4_in[2740]),
   .I5(level4_in[2741])
);

LUT6 #(
   .INIT(64'h8c26726f8c26726f)  
) LUT6_inst8233 (
   .O(to_level3[457]),
   .I0(level4_in[2742]),
   .I1(level4_in[2743]),
   .I2(level4_in[2744]),
   .I3(level4_in[2745]),
   .I4(level4_in[2746]),
   .I5(level4_in[2747])
);

LUT6 #(
   .INIT(64'hfbe42fbffbe42fbf)  
) LUT6_inst8234 (
   .O(to_level3[458]),
   .I0(level4_in[2748]),
   .I1(level4_in[2749]),
   .I2(level4_in[2750]),
   .I3(level4_in[2751]),
   .I4(level4_in[2752]),
   .I5(level4_in[2753])
);

LUT6 #(
   .INIT(64'h0ee0f9cd0ee0f9cd)  
) LUT6_inst8235 (
   .O(to_level3[459]),
   .I0(level4_in[2754]),
   .I1(level4_in[2755]),
   .I2(level4_in[2756]),
   .I3(level4_in[2757]),
   .I4(level4_in[2758]),
   .I5(level4_in[2759])
);

LUT6 #(
   .INIT(64'hfb53f02afb53f02a)  
) LUT6_inst8236 (
   .O(to_level3[460]),
   .I0(level4_in[2760]),
   .I1(level4_in[2761]),
   .I2(level4_in[2762]),
   .I3(level4_in[2763]),
   .I4(level4_in[2764]),
   .I5(level4_in[2765])
);

LUT6 #(
   .INIT(64'hd9e227fbd9e227fb)  
) LUT6_inst8237 (
   .O(to_level3[461]),
   .I0(level4_in[2766]),
   .I1(level4_in[2767]),
   .I2(level4_in[2768]),
   .I3(level4_in[2769]),
   .I4(level4_in[2770]),
   .I5(level4_in[2771])
);

LUT6 #(
   .INIT(64'h57c21c9957c21c99)  
) LUT6_inst8238 (
   .O(to_level3[462]),
   .I0(level4_in[2772]),
   .I1(level4_in[2773]),
   .I2(level4_in[2774]),
   .I3(level4_in[2775]),
   .I4(level4_in[2776]),
   .I5(level4_in[2777])
);

LUT6 #(
   .INIT(64'h5c561fa95c561fa9)  
) LUT6_inst8239 (
   .O(to_level3[463]),
   .I0(level4_in[2778]),
   .I1(level4_in[2779]),
   .I2(level4_in[2780]),
   .I3(level4_in[2781]),
   .I4(level4_in[2782]),
   .I5(level4_in[2783])
);

LUT6 #(
   .INIT(64'h09aa64df09aa64df)  
) LUT6_inst8240 (
   .O(to_level3[464]),
   .I0(level4_in[2784]),
   .I1(level4_in[2785]),
   .I2(level4_in[2786]),
   .I3(level4_in[2787]),
   .I4(level4_in[2788]),
   .I5(level4_in[2789])
);

LUT6 #(
   .INIT(64'h5f698cb95f698cb9)  
) LUT6_inst8241 (
   .O(to_level3[465]),
   .I0(level4_in[2790]),
   .I1(level4_in[2791]),
   .I2(level4_in[2792]),
   .I3(level4_in[2793]),
   .I4(level4_in[2794]),
   .I5(level4_in[2795])
);

LUT6 #(
   .INIT(64'hc698597cc698597c)  
) LUT6_inst8242 (
   .O(to_level3[466]),
   .I0(level4_in[2796]),
   .I1(level4_in[2797]),
   .I2(level4_in[2798]),
   .I3(level4_in[2799]),
   .I4(level4_in[2800]),
   .I5(level4_in[2801])
);

LUT6 #(
   .INIT(64'he5be1ecae5be1eca)  
) LUT6_inst8243 (
   .O(to_level3[467]),
   .I0(level4_in[2802]),
   .I1(level4_in[2803]),
   .I2(level4_in[2804]),
   .I3(level4_in[2805]),
   .I4(level4_in[2806]),
   .I5(level4_in[2807])
);

LUT6 #(
   .INIT(64'h43a6a68843a6a688)  
) LUT6_inst8244 (
   .O(to_level3[468]),
   .I0(level4_in[2808]),
   .I1(level4_in[2809]),
   .I2(level4_in[2810]),
   .I3(level4_in[2811]),
   .I4(level4_in[2812]),
   .I5(level4_in[2813])
);

LUT6 #(
   .INIT(64'h8b5d841c8b5d841c)  
) LUT6_inst8245 (
   .O(to_level3[469]),
   .I0(level4_in[2814]),
   .I1(level4_in[2815]),
   .I2(level4_in[2816]),
   .I3(level4_in[2817]),
   .I4(level4_in[2818]),
   .I5(level4_in[2819])
);

LUT6 #(
   .INIT(64'h4674a83e4674a83e)  
) LUT6_inst8246 (
   .O(to_level3[470]),
   .I0(level4_in[2820]),
   .I1(level4_in[2821]),
   .I2(level4_in[2822]),
   .I3(level4_in[2823]),
   .I4(level4_in[2824]),
   .I5(level4_in[2825])
);

LUT6 #(
   .INIT(64'h81d6a7d181d6a7d1)  
) LUT6_inst8247 (
   .O(to_level3[471]),
   .I0(level4_in[2826]),
   .I1(level4_in[2827]),
   .I2(level4_in[2828]),
   .I3(level4_in[2829]),
   .I4(level4_in[2830]),
   .I5(level4_in[2831])
);

LUT6 #(
   .INIT(64'hcb278c15cb278c15)  
) LUT6_inst8248 (
   .O(to_level3[472]),
   .I0(level4_in[2832]),
   .I1(level4_in[2833]),
   .I2(level4_in[2834]),
   .I3(level4_in[2835]),
   .I4(level4_in[2836]),
   .I5(level4_in[2837])
);

LUT6 #(
   .INIT(64'hc0969214c0969214)  
) LUT6_inst8249 (
   .O(to_level3[473]),
   .I0(level4_in[2838]),
   .I1(level4_in[2839]),
   .I2(level4_in[2840]),
   .I3(level4_in[2841]),
   .I4(level4_in[2842]),
   .I5(level4_in[2843])
);

LUT6 #(
   .INIT(64'hfebd3569febd3569)  
) LUT6_inst8250 (
   .O(to_level3[474]),
   .I0(level4_in[2844]),
   .I1(level4_in[2845]),
   .I2(level4_in[2846]),
   .I3(level4_in[2847]),
   .I4(level4_in[2848]),
   .I5(level4_in[2849])
);

LUT6 #(
   .INIT(64'h2ca4db312ca4db31)  
) LUT6_inst8251 (
   .O(to_level3[475]),
   .I0(level4_in[2850]),
   .I1(level4_in[2851]),
   .I2(level4_in[2852]),
   .I3(level4_in[2853]),
   .I4(level4_in[2854]),
   .I5(level4_in[2855])
);

LUT6 #(
   .INIT(64'h78fa8be678fa8be6)  
) LUT6_inst8252 (
   .O(to_level3[476]),
   .I0(level4_in[2856]),
   .I1(level4_in[2857]),
   .I2(level4_in[2858]),
   .I3(level4_in[2859]),
   .I4(level4_in[2860]),
   .I5(level4_in[2861])
);

LUT6 #(
   .INIT(64'h6528817365288173)  
) LUT6_inst8253 (
   .O(to_level3[477]),
   .I0(level4_in[2862]),
   .I1(level4_in[2863]),
   .I2(level4_in[2864]),
   .I3(level4_in[2865]),
   .I4(level4_in[2866]),
   .I5(level4_in[2867])
);

LUT6 #(
   .INIT(64'h96c17d4396c17d43)  
) LUT6_inst8254 (
   .O(to_level3[478]),
   .I0(level4_in[2868]),
   .I1(level4_in[2869]),
   .I2(level4_in[2870]),
   .I3(level4_in[2871]),
   .I4(level4_in[2872]),
   .I5(level4_in[2873])
);

LUT6 #(
   .INIT(64'h773744eb773744eb)  
) LUT6_inst8255 (
   .O(to_level3[479]),
   .I0(level4_in[2874]),
   .I1(level4_in[2875]),
   .I2(level4_in[2876]),
   .I3(level4_in[2877]),
   .I4(level4_in[2878]),
   .I5(level4_in[2879])
);

LUT6 #(
   .INIT(64'h261f341b261f341b)  
) LUT6_inst8256 (
   .O(to_level3[480]),
   .I0(level4_in[2880]),
   .I1(level4_in[2881]),
   .I2(level4_in[2882]),
   .I3(level4_in[2883]),
   .I4(level4_in[2884]),
   .I5(level4_in[2885])
);

LUT6 #(
   .INIT(64'h733c8d9b733c8d9b)  
) LUT6_inst8257 (
   .O(to_level3[481]),
   .I0(level4_in[2886]),
   .I1(level4_in[2887]),
   .I2(level4_in[2888]),
   .I3(level4_in[2889]),
   .I4(level4_in[2890]),
   .I5(level4_in[2891])
);

LUT6 #(
   .INIT(64'hfe3657d6fe3657d6)  
) LUT6_inst8258 (
   .O(to_level3[482]),
   .I0(level4_in[2892]),
   .I1(level4_in[2893]),
   .I2(level4_in[2894]),
   .I3(level4_in[2895]),
   .I4(level4_in[2896]),
   .I5(level4_in[2897])
);

LUT6 #(
   .INIT(64'h17d5bca217d5bca2)  
) LUT6_inst8259 (
   .O(to_level3[483]),
   .I0(level4_in[2898]),
   .I1(level4_in[2899]),
   .I2(level4_in[2900]),
   .I3(level4_in[2901]),
   .I4(level4_in[2902]),
   .I5(level4_in[2903])
);

LUT6 #(
   .INIT(64'ha6c3d644a6c3d644)  
) LUT6_inst8260 (
   .O(to_level3[484]),
   .I0(level4_in[2904]),
   .I1(level4_in[2905]),
   .I2(level4_in[2906]),
   .I3(level4_in[2907]),
   .I4(level4_in[2908]),
   .I5(level4_in[2909])
);

LUT6 #(
   .INIT(64'h3b283c703b283c70)  
) LUT6_inst8261 (
   .O(to_level3[485]),
   .I0(level4_in[2910]),
   .I1(level4_in[2911]),
   .I2(level4_in[2912]),
   .I3(level4_in[2913]),
   .I4(level4_in[2914]),
   .I5(level4_in[2915])
);

LUT6 #(
   .INIT(64'hd7dc358ad7dc358a)  
) LUT6_inst8262 (
   .O(to_level3[486]),
   .I0(level4_in[2916]),
   .I1(level4_in[2917]),
   .I2(level4_in[2918]),
   .I3(level4_in[2919]),
   .I4(level4_in[2920]),
   .I5(level4_in[2921])
);

LUT6 #(
   .INIT(64'h97ef86c997ef86c9)  
) LUT6_inst8263 (
   .O(to_level3[487]),
   .I0(level4_in[2922]),
   .I1(level4_in[2923]),
   .I2(level4_in[2924]),
   .I3(level4_in[2925]),
   .I4(level4_in[2926]),
   .I5(level4_in[2927])
);

LUT6 #(
   .INIT(64'h7d49e8f47d49e8f4)  
) LUT6_inst8264 (
   .O(to_level3[488]),
   .I0(level4_in[2928]),
   .I1(level4_in[2929]),
   .I2(level4_in[2930]),
   .I3(level4_in[2931]),
   .I4(level4_in[2932]),
   .I5(level4_in[2933])
);

LUT6 #(
   .INIT(64'h807691c6807691c6)  
) LUT6_inst8265 (
   .O(to_level3[489]),
   .I0(level4_in[2934]),
   .I1(level4_in[2935]),
   .I2(level4_in[2936]),
   .I3(level4_in[2937]),
   .I4(level4_in[2938]),
   .I5(level4_in[2939])
);

LUT6 #(
   .INIT(64'hc99cd998c99cd998)  
) LUT6_inst8266 (
   .O(to_level3[490]),
   .I0(level4_in[2940]),
   .I1(level4_in[2941]),
   .I2(level4_in[2942]),
   .I3(level4_in[2943]),
   .I4(level4_in[2944]),
   .I5(level4_in[2945])
);

LUT6 #(
   .INIT(64'h631d8554631d8554)  
) LUT6_inst8267 (
   .O(to_level3[491]),
   .I0(level4_in[2946]),
   .I1(level4_in[2947]),
   .I2(level4_in[2948]),
   .I3(level4_in[2949]),
   .I4(level4_in[2950]),
   .I5(level4_in[2951])
);

LUT6 #(
   .INIT(64'h542e532c542e532c)  
) LUT6_inst8268 (
   .O(to_level3[492]),
   .I0(level4_in[2952]),
   .I1(level4_in[2953]),
   .I2(level4_in[2954]),
   .I3(level4_in[2955]),
   .I4(level4_in[2956]),
   .I5(level4_in[2957])
);

LUT6 #(
   .INIT(64'h6cdb1cef6cdb1cef)  
) LUT6_inst8269 (
   .O(to_level3[493]),
   .I0(level4_in[2958]),
   .I1(level4_in[2959]),
   .I2(level4_in[2960]),
   .I3(level4_in[2961]),
   .I4(level4_in[2962]),
   .I5(level4_in[2963])
);

LUT6 #(
   .INIT(64'h4f766ffc4f766ffc)  
) LUT6_inst8270 (
   .O(to_level3[494]),
   .I0(level4_in[2964]),
   .I1(level4_in[2965]),
   .I2(level4_in[2966]),
   .I3(level4_in[2967]),
   .I4(level4_in[2968]),
   .I5(level4_in[2969])
);

LUT6 #(
   .INIT(64'he00fb5e7e00fb5e7)  
) LUT6_inst8271 (
   .O(to_level3[495]),
   .I0(level4_in[2970]),
   .I1(level4_in[2971]),
   .I2(level4_in[2972]),
   .I3(level4_in[2973]),
   .I4(level4_in[2974]),
   .I5(level4_in[2975])
);

LUT6 #(
   .INIT(64'h9906798e9906798e)  
) LUT6_inst8272 (
   .O(to_level3[496]),
   .I0(level4_in[2976]),
   .I1(level4_in[2977]),
   .I2(level4_in[2978]),
   .I3(level4_in[2979]),
   .I4(level4_in[2980]),
   .I5(level4_in[2981])
);

LUT6 #(
   .INIT(64'h9a0398b19a0398b1)  
) LUT6_inst8273 (
   .O(to_level3[497]),
   .I0(level4_in[2982]),
   .I1(level4_in[2983]),
   .I2(level4_in[2984]),
   .I3(level4_in[2985]),
   .I4(level4_in[2986]),
   .I5(level4_in[2987])
);

LUT6 #(
   .INIT(64'hdab35f20dab35f20)  
) LUT6_inst8274 (
   .O(to_level3[498]),
   .I0(level4_in[2988]),
   .I1(level4_in[2989]),
   .I2(level4_in[2990]),
   .I3(level4_in[2991]),
   .I4(level4_in[2992]),
   .I5(level4_in[2993])
);

LUT6 #(
   .INIT(64'h63afb2d863afb2d8)  
) LUT6_inst8275 (
   .O(to_level3[499]),
   .I0(level4_in[2994]),
   .I1(level4_in[2995]),
   .I2(level4_in[2996]),
   .I3(level4_in[2997]),
   .I4(level4_in[2998]),
   .I5(level4_in[2999])
);

LUT6 #(
   .INIT(64'hadbf297dadbf297d)  
) LUT6_inst8276 (
   .O(to_level3[500]),
   .I0(level4_in[3000]),
   .I1(level4_in[3001]),
   .I2(level4_in[3002]),
   .I3(level4_in[3003]),
   .I4(level4_in[3004]),
   .I5(level4_in[3005])
);

LUT6 #(
   .INIT(64'hdd053ff0dd053ff0)  
) LUT6_inst8277 (
   .O(to_level3[501]),
   .I0(level4_in[3006]),
   .I1(level4_in[3007]),
   .I2(level4_in[3008]),
   .I3(level4_in[3009]),
   .I4(level4_in[3010]),
   .I5(level4_in[3011])
);

LUT6 #(
   .INIT(64'hadb4b14eadb4b14e)  
) LUT6_inst8278 (
   .O(to_level3[502]),
   .I0(level4_in[3012]),
   .I1(level4_in[3013]),
   .I2(level4_in[3014]),
   .I3(level4_in[3015]),
   .I4(level4_in[3016]),
   .I5(level4_in[3017])
);

LUT6 #(
   .INIT(64'h0a0e622a0a0e622a)  
) LUT6_inst8279 (
   .O(to_level3[503]),
   .I0(level4_in[3018]),
   .I1(level4_in[3019]),
   .I2(level4_in[3020]),
   .I3(level4_in[3021]),
   .I4(level4_in[3022]),
   .I5(level4_in[3023])
);

LUT6 #(
   .INIT(64'hb92e8ffcb92e8ffc)  
) LUT6_inst8280 (
   .O(to_level3[504]),
   .I0(level4_in[3024]),
   .I1(level4_in[3025]),
   .I2(level4_in[3026]),
   .I3(level4_in[3027]),
   .I4(level4_in[3028]),
   .I5(level4_in[3029])
);

LUT6 #(
   .INIT(64'hca0eb4f2ca0eb4f2)  
) LUT6_inst8281 (
   .O(to_level3[505]),
   .I0(level4_in[3030]),
   .I1(level4_in[3031]),
   .I2(level4_in[3032]),
   .I3(level4_in[3033]),
   .I4(level4_in[3034]),
   .I5(level4_in[3035])
);

LUT6 #(
   .INIT(64'h0313e5330313e533)  
) LUT6_inst8282 (
   .O(to_level3[506]),
   .I0(level4_in[3036]),
   .I1(level4_in[3037]),
   .I2(level4_in[3038]),
   .I3(level4_in[3039]),
   .I4(level4_in[3040]),
   .I5(level4_in[3041])
);

LUT6 #(
   .INIT(64'hd4562974d4562974)  
) LUT6_inst8283 (
   .O(to_level3[507]),
   .I0(level4_in[3042]),
   .I1(level4_in[3043]),
   .I2(level4_in[3044]),
   .I3(level4_in[3045]),
   .I4(level4_in[3046]),
   .I5(level4_in[3047])
);

LUT6 #(
   .INIT(64'h187125a0187125a0)  
) LUT6_inst8284 (
   .O(to_level3[508]),
   .I0(level4_in[3048]),
   .I1(level4_in[3049]),
   .I2(level4_in[3050]),
   .I3(level4_in[3051]),
   .I4(level4_in[3052]),
   .I5(level4_in[3053])
);

LUT6 #(
   .INIT(64'hfd352b9cfd352b9c)  
) LUT6_inst8285 (
   .O(to_level3[509]),
   .I0(level4_in[3054]),
   .I1(level4_in[3055]),
   .I2(level4_in[3056]),
   .I3(level4_in[3057]),
   .I4(level4_in[3058]),
   .I5(level4_in[3059])
);

LUT6 #(
   .INIT(64'h1964ab8a1964ab8a)  
) LUT6_inst8286 (
   .O(to_level3[510]),
   .I0(level4_in[3060]),
   .I1(level4_in[3061]),
   .I2(level4_in[3062]),
   .I3(level4_in[3063]),
   .I4(level4_in[3064]),
   .I5(level4_in[3065])
);

LUT6 #(
   .INIT(64'he5e9b60ce5e9b60c)  
) LUT6_inst8287 (
   .O(to_level3[511]),
   .I0(level4_in[3066]),
   .I1(level4_in[3067]),
   .I2(level4_in[3068]),
   .I3(level4_in[3069]),
   .I4(level4_in[3070]),
   .I5(level4_in[3071])
);

LUT6 #(
   .INIT(64'hc800fdfdc800fdfd)  
) LUT6_inst8288 (
   .O(to_level3[512]),
   .I0(level4_in[3072]),
   .I1(level4_in[3073]),
   .I2(level4_in[3074]),
   .I3(level4_in[3075]),
   .I4(level4_in[3076]),
   .I5(level4_in[3077])
);

LUT6 #(
   .INIT(64'hb308e086b308e086)  
) LUT6_inst8289 (
   .O(to_level3[513]),
   .I0(level4_in[3078]),
   .I1(level4_in[3079]),
   .I2(level4_in[3080]),
   .I3(level4_in[3081]),
   .I4(level4_in[3082]),
   .I5(level4_in[3083])
);

LUT6 #(
   .INIT(64'hd1a01e40d1a01e40)  
) LUT6_inst8290 (
   .O(to_level3[514]),
   .I0(level4_in[3084]),
   .I1(level4_in[3085]),
   .I2(level4_in[3086]),
   .I3(level4_in[3087]),
   .I4(level4_in[3088]),
   .I5(level4_in[3089])
);

LUT6 #(
   .INIT(64'hf85455c9f85455c9)  
) LUT6_inst8291 (
   .O(to_level3[515]),
   .I0(level4_in[3090]),
   .I1(level4_in[3091]),
   .I2(level4_in[3092]),
   .I3(level4_in[3093]),
   .I4(level4_in[3094]),
   .I5(level4_in[3095])
);

LUT6 #(
   .INIT(64'hc01a7bd7c01a7bd7)  
) LUT6_inst8292 (
   .O(to_level3[516]),
   .I0(level4_in[3096]),
   .I1(level4_in[3097]),
   .I2(level4_in[3098]),
   .I3(level4_in[3099]),
   .I4(level4_in[3100]),
   .I5(level4_in[3101])
);

LUT6 #(
   .INIT(64'h812edff7812edff7)  
) LUT6_inst8293 (
   .O(to_level3[517]),
   .I0(level4_in[3102]),
   .I1(level4_in[3103]),
   .I2(level4_in[3104]),
   .I3(level4_in[3105]),
   .I4(level4_in[3106]),
   .I5(level4_in[3107])
);

LUT6 #(
   .INIT(64'h31bce65231bce652)  
) LUT6_inst8294 (
   .O(to_level3[518]),
   .I0(level4_in[3108]),
   .I1(level4_in[3109]),
   .I2(level4_in[3110]),
   .I3(level4_in[3111]),
   .I4(level4_in[3112]),
   .I5(level4_in[3113])
);

LUT6 #(
   .INIT(64'hfa4a6062fa4a6062)  
) LUT6_inst8295 (
   .O(to_level3[519]),
   .I0(level4_in[3114]),
   .I1(level4_in[3115]),
   .I2(level4_in[3116]),
   .I3(level4_in[3117]),
   .I4(level4_in[3118]),
   .I5(level4_in[3119])
);

LUT6 #(
   .INIT(64'h06664ce306664ce3)  
) LUT6_inst8296 (
   .O(to_level3[520]),
   .I0(level4_in[3120]),
   .I1(level4_in[3121]),
   .I2(level4_in[3122]),
   .I3(level4_in[3123]),
   .I4(level4_in[3124]),
   .I5(level4_in[3125])
);

LUT6 #(
   .INIT(64'h9e494ee59e494ee5)  
) LUT6_inst8297 (
   .O(to_level3[521]),
   .I0(level4_in[3126]),
   .I1(level4_in[3127]),
   .I2(level4_in[3128]),
   .I3(level4_in[3129]),
   .I4(level4_in[3130]),
   .I5(level4_in[3131])
);

LUT6 #(
   .INIT(64'h24d3162e24d3162e)  
) LUT6_inst8298 (
   .O(to_level3[522]),
   .I0(level4_in[3132]),
   .I1(level4_in[3133]),
   .I2(level4_in[3134]),
   .I3(level4_in[3135]),
   .I4(level4_in[3136]),
   .I5(level4_in[3137])
);

LUT6 #(
   .INIT(64'h8d861b0e8d861b0e)  
) LUT6_inst8299 (
   .O(to_level3[523]),
   .I0(level4_in[3138]),
   .I1(level4_in[3139]),
   .I2(level4_in[3140]),
   .I3(level4_in[3141]),
   .I4(level4_in[3142]),
   .I5(level4_in[3143])
);

LUT6 #(
   .INIT(64'h4aa4ca694aa4ca69)  
) LUT6_inst8300 (
   .O(to_level3[524]),
   .I0(level4_in[3144]),
   .I1(level4_in[3145]),
   .I2(level4_in[3146]),
   .I3(level4_in[3147]),
   .I4(level4_in[3148]),
   .I5(level4_in[3149])
);

LUT6 #(
   .INIT(64'h075fe1f9075fe1f9)  
) LUT6_inst8301 (
   .O(to_level3[525]),
   .I0(level4_in[3150]),
   .I1(level4_in[3151]),
   .I2(level4_in[3152]),
   .I3(level4_in[3153]),
   .I4(level4_in[3154]),
   .I5(level4_in[3155])
);

LUT6 #(
   .INIT(64'h5b5affd25b5affd2)  
) LUT6_inst8302 (
   .O(to_level3[526]),
   .I0(level4_in[3156]),
   .I1(level4_in[3157]),
   .I2(level4_in[3158]),
   .I3(level4_in[3159]),
   .I4(level4_in[3160]),
   .I5(level4_in[3161])
);

LUT6 #(
   .INIT(64'h471e99a6471e99a6)  
) LUT6_inst8303 (
   .O(to_level3[527]),
   .I0(level4_in[3162]),
   .I1(level4_in[3163]),
   .I2(level4_in[3164]),
   .I3(level4_in[3165]),
   .I4(level4_in[3166]),
   .I5(level4_in[3167])
);

LUT6 #(
   .INIT(64'h4cbe7d6d4cbe7d6d)  
) LUT6_inst8304 (
   .O(to_level3[528]),
   .I0(level4_in[3168]),
   .I1(level4_in[3169]),
   .I2(level4_in[3170]),
   .I3(level4_in[3171]),
   .I4(level4_in[3172]),
   .I5(level4_in[3173])
);

LUT6 #(
   .INIT(64'hed62c84aed62c84a)  
) LUT6_inst8305 (
   .O(to_level3[529]),
   .I0(level4_in[3174]),
   .I1(level4_in[3175]),
   .I2(level4_in[3176]),
   .I3(level4_in[3177]),
   .I4(level4_in[3178]),
   .I5(level4_in[3179])
);

LUT6 #(
   .INIT(64'h8aae6f3c8aae6f3c)  
) LUT6_inst8306 (
   .O(to_level3[530]),
   .I0(level4_in[3180]),
   .I1(level4_in[3181]),
   .I2(level4_in[3182]),
   .I3(level4_in[3183]),
   .I4(level4_in[3184]),
   .I5(level4_in[3185])
);

LUT6 #(
   .INIT(64'hc51ed8d3c51ed8d3)  
) LUT6_inst8307 (
   .O(to_level3[531]),
   .I0(level4_in[3186]),
   .I1(level4_in[3187]),
   .I2(level4_in[3188]),
   .I3(level4_in[3189]),
   .I4(level4_in[3190]),
   .I5(level4_in[3191])
);

LUT6 #(
   .INIT(64'h94a5676794a56767)  
) LUT6_inst8308 (
   .O(to_level3[532]),
   .I0(level4_in[3192]),
   .I1(level4_in[3193]),
   .I2(level4_in[3194]),
   .I3(level4_in[3195]),
   .I4(level4_in[3196]),
   .I5(level4_in[3197])
);

LUT6 #(
   .INIT(64'h45ac50c345ac50c3)  
) LUT6_inst8309 (
   .O(to_level3[533]),
   .I0(level4_in[3198]),
   .I1(level4_in[3199]),
   .I2(level4_in[3200]),
   .I3(level4_in[3201]),
   .I4(level4_in[3202]),
   .I5(level4_in[3203])
);

LUT6 #(
   .INIT(64'h28759fab28759fab)  
) LUT6_inst8310 (
   .O(to_level3[534]),
   .I0(level4_in[3204]),
   .I1(level4_in[3205]),
   .I2(level4_in[3206]),
   .I3(level4_in[3207]),
   .I4(level4_in[3208]),
   .I5(level4_in[3209])
);

LUT6 #(
   .INIT(64'h55ede2dd55ede2dd)  
) LUT6_inst8311 (
   .O(to_level3[535]),
   .I0(level4_in[3210]),
   .I1(level4_in[3211]),
   .I2(level4_in[3212]),
   .I3(level4_in[3213]),
   .I4(level4_in[3214]),
   .I5(level4_in[3215])
);

LUT6 #(
   .INIT(64'hdbb2eabedbb2eabe)  
) LUT6_inst8312 (
   .O(to_level3[536]),
   .I0(level4_in[3216]),
   .I1(level4_in[3217]),
   .I2(level4_in[3218]),
   .I3(level4_in[3219]),
   .I4(level4_in[3220]),
   .I5(level4_in[3221])
);

LUT6 #(
   .INIT(64'hea7e811dea7e811d)  
) LUT6_inst8313 (
   .O(to_level3[537]),
   .I0(level4_in[3222]),
   .I1(level4_in[3223]),
   .I2(level4_in[3224]),
   .I3(level4_in[3225]),
   .I4(level4_in[3226]),
   .I5(level4_in[3227])
);

LUT6 #(
   .INIT(64'hc39c254fc39c254f)  
) LUT6_inst8314 (
   .O(to_level3[538]),
   .I0(level4_in[3228]),
   .I1(level4_in[3229]),
   .I2(level4_in[3230]),
   .I3(level4_in[3231]),
   .I4(level4_in[3232]),
   .I5(level4_in[3233])
);

LUT6 #(
   .INIT(64'h6dd88f6f6dd88f6f)  
) LUT6_inst8315 (
   .O(to_level3[539]),
   .I0(level4_in[3234]),
   .I1(level4_in[3235]),
   .I2(level4_in[3236]),
   .I3(level4_in[3237]),
   .I4(level4_in[3238]),
   .I5(level4_in[3239])
);

LUT6 #(
   .INIT(64'h5238f04a5238f04a)  
) LUT6_inst8316 (
   .O(to_level3[540]),
   .I0(level4_in[3240]),
   .I1(level4_in[3241]),
   .I2(level4_in[3242]),
   .I3(level4_in[3243]),
   .I4(level4_in[3244]),
   .I5(level4_in[3245])
);

LUT6 #(
   .INIT(64'h9973a2519973a251)  
) LUT6_inst8317 (
   .O(to_level3[541]),
   .I0(level4_in[3246]),
   .I1(level4_in[3247]),
   .I2(level4_in[3248]),
   .I3(level4_in[3249]),
   .I4(level4_in[3250]),
   .I5(level4_in[3251])
);

LUT6 #(
   .INIT(64'hbddb24d8bddb24d8)  
) LUT6_inst8318 (
   .O(to_level3[542]),
   .I0(level4_in[3252]),
   .I1(level4_in[3253]),
   .I2(level4_in[3254]),
   .I3(level4_in[3255]),
   .I4(level4_in[3256]),
   .I5(level4_in[3257])
);

LUT6 #(
   .INIT(64'h34a6823334a68233)  
) LUT6_inst8319 (
   .O(to_level3[543]),
   .I0(level4_in[3258]),
   .I1(level4_in[3259]),
   .I2(level4_in[3260]),
   .I3(level4_in[3261]),
   .I4(level4_in[3262]),
   .I5(level4_in[3263])
);

LUT6 #(
   .INIT(64'h8cc2b3a48cc2b3a4)  
) LUT6_inst8320 (
   .O(to_level3[544]),
   .I0(level4_in[3264]),
   .I1(level4_in[3265]),
   .I2(level4_in[3266]),
   .I3(level4_in[3267]),
   .I4(level4_in[3268]),
   .I5(level4_in[3269])
);

LUT6 #(
   .INIT(64'h273d6379273d6379)  
) LUT6_inst8321 (
   .O(to_level3[545]),
   .I0(level4_in[3270]),
   .I1(level4_in[3271]),
   .I2(level4_in[3272]),
   .I3(level4_in[3273]),
   .I4(level4_in[3274]),
   .I5(level4_in[3275])
);

LUT6 #(
   .INIT(64'h5c7ffcb75c7ffcb7)  
) LUT6_inst8322 (
   .O(to_level3[546]),
   .I0(level4_in[3276]),
   .I1(level4_in[3277]),
   .I2(level4_in[3278]),
   .I3(level4_in[3279]),
   .I4(level4_in[3280]),
   .I5(level4_in[3281])
);

LUT6 #(
   .INIT(64'hc9067d63c9067d63)  
) LUT6_inst8323 (
   .O(to_level3[547]),
   .I0(level4_in[3282]),
   .I1(level4_in[3283]),
   .I2(level4_in[3284]),
   .I3(level4_in[3285]),
   .I4(level4_in[3286]),
   .I5(level4_in[3287])
);

LUT6 #(
   .INIT(64'h91f2c90391f2c903)  
) LUT6_inst8324 (
   .O(to_level3[548]),
   .I0(level4_in[3288]),
   .I1(level4_in[3289]),
   .I2(level4_in[3290]),
   .I3(level4_in[3291]),
   .I4(level4_in[3292]),
   .I5(level4_in[3293])
);

LUT6 #(
   .INIT(64'h0aa8f5e20aa8f5e2)  
) LUT6_inst8325 (
   .O(to_level3[549]),
   .I0(level4_in[3294]),
   .I1(level4_in[3295]),
   .I2(level4_in[3296]),
   .I3(level4_in[3297]),
   .I4(level4_in[3298]),
   .I5(level4_in[3299])
);

LUT6 #(
   .INIT(64'hdba1770ddba1770d)  
) LUT6_inst8326 (
   .O(to_level3[550]),
   .I0(level4_in[3300]),
   .I1(level4_in[3301]),
   .I2(level4_in[3302]),
   .I3(level4_in[3303]),
   .I4(level4_in[3304]),
   .I5(level4_in[3305])
);

LUT6 #(
   .INIT(64'h4cf02bda4cf02bda)  
) LUT6_inst8327 (
   .O(to_level3[551]),
   .I0(level4_in[3306]),
   .I1(level4_in[3307]),
   .I2(level4_in[3308]),
   .I3(level4_in[3309]),
   .I4(level4_in[3310]),
   .I5(level4_in[3311])
);

LUT6 #(
   .INIT(64'hbfa53352bfa53352)  
) LUT6_inst8328 (
   .O(to_level3[552]),
   .I0(level4_in[3312]),
   .I1(level4_in[3313]),
   .I2(level4_in[3314]),
   .I3(level4_in[3315]),
   .I4(level4_in[3316]),
   .I5(level4_in[3317])
);

LUT6 #(
   .INIT(64'hceb8b1d6ceb8b1d6)  
) LUT6_inst8329 (
   .O(to_level3[553]),
   .I0(level4_in[3318]),
   .I1(level4_in[3319]),
   .I2(level4_in[3320]),
   .I3(level4_in[3321]),
   .I4(level4_in[3322]),
   .I5(level4_in[3323])
);

LUT6 #(
   .INIT(64'h48d1ef6b48d1ef6b)  
) LUT6_inst8330 (
   .O(to_level3[554]),
   .I0(level4_in[3324]),
   .I1(level4_in[3325]),
   .I2(level4_in[3326]),
   .I3(level4_in[3327]),
   .I4(level4_in[3328]),
   .I5(level4_in[3329])
);

LUT6 #(
   .INIT(64'h9474b6059474b605)  
) LUT6_inst8331 (
   .O(to_level3[555]),
   .I0(level4_in[3330]),
   .I1(level4_in[3331]),
   .I2(level4_in[3332]),
   .I3(level4_in[3333]),
   .I4(level4_in[3334]),
   .I5(level4_in[3335])
);

LUT6 #(
   .INIT(64'he7ef702be7ef702b)  
) LUT6_inst8332 (
   .O(to_level3[556]),
   .I0(level4_in[3336]),
   .I1(level4_in[3337]),
   .I2(level4_in[3338]),
   .I3(level4_in[3339]),
   .I4(level4_in[3340]),
   .I5(level4_in[3341])
);

LUT6 #(
   .INIT(64'hc499b032c499b032)  
) LUT6_inst8333 (
   .O(to_level3[557]),
   .I0(level4_in[3342]),
   .I1(level4_in[3343]),
   .I2(level4_in[3344]),
   .I3(level4_in[3345]),
   .I4(level4_in[3346]),
   .I5(level4_in[3347])
);

LUT6 #(
   .INIT(64'ha797e753a797e753)  
) LUT6_inst8334 (
   .O(to_level3[558]),
   .I0(level4_in[3348]),
   .I1(level4_in[3349]),
   .I2(level4_in[3350]),
   .I3(level4_in[3351]),
   .I4(level4_in[3352]),
   .I5(level4_in[3353])
);

LUT6 #(
   .INIT(64'h9ccbd51f9ccbd51f)  
) LUT6_inst8335 (
   .O(to_level3[559]),
   .I0(level4_in[3354]),
   .I1(level4_in[3355]),
   .I2(level4_in[3356]),
   .I3(level4_in[3357]),
   .I4(level4_in[3358]),
   .I5(level4_in[3359])
);

LUT6 #(
   .INIT(64'h2ecc7ba72ecc7ba7)  
) LUT6_inst8336 (
   .O(to_level3[560]),
   .I0(level4_in[3360]),
   .I1(level4_in[3361]),
   .I2(level4_in[3362]),
   .I3(level4_in[3363]),
   .I4(level4_in[3364]),
   .I5(level4_in[3365])
);

LUT6 #(
   .INIT(64'h61a1356161a13561)  
) LUT6_inst8337 (
   .O(to_level3[561]),
   .I0(level4_in[3366]),
   .I1(level4_in[3367]),
   .I2(level4_in[3368]),
   .I3(level4_in[3369]),
   .I4(level4_in[3370]),
   .I5(level4_in[3371])
);

LUT6 #(
   .INIT(64'he0a491c8e0a491c8)  
) LUT6_inst8338 (
   .O(to_level3[562]),
   .I0(level4_in[3372]),
   .I1(level4_in[3373]),
   .I2(level4_in[3374]),
   .I3(level4_in[3375]),
   .I4(level4_in[3376]),
   .I5(level4_in[3377])
);

LUT6 #(
   .INIT(64'h034598e6034598e6)  
) LUT6_inst8339 (
   .O(to_level3[563]),
   .I0(level4_in[3378]),
   .I1(level4_in[3379]),
   .I2(level4_in[3380]),
   .I3(level4_in[3381]),
   .I4(level4_in[3382]),
   .I5(level4_in[3383])
);

LUT6 #(
   .INIT(64'h50a35ba150a35ba1)  
) LUT6_inst8340 (
   .O(to_level3[564]),
   .I0(level4_in[3384]),
   .I1(level4_in[3385]),
   .I2(level4_in[3386]),
   .I3(level4_in[3387]),
   .I4(level4_in[3388]),
   .I5(level4_in[3389])
);

LUT6 #(
   .INIT(64'hde4cf191de4cf191)  
) LUT6_inst8341 (
   .O(to_level3[565]),
   .I0(level4_in[3390]),
   .I1(level4_in[3391]),
   .I2(level4_in[3392]),
   .I3(level4_in[3393]),
   .I4(level4_in[3394]),
   .I5(level4_in[3395])
);

LUT6 #(
   .INIT(64'he0e25b6de0e25b6d)  
) LUT6_inst8342 (
   .O(to_level3[566]),
   .I0(level4_in[3396]),
   .I1(level4_in[3397]),
   .I2(level4_in[3398]),
   .I3(level4_in[3399]),
   .I4(level4_in[3400]),
   .I5(level4_in[3401])
);

LUT6 #(
   .INIT(64'had9d5fe5ad9d5fe5)  
) LUT6_inst8343 (
   .O(to_level3[567]),
   .I0(level4_in[3402]),
   .I1(level4_in[3403]),
   .I2(level4_in[3404]),
   .I3(level4_in[3405]),
   .I4(level4_in[3406]),
   .I5(level4_in[3407])
);

LUT6 #(
   .INIT(64'h3affd4a53affd4a5)  
) LUT6_inst8344 (
   .O(to_level3[568]),
   .I0(level4_in[3408]),
   .I1(level4_in[3409]),
   .I2(level4_in[3410]),
   .I3(level4_in[3411]),
   .I4(level4_in[3412]),
   .I5(level4_in[3413])
);

LUT6 #(
   .INIT(64'h3920229f3920229f)  
) LUT6_inst8345 (
   .O(to_level3[569]),
   .I0(level4_in[3414]),
   .I1(level4_in[3415]),
   .I2(level4_in[3416]),
   .I3(level4_in[3417]),
   .I4(level4_in[3418]),
   .I5(level4_in[3419])
);

LUT6 #(
   .INIT(64'h48531e9648531e96)  
) LUT6_inst8346 (
   .O(to_level3[570]),
   .I0(level4_in[3420]),
   .I1(level4_in[3421]),
   .I2(level4_in[3422]),
   .I3(level4_in[3423]),
   .I4(level4_in[3424]),
   .I5(level4_in[3425])
);

LUT6 #(
   .INIT(64'hf264063cf264063c)  
) LUT6_inst8347 (
   .O(to_level3[571]),
   .I0(level4_in[3426]),
   .I1(level4_in[3427]),
   .I2(level4_in[3428]),
   .I3(level4_in[3429]),
   .I4(level4_in[3430]),
   .I5(level4_in[3431])
);

LUT6 #(
   .INIT(64'h704916ef704916ef)  
) LUT6_inst8348 (
   .O(to_level3[572]),
   .I0(level4_in[3432]),
   .I1(level4_in[3433]),
   .I2(level4_in[3434]),
   .I3(level4_in[3435]),
   .I4(level4_in[3436]),
   .I5(level4_in[3437])
);

LUT6 #(
   .INIT(64'h850c4fe9850c4fe9)  
) LUT6_inst8349 (
   .O(to_level3[573]),
   .I0(level4_in[3438]),
   .I1(level4_in[3439]),
   .I2(level4_in[3440]),
   .I3(level4_in[3441]),
   .I4(level4_in[3442]),
   .I5(level4_in[3443])
);

LUT6 #(
   .INIT(64'hbe301247be301247)  
) LUT6_inst8350 (
   .O(to_level3[574]),
   .I0(level4_in[3444]),
   .I1(level4_in[3445]),
   .I2(level4_in[3446]),
   .I3(level4_in[3447]),
   .I4(level4_in[3448]),
   .I5(level4_in[3449])
);

LUT6 #(
   .INIT(64'h7e86c3a87e86c3a8)  
) LUT6_inst8351 (
   .O(to_level3[575]),
   .I0(level4_in[3450]),
   .I1(level4_in[3451]),
   .I2(level4_in[3452]),
   .I3(level4_in[3453]),
   .I4(level4_in[3454]),
   .I5(level4_in[3455])
);

LUT6 #(
   .INIT(64'hab7f7f3aab7f7f3a)  
) LUT6_inst8352 (
   .O(to_level3[576]),
   .I0(level4_in[3456]),
   .I1(level4_in[3457]),
   .I2(level4_in[3458]),
   .I3(level4_in[3459]),
   .I4(level4_in[3460]),
   .I5(level4_in[3461])
);

LUT6 #(
   .INIT(64'hc9d7518ec9d7518e)  
) LUT6_inst8353 (
   .O(to_level3[577]),
   .I0(level4_in[3462]),
   .I1(level4_in[3463]),
   .I2(level4_in[3464]),
   .I3(level4_in[3465]),
   .I4(level4_in[3466]),
   .I5(level4_in[3467])
);

LUT6 #(
   .INIT(64'hbbde0a34bbde0a34)  
) LUT6_inst8354 (
   .O(to_level3[578]),
   .I0(level4_in[3468]),
   .I1(level4_in[3469]),
   .I2(level4_in[3470]),
   .I3(level4_in[3471]),
   .I4(level4_in[3472]),
   .I5(level4_in[3473])
);

LUT6 #(
   .INIT(64'h93056ca993056ca9)  
) LUT6_inst8355 (
   .O(to_level3[579]),
   .I0(level4_in[3474]),
   .I1(level4_in[3475]),
   .I2(level4_in[3476]),
   .I3(level4_in[3477]),
   .I4(level4_in[3478]),
   .I5(level4_in[3479])
);

LUT6 #(
   .INIT(64'h4667e8054667e805)  
) LUT6_inst8356 (
   .O(to_level3[580]),
   .I0(level4_in[3480]),
   .I1(level4_in[3481]),
   .I2(level4_in[3482]),
   .I3(level4_in[3483]),
   .I4(level4_in[3484]),
   .I5(level4_in[3485])
);

LUT6 #(
   .INIT(64'hb0b0a95cb0b0a95c)  
) LUT6_inst8357 (
   .O(to_level3[581]),
   .I0(level4_in[3486]),
   .I1(level4_in[3487]),
   .I2(level4_in[3488]),
   .I3(level4_in[3489]),
   .I4(level4_in[3490]),
   .I5(level4_in[3491])
);

LUT6 #(
   .INIT(64'hcfc8f5a2cfc8f5a2)  
) LUT6_inst8358 (
   .O(to_level3[582]),
   .I0(level4_in[3492]),
   .I1(level4_in[3493]),
   .I2(level4_in[3494]),
   .I3(level4_in[3495]),
   .I4(level4_in[3496]),
   .I5(level4_in[3497])
);

LUT6 #(
   .INIT(64'h970dd15c970dd15c)  
) LUT6_inst8359 (
   .O(to_level3[583]),
   .I0(level4_in[3498]),
   .I1(level4_in[3499]),
   .I2(level4_in[3500]),
   .I3(level4_in[3501]),
   .I4(level4_in[3502]),
   .I5(level4_in[3503])
);

LUT6 #(
   .INIT(64'hc232b78bc232b78b)  
) LUT6_inst8360 (
   .O(to_level3[584]),
   .I0(level4_in[3504]),
   .I1(level4_in[3505]),
   .I2(level4_in[3506]),
   .I3(level4_in[3507]),
   .I4(level4_in[3508]),
   .I5(level4_in[3509])
);

LUT6 #(
   .INIT(64'h3bef05c43bef05c4)  
) LUT6_inst8361 (
   .O(to_level3[585]),
   .I0(level4_in[3510]),
   .I1(level4_in[3511]),
   .I2(level4_in[3512]),
   .I3(level4_in[3513]),
   .I4(level4_in[3514]),
   .I5(level4_in[3515])
);

LUT6 #(
   .INIT(64'h3ca27f973ca27f97)  
) LUT6_inst8362 (
   .O(to_level3[586]),
   .I0(level4_in[3516]),
   .I1(level4_in[3517]),
   .I2(level4_in[3518]),
   .I3(level4_in[3519]),
   .I4(level4_in[3520]),
   .I5(level4_in[3521])
);

LUT6 #(
   .INIT(64'ha4e2a063a4e2a063)  
) LUT6_inst8363 (
   .O(to_level3[587]),
   .I0(level4_in[3522]),
   .I1(level4_in[3523]),
   .I2(level4_in[3524]),
   .I3(level4_in[3525]),
   .I4(level4_in[3526]),
   .I5(level4_in[3527])
);

LUT6 #(
   .INIT(64'h65188e7c65188e7c)  
) LUT6_inst8364 (
   .O(to_level3[588]),
   .I0(level4_in[3528]),
   .I1(level4_in[3529]),
   .I2(level4_in[3530]),
   .I3(level4_in[3531]),
   .I4(level4_in[3532]),
   .I5(level4_in[3533])
);

LUT6 #(
   .INIT(64'hddc4a3d4ddc4a3d4)  
) LUT6_inst8365 (
   .O(to_level3[589]),
   .I0(level4_in[3534]),
   .I1(level4_in[3535]),
   .I2(level4_in[3536]),
   .I3(level4_in[3537]),
   .I4(level4_in[3538]),
   .I5(level4_in[3539])
);

LUT6 #(
   .INIT(64'h5b58519a5b58519a)  
) LUT6_inst8366 (
   .O(to_level3[590]),
   .I0(level4_in[3540]),
   .I1(level4_in[3541]),
   .I2(level4_in[3542]),
   .I3(level4_in[3543]),
   .I4(level4_in[3544]),
   .I5(level4_in[3545])
);

LUT6 #(
   .INIT(64'he920a25ce920a25c)  
) LUT6_inst8367 (
   .O(to_level3[591]),
   .I0(level4_in[3546]),
   .I1(level4_in[3547]),
   .I2(level4_in[3548]),
   .I3(level4_in[3549]),
   .I4(level4_in[3550]),
   .I5(level4_in[3551])
);

LUT6 #(
   .INIT(64'h797a8c45797a8c45)  
) LUT6_inst8368 (
   .O(to_level3[592]),
   .I0(level4_in[3552]),
   .I1(level4_in[3553]),
   .I2(level4_in[3554]),
   .I3(level4_in[3555]),
   .I4(level4_in[3556]),
   .I5(level4_in[3557])
);

LUT6 #(
   .INIT(64'h30e80a4e30e80a4e)  
) LUT6_inst8369 (
   .O(to_level3[593]),
   .I0(level4_in[3558]),
   .I1(level4_in[3559]),
   .I2(level4_in[3560]),
   .I3(level4_in[3561]),
   .I4(level4_in[3562]),
   .I5(level4_in[3563])
);

LUT6 #(
   .INIT(64'h36bf01f036bf01f0)  
) LUT6_inst8370 (
   .O(to_level3[594]),
   .I0(level4_in[3564]),
   .I1(level4_in[3565]),
   .I2(level4_in[3566]),
   .I3(level4_in[3567]),
   .I4(level4_in[3568]),
   .I5(level4_in[3569])
);

LUT6 #(
   .INIT(64'h685e2d29685e2d29)  
) LUT6_inst8371 (
   .O(to_level3[595]),
   .I0(level4_in[3570]),
   .I1(level4_in[3571]),
   .I2(level4_in[3572]),
   .I3(level4_in[3573]),
   .I4(level4_in[3574]),
   .I5(level4_in[3575])
);

LUT6 #(
   .INIT(64'hfbd13d25fbd13d25)  
) LUT6_inst8372 (
   .O(to_level3[596]),
   .I0(level4_in[3576]),
   .I1(level4_in[3577]),
   .I2(level4_in[3578]),
   .I3(level4_in[3579]),
   .I4(level4_in[3580]),
   .I5(level4_in[3581])
);

LUT6 #(
   .INIT(64'hb10e4e82b10e4e82)  
) LUT6_inst8373 (
   .O(to_level3[597]),
   .I0(level4_in[3582]),
   .I1(level4_in[3583]),
   .I2(level4_in[3584]),
   .I3(level4_in[3585]),
   .I4(level4_in[3586]),
   .I5(level4_in[3587])
);

LUT6 #(
   .INIT(64'h0f0520b00f0520b0)  
) LUT6_inst8374 (
   .O(to_level3[598]),
   .I0(level4_in[3588]),
   .I1(level4_in[3589]),
   .I2(level4_in[3590]),
   .I3(level4_in[3591]),
   .I4(level4_in[3592]),
   .I5(level4_in[3593])
);

LUT6 #(
   .INIT(64'h0a58d58c0a58d58c)  
) LUT6_inst8375 (
   .O(to_level3[599]),
   .I0(level4_in[3594]),
   .I1(level4_in[3595]),
   .I2(level4_in[3596]),
   .I3(level4_in[3597]),
   .I4(level4_in[3598]),
   .I5(level4_in[3599])
);

LUT6 #(
   .INIT(64'hf00f78dbf00f78db)  
) LUT6_inst8376 (
   .O(to_level3[600]),
   .I0(level4_in[3600]),
   .I1(level4_in[3601]),
   .I2(level4_in[3602]),
   .I3(level4_in[3603]),
   .I4(level4_in[3604]),
   .I5(level4_in[3605])
);

LUT6 #(
   .INIT(64'hd21ea0a2d21ea0a2)  
) LUT6_inst8377 (
   .O(to_level3[601]),
   .I0(level4_in[3606]),
   .I1(level4_in[3607]),
   .I2(level4_in[3608]),
   .I3(level4_in[3609]),
   .I4(level4_in[3610]),
   .I5(level4_in[3611])
);

LUT6 #(
   .INIT(64'hab70cb53ab70cb53)  
) LUT6_inst8378 (
   .O(to_level3[602]),
   .I0(level4_in[3612]),
   .I1(level4_in[3613]),
   .I2(level4_in[3614]),
   .I3(level4_in[3615]),
   .I4(level4_in[3616]),
   .I5(level4_in[3617])
);

LUT6 #(
   .INIT(64'h9b15d8f59b15d8f5)  
) LUT6_inst8379 (
   .O(to_level3[603]),
   .I0(level4_in[3618]),
   .I1(level4_in[3619]),
   .I2(level4_in[3620]),
   .I3(level4_in[3621]),
   .I4(level4_in[3622]),
   .I5(level4_in[3623])
);

LUT6 #(
   .INIT(64'h6ddea2a76ddea2a7)  
) LUT6_inst8380 (
   .O(to_level3[604]),
   .I0(level4_in[3624]),
   .I1(level4_in[3625]),
   .I2(level4_in[3626]),
   .I3(level4_in[3627]),
   .I4(level4_in[3628]),
   .I5(level4_in[3629])
);

LUT6 #(
   .INIT(64'hca0a0e50ca0a0e50)  
) LUT6_inst8381 (
   .O(to_level3[605]),
   .I0(level4_in[3630]),
   .I1(level4_in[3631]),
   .I2(level4_in[3632]),
   .I3(level4_in[3633]),
   .I4(level4_in[3634]),
   .I5(level4_in[3635])
);

LUT6 #(
   .INIT(64'h149e9f10149e9f10)  
) LUT6_inst8382 (
   .O(to_level3[606]),
   .I0(level4_in[3636]),
   .I1(level4_in[3637]),
   .I2(level4_in[3638]),
   .I3(level4_in[3639]),
   .I4(level4_in[3640]),
   .I5(level4_in[3641])
);

LUT6 #(
   .INIT(64'heca49377eca49377)  
) LUT6_inst8383 (
   .O(to_level3[607]),
   .I0(level4_in[3642]),
   .I1(level4_in[3643]),
   .I2(level4_in[3644]),
   .I3(level4_in[3645]),
   .I4(level4_in[3646]),
   .I5(level4_in[3647])
);

LUT6 #(
   .INIT(64'h2f507cca2f507cca)  
) LUT6_inst8384 (
   .O(to_level3[608]),
   .I0(level4_in[3648]),
   .I1(level4_in[3649]),
   .I2(level4_in[3650]),
   .I3(level4_in[3651]),
   .I4(level4_in[3652]),
   .I5(level4_in[3653])
);

LUT6 #(
   .INIT(64'hc40fa3fec40fa3fe)  
) LUT6_inst8385 (
   .O(to_level3[609]),
   .I0(level4_in[3654]),
   .I1(level4_in[3655]),
   .I2(level4_in[3656]),
   .I3(level4_in[3657]),
   .I4(level4_in[3658]),
   .I5(level4_in[3659])
);

LUT6 #(
   .INIT(64'hf7e762e0f7e762e0)  
) LUT6_inst8386 (
   .O(to_level3[610]),
   .I0(level4_in[3660]),
   .I1(level4_in[3661]),
   .I2(level4_in[3662]),
   .I3(level4_in[3663]),
   .I4(level4_in[3664]),
   .I5(level4_in[3665])
);

LUT6 #(
   .INIT(64'h826a1ea5826a1ea5)  
) LUT6_inst8387 (
   .O(to_level3[611]),
   .I0(level4_in[3666]),
   .I1(level4_in[3667]),
   .I2(level4_in[3668]),
   .I3(level4_in[3669]),
   .I4(level4_in[3670]),
   .I5(level4_in[3671])
);

LUT6 #(
   .INIT(64'he79203e5e79203e5)  
) LUT6_inst8388 (
   .O(to_level3[612]),
   .I0(level4_in[3672]),
   .I1(level4_in[3673]),
   .I2(level4_in[3674]),
   .I3(level4_in[3675]),
   .I4(level4_in[3676]),
   .I5(level4_in[3677])
);

LUT6 #(
   .INIT(64'hdf7f0480df7f0480)  
) LUT6_inst8389 (
   .O(to_level3[613]),
   .I0(level4_in[3678]),
   .I1(level4_in[3679]),
   .I2(level4_in[3680]),
   .I3(level4_in[3681]),
   .I4(level4_in[3682]),
   .I5(level4_in[3683])
);

LUT6 #(
   .INIT(64'h283a976d283a976d)  
) LUT6_inst8390 (
   .O(to_level3[614]),
   .I0(level4_in[3684]),
   .I1(level4_in[3685]),
   .I2(level4_in[3686]),
   .I3(level4_in[3687]),
   .I4(level4_in[3688]),
   .I5(level4_in[3689])
);

LUT6 #(
   .INIT(64'h06a9adf206a9adf2)  
) LUT6_inst8391 (
   .O(to_level3[615]),
   .I0(level4_in[3690]),
   .I1(level4_in[3691]),
   .I2(level4_in[3692]),
   .I3(level4_in[3693]),
   .I4(level4_in[3694]),
   .I5(level4_in[3695])
);

LUT6 #(
   .INIT(64'h4917e2784917e278)  
) LUT6_inst8392 (
   .O(to_level3[616]),
   .I0(level4_in[3696]),
   .I1(level4_in[3697]),
   .I2(level4_in[3698]),
   .I3(level4_in[3699]),
   .I4(level4_in[3700]),
   .I5(level4_in[3701])
);

LUT6 #(
   .INIT(64'h1ee645b81ee645b8)  
) LUT6_inst8393 (
   .O(to_level3[617]),
   .I0(level4_in[3702]),
   .I1(level4_in[3703]),
   .I2(level4_in[3704]),
   .I3(level4_in[3705]),
   .I4(level4_in[3706]),
   .I5(level4_in[3707])
);

LUT6 #(
   .INIT(64'h2d7edfbf2d7edfbf)  
) LUT6_inst8394 (
   .O(to_level3[618]),
   .I0(level4_in[3708]),
   .I1(level4_in[3709]),
   .I2(level4_in[3710]),
   .I3(level4_in[3711]),
   .I4(level4_in[3712]),
   .I5(level4_in[3713])
);

LUT6 #(
   .INIT(64'he709e251e709e251)  
) LUT6_inst8395 (
   .O(to_level3[619]),
   .I0(level4_in[3714]),
   .I1(level4_in[3715]),
   .I2(level4_in[3716]),
   .I3(level4_in[3717]),
   .I4(level4_in[3718]),
   .I5(level4_in[3719])
);

LUT6 #(
   .INIT(64'hef4b1e66ef4b1e66)  
) LUT6_inst8396 (
   .O(to_level3[620]),
   .I0(level4_in[3720]),
   .I1(level4_in[3721]),
   .I2(level4_in[3722]),
   .I3(level4_in[3723]),
   .I4(level4_in[3724]),
   .I5(level4_in[3725])
);

LUT6 #(
   .INIT(64'h5ce8c4ea5ce8c4ea)  
) LUT6_inst8397 (
   .O(to_level3[621]),
   .I0(level4_in[3726]),
   .I1(level4_in[3727]),
   .I2(level4_in[3728]),
   .I3(level4_in[3729]),
   .I4(level4_in[3730]),
   .I5(level4_in[3731])
);

LUT6 #(
   .INIT(64'h71a577b071a577b0)  
) LUT6_inst8398 (
   .O(to_level3[622]),
   .I0(level4_in[3732]),
   .I1(level4_in[3733]),
   .I2(level4_in[3734]),
   .I3(level4_in[3735]),
   .I4(level4_in[3736]),
   .I5(level4_in[3737])
);

LUT6 #(
   .INIT(64'h67490b7767490b77)  
) LUT6_inst8399 (
   .O(to_level3[623]),
   .I0(level4_in[3738]),
   .I1(level4_in[3739]),
   .I2(level4_in[3740]),
   .I3(level4_in[3741]),
   .I4(level4_in[3742]),
   .I5(level4_in[3743])
);

LUT6 #(
   .INIT(64'h36b2eb8136b2eb81)  
) LUT6_inst8400 (
   .O(to_level3[624]),
   .I0(level4_in[3744]),
   .I1(level4_in[3745]),
   .I2(level4_in[3746]),
   .I3(level4_in[3747]),
   .I4(level4_in[3748]),
   .I5(level4_in[3749])
);

LUT6 #(
   .INIT(64'h6453600c6453600c)  
) LUT6_inst8401 (
   .O(to_level3[625]),
   .I0(level4_in[3750]),
   .I1(level4_in[3751]),
   .I2(level4_in[3752]),
   .I3(level4_in[3753]),
   .I4(level4_in[3754]),
   .I5(level4_in[3755])
);

LUT6 #(
   .INIT(64'h8608d8fc8608d8fc)  
) LUT6_inst8402 (
   .O(to_level3[626]),
   .I0(level4_in[3756]),
   .I1(level4_in[3757]),
   .I2(level4_in[3758]),
   .I3(level4_in[3759]),
   .I4(level4_in[3760]),
   .I5(level4_in[3761])
);

LUT6 #(
   .INIT(64'hfe5392a9fe5392a9)  
) LUT6_inst8403 (
   .O(to_level3[627]),
   .I0(level4_in[3762]),
   .I1(level4_in[3763]),
   .I2(level4_in[3764]),
   .I3(level4_in[3765]),
   .I4(level4_in[3766]),
   .I5(level4_in[3767])
);

LUT6 #(
   .INIT(64'h915b182c915b182c)  
) LUT6_inst8404 (
   .O(to_level3[628]),
   .I0(level4_in[3768]),
   .I1(level4_in[3769]),
   .I2(level4_in[3770]),
   .I3(level4_in[3771]),
   .I4(level4_in[3772]),
   .I5(level4_in[3773])
);

LUT6 #(
   .INIT(64'h192c5fb2192c5fb2)  
) LUT6_inst8405 (
   .O(to_level3[629]),
   .I0(level4_in[3774]),
   .I1(level4_in[3775]),
   .I2(level4_in[3776]),
   .I3(level4_in[3777]),
   .I4(level4_in[3778]),
   .I5(level4_in[3779])
);

LUT6 #(
   .INIT(64'ha00817ada00817ad)  
) LUT6_inst8406 (
   .O(to_level3[630]),
   .I0(level4_in[3780]),
   .I1(level4_in[3781]),
   .I2(level4_in[3782]),
   .I3(level4_in[3783]),
   .I4(level4_in[3784]),
   .I5(level4_in[3785])
);

LUT6 #(
   .INIT(64'h98297deb98297deb)  
) LUT6_inst8407 (
   .O(to_level3[631]),
   .I0(level4_in[3786]),
   .I1(level4_in[3787]),
   .I2(level4_in[3788]),
   .I3(level4_in[3789]),
   .I4(level4_in[3790]),
   .I5(level4_in[3791])
);

LUT6 #(
   .INIT(64'h460bd059460bd059)  
) LUT6_inst8408 (
   .O(to_level3[632]),
   .I0(level4_in[3792]),
   .I1(level4_in[3793]),
   .I2(level4_in[3794]),
   .I3(level4_in[3795]),
   .I4(level4_in[3796]),
   .I5(level4_in[3797])
);

LUT6 #(
   .INIT(64'hff713651ff713651)  
) LUT6_inst8409 (
   .O(to_level3[633]),
   .I0(level4_in[3798]),
   .I1(level4_in[3799]),
   .I2(level4_in[3800]),
   .I3(level4_in[3801]),
   .I4(level4_in[3802]),
   .I5(level4_in[3803])
);

LUT6 #(
   .INIT(64'h172e769f172e769f)  
) LUT6_inst8410 (
   .O(to_level3[634]),
   .I0(level4_in[3804]),
   .I1(level4_in[3805]),
   .I2(level4_in[3806]),
   .I3(level4_in[3807]),
   .I4(level4_in[3808]),
   .I5(level4_in[3809])
);

LUT6 #(
   .INIT(64'h75f511d475f511d4)  
) LUT6_inst8411 (
   .O(to_level3[635]),
   .I0(level4_in[3810]),
   .I1(level4_in[3811]),
   .I2(level4_in[3812]),
   .I3(level4_in[3813]),
   .I4(level4_in[3814]),
   .I5(level4_in[3815])
);

LUT6 #(
   .INIT(64'h72f0bdae72f0bdae)  
) LUT6_inst8412 (
   .O(to_level3[636]),
   .I0(level4_in[3816]),
   .I1(level4_in[3817]),
   .I2(level4_in[3818]),
   .I3(level4_in[3819]),
   .I4(level4_in[3820]),
   .I5(level4_in[3821])
);

LUT6 #(
   .INIT(64'h829829d0829829d0)  
) LUT6_inst8413 (
   .O(to_level3[637]),
   .I0(level4_in[3822]),
   .I1(level4_in[3823]),
   .I2(level4_in[3824]),
   .I3(level4_in[3825]),
   .I4(level4_in[3826]),
   .I5(level4_in[3827])
);

LUT6 #(
   .INIT(64'hfa1ec55efa1ec55e)  
) LUT6_inst8414 (
   .O(to_level3[638]),
   .I0(level4_in[3828]),
   .I1(level4_in[3829]),
   .I2(level4_in[3830]),
   .I3(level4_in[3831]),
   .I4(level4_in[3832]),
   .I5(level4_in[3833])
);

LUT6 #(
   .INIT(64'h89292cb989292cb9)  
) LUT6_inst8415 (
   .O(to_level3[639]),
   .I0(level4_in[3834]),
   .I1(level4_in[3835]),
   .I2(level4_in[3836]),
   .I3(level4_in[3837]),
   .I4(level4_in[3838]),
   .I5(level4_in[3839])
);

LUT6 #(
   .INIT(64'h3361b37e3361b37e)  
) LUT6_inst8416 (
   .O(to_level3[640]),
   .I0(level4_in[3840]),
   .I1(level4_in[3841]),
   .I2(level4_in[3842]),
   .I3(level4_in[3843]),
   .I4(level4_in[3844]),
   .I5(level4_in[3845])
);

LUT6 #(
   .INIT(64'h31ef83c431ef83c4)  
) LUT6_inst8417 (
   .O(to_level3[641]),
   .I0(level4_in[3846]),
   .I1(level4_in[3847]),
   .I2(level4_in[3848]),
   .I3(level4_in[3849]),
   .I4(level4_in[3850]),
   .I5(level4_in[3851])
);

LUT6 #(
   .INIT(64'h5ac33ef75ac33ef7)  
) LUT6_inst8418 (
   .O(to_level3[642]),
   .I0(level4_in[3852]),
   .I1(level4_in[3853]),
   .I2(level4_in[3854]),
   .I3(level4_in[3855]),
   .I4(level4_in[3856]),
   .I5(level4_in[3857])
);

LUT6 #(
   .INIT(64'hbe41cc82be41cc82)  
) LUT6_inst8419 (
   .O(to_level3[643]),
   .I0(level4_in[3858]),
   .I1(level4_in[3859]),
   .I2(level4_in[3860]),
   .I3(level4_in[3861]),
   .I4(level4_in[3862]),
   .I5(level4_in[3863])
);

LUT6 #(
   .INIT(64'h9fbd34de9fbd34de)  
) LUT6_inst8420 (
   .O(to_level3[644]),
   .I0(level4_in[3864]),
   .I1(level4_in[3865]),
   .I2(level4_in[3866]),
   .I3(level4_in[3867]),
   .I4(level4_in[3868]),
   .I5(level4_in[3869])
);

LUT6 #(
   .INIT(64'h7e1f41867e1f4186)  
) LUT6_inst8421 (
   .O(to_level3[645]),
   .I0(level4_in[3870]),
   .I1(level4_in[3871]),
   .I2(level4_in[3872]),
   .I3(level4_in[3873]),
   .I4(level4_in[3874]),
   .I5(level4_in[3875])
);

LUT6 #(
   .INIT(64'h1f1069571f106957)  
) LUT6_inst8422 (
   .O(to_level3[646]),
   .I0(level4_in[3876]),
   .I1(level4_in[3877]),
   .I2(level4_in[3878]),
   .I3(level4_in[3879]),
   .I4(level4_in[3880]),
   .I5(level4_in[3881])
);

LUT6 #(
   .INIT(64'hc1e0a8d5c1e0a8d5)  
) LUT6_inst8423 (
   .O(to_level3[647]),
   .I0(level4_in[3882]),
   .I1(level4_in[3883]),
   .I2(level4_in[3884]),
   .I3(level4_in[3885]),
   .I4(level4_in[3886]),
   .I5(level4_in[3887])
);

LUT6 #(
   .INIT(64'h6e8d0e436e8d0e43)  
) LUT6_inst8424 (
   .O(to_level3[648]),
   .I0(level4_in[3888]),
   .I1(level4_in[3889]),
   .I2(level4_in[3890]),
   .I3(level4_in[3891]),
   .I4(level4_in[3892]),
   .I5(level4_in[3893])
);

LUT6 #(
   .INIT(64'h73e8a9ec73e8a9ec)  
) LUT6_inst8425 (
   .O(to_level3[649]),
   .I0(level4_in[3894]),
   .I1(level4_in[3895]),
   .I2(level4_in[3896]),
   .I3(level4_in[3897]),
   .I4(level4_in[3898]),
   .I5(level4_in[3899])
);

LUT6 #(
   .INIT(64'h23414bfa23414bfa)  
) LUT6_inst8426 (
   .O(to_level3[650]),
   .I0(level4_in[3900]),
   .I1(level4_in[3901]),
   .I2(level4_in[3902]),
   .I3(level4_in[3903]),
   .I4(level4_in[3904]),
   .I5(level4_in[3905])
);

LUT6 #(
   .INIT(64'h65f3a7ea65f3a7ea)  
) LUT6_inst8427 (
   .O(to_level3[651]),
   .I0(level4_in[3906]),
   .I1(level4_in[3907]),
   .I2(level4_in[3908]),
   .I3(level4_in[3909]),
   .I4(level4_in[3910]),
   .I5(level4_in[3911])
);

LUT6 #(
   .INIT(64'h8d9f4b348d9f4b34)  
) LUT6_inst8428 (
   .O(to_level3[652]),
   .I0(level4_in[3912]),
   .I1(level4_in[3913]),
   .I2(level4_in[3914]),
   .I3(level4_in[3915]),
   .I4(level4_in[3916]),
   .I5(level4_in[3917])
);

LUT6 #(
   .INIT(64'h5b215e9e5b215e9e)  
) LUT6_inst8429 (
   .O(to_level3[653]),
   .I0(level4_in[3918]),
   .I1(level4_in[3919]),
   .I2(level4_in[3920]),
   .I3(level4_in[3921]),
   .I4(level4_in[3922]),
   .I5(level4_in[3923])
);

LUT6 #(
   .INIT(64'h35ab43d035ab43d0)  
) LUT6_inst8430 (
   .O(to_level3[654]),
   .I0(level4_in[3924]),
   .I1(level4_in[3925]),
   .I2(level4_in[3926]),
   .I3(level4_in[3927]),
   .I4(level4_in[3928]),
   .I5(level4_in[3929])
);

LUT6 #(
   .INIT(64'h316e2aaa316e2aaa)  
) LUT6_inst8431 (
   .O(to_level3[655]),
   .I0(level4_in[3930]),
   .I1(level4_in[3931]),
   .I2(level4_in[3932]),
   .I3(level4_in[3933]),
   .I4(level4_in[3934]),
   .I5(level4_in[3935])
);

LUT6 #(
   .INIT(64'h9fdea1869fdea186)  
) LUT6_inst8432 (
   .O(to_level3[656]),
   .I0(level4_in[3936]),
   .I1(level4_in[3937]),
   .I2(level4_in[3938]),
   .I3(level4_in[3939]),
   .I4(level4_in[3940]),
   .I5(level4_in[3941])
);

LUT6 #(
   .INIT(64'h38fc61b538fc61b5)  
) LUT6_inst8433 (
   .O(to_level3[657]),
   .I0(level4_in[3942]),
   .I1(level4_in[3943]),
   .I2(level4_in[3944]),
   .I3(level4_in[3945]),
   .I4(level4_in[3946]),
   .I5(level4_in[3947])
);

LUT6 #(
   .INIT(64'hfbba30d7fbba30d7)  
) LUT6_inst8434 (
   .O(to_level3[658]),
   .I0(level4_in[3948]),
   .I1(level4_in[3949]),
   .I2(level4_in[3950]),
   .I3(level4_in[3951]),
   .I4(level4_in[3952]),
   .I5(level4_in[3953])
);

LUT6 #(
   .INIT(64'hcf6e0fadcf6e0fad)  
) LUT6_inst8435 (
   .O(to_level3[659]),
   .I0(level4_in[3954]),
   .I1(level4_in[3955]),
   .I2(level4_in[3956]),
   .I3(level4_in[3957]),
   .I4(level4_in[3958]),
   .I5(level4_in[3959])
);

LUT6 #(
   .INIT(64'h5a4a25c05a4a25c0)  
) LUT6_inst8436 (
   .O(to_level3[660]),
   .I0(level4_in[3960]),
   .I1(level4_in[3961]),
   .I2(level4_in[3962]),
   .I3(level4_in[3963]),
   .I4(level4_in[3964]),
   .I5(level4_in[3965])
);

LUT6 #(
   .INIT(64'h0f914e490f914e49)  
) LUT6_inst8437 (
   .O(to_level3[661]),
   .I0(level4_in[3966]),
   .I1(level4_in[3967]),
   .I2(level4_in[3968]),
   .I3(level4_in[3969]),
   .I4(level4_in[3970]),
   .I5(level4_in[3971])
);

LUT6 #(
   .INIT(64'hfc044a6efc044a6e)  
) LUT6_inst8438 (
   .O(to_level3[662]),
   .I0(level4_in[3972]),
   .I1(level4_in[3973]),
   .I2(level4_in[3974]),
   .I3(level4_in[3975]),
   .I4(level4_in[3976]),
   .I5(level4_in[3977])
);

LUT6 #(
   .INIT(64'h8029611d8029611d)  
) LUT6_inst8439 (
   .O(to_level3[663]),
   .I0(level4_in[3978]),
   .I1(level4_in[3979]),
   .I2(level4_in[3980]),
   .I3(level4_in[3981]),
   .I4(level4_in[3982]),
   .I5(level4_in[3983])
);

LUT6 #(
   .INIT(64'h382e274b382e274b)  
) LUT6_inst8440 (
   .O(to_level3[664]),
   .I0(level4_in[3984]),
   .I1(level4_in[3985]),
   .I2(level4_in[3986]),
   .I3(level4_in[3987]),
   .I4(level4_in[3988]),
   .I5(level4_in[3989])
);

LUT6 #(
   .INIT(64'haa54ffd5aa54ffd5)  
) LUT6_inst8441 (
   .O(to_level3[665]),
   .I0(level4_in[3990]),
   .I1(level4_in[3991]),
   .I2(level4_in[3992]),
   .I3(level4_in[3993]),
   .I4(level4_in[3994]),
   .I5(level4_in[3995])
);

LUT6 #(
   .INIT(64'hb6782995b6782995)  
) LUT6_inst8442 (
   .O(to_level3[666]),
   .I0(level4_in[3996]),
   .I1(level4_in[3997]),
   .I2(level4_in[3998]),
   .I3(level4_in[3999]),
   .I4(level4_in[4000]),
   .I5(level4_in[4001])
);

LUT6 #(
   .INIT(64'ha83cd8e2a83cd8e2)  
) LUT6_inst8443 (
   .O(to_level3[667]),
   .I0(level4_in[4002]),
   .I1(level4_in[4003]),
   .I2(level4_in[4004]),
   .I3(level4_in[4005]),
   .I4(level4_in[4006]),
   .I5(level4_in[4007])
);

LUT6 #(
   .INIT(64'ha9da820da9da820d)  
) LUT6_inst8444 (
   .O(to_level3[668]),
   .I0(level4_in[4008]),
   .I1(level4_in[4009]),
   .I2(level4_in[4010]),
   .I3(level4_in[4011]),
   .I4(level4_in[4012]),
   .I5(level4_in[4013])
);

LUT6 #(
   .INIT(64'hd7dea872d7dea872)  
) LUT6_inst8445 (
   .O(to_level3[669]),
   .I0(level4_in[4014]),
   .I1(level4_in[4015]),
   .I2(level4_in[4016]),
   .I3(level4_in[4017]),
   .I4(level4_in[4018]),
   .I5(level4_in[4019])
);

LUT6 #(
   .INIT(64'h9afbce2b9afbce2b)  
) LUT6_inst8446 (
   .O(to_level3[670]),
   .I0(level4_in[4020]),
   .I1(level4_in[4021]),
   .I2(level4_in[4022]),
   .I3(level4_in[4023]),
   .I4(level4_in[4024]),
   .I5(level4_in[4025])
);

LUT6 #(
   .INIT(64'h8e3078988e307898)  
) LUT6_inst8447 (
   .O(to_level3[671]),
   .I0(level4_in[4026]),
   .I1(level4_in[4027]),
   .I2(level4_in[4028]),
   .I3(level4_in[4029]),
   .I4(level4_in[4030]),
   .I5(level4_in[4031])
);

LUT6 #(
   .INIT(64'hf1cb7f7ef1cb7f7e)  
) LUT6_inst8448 (
   .O(to_level3[672]),
   .I0(level4_in[4032]),
   .I1(level4_in[4033]),
   .I2(level4_in[4034]),
   .I3(level4_in[4035]),
   .I4(level4_in[4036]),
   .I5(level4_in[4037])
);

LUT6 #(
   .INIT(64'h5aa22c3a5aa22c3a)  
) LUT6_inst8449 (
   .O(to_level3[673]),
   .I0(level4_in[4038]),
   .I1(level4_in[4039]),
   .I2(level4_in[4040]),
   .I3(level4_in[4041]),
   .I4(level4_in[4042]),
   .I5(level4_in[4043])
);

LUT6 #(
   .INIT(64'hee8d9972ee8d9972)  
) LUT6_inst8450 (
   .O(to_level3[674]),
   .I0(level4_in[4044]),
   .I1(level4_in[4045]),
   .I2(level4_in[4046]),
   .I3(level4_in[4047]),
   .I4(level4_in[4048]),
   .I5(level4_in[4049])
);

LUT6 #(
   .INIT(64'h42c29f6842c29f68)  
) LUT6_inst8451 (
   .O(to_level3[675]),
   .I0(level4_in[4050]),
   .I1(level4_in[4051]),
   .I2(level4_in[4052]),
   .I3(level4_in[4053]),
   .I4(level4_in[4054]),
   .I5(level4_in[4055])
);

LUT6 #(
   .INIT(64'h68c3a5e968c3a5e9)  
) LUT6_inst8452 (
   .O(to_level3[676]),
   .I0(level4_in[4056]),
   .I1(level4_in[4057]),
   .I2(level4_in[4058]),
   .I3(level4_in[4059]),
   .I4(level4_in[4060]),
   .I5(level4_in[4061])
);

LUT6 #(
   .INIT(64'hb9bb8a79b9bb8a79)  
) LUT6_inst8453 (
   .O(to_level3[677]),
   .I0(level4_in[4062]),
   .I1(level4_in[4063]),
   .I2(level4_in[4064]),
   .I3(level4_in[4065]),
   .I4(level4_in[4066]),
   .I5(level4_in[4067])
);

LUT6 #(
   .INIT(64'hce8585aace8585aa)  
) LUT6_inst8454 (
   .O(to_level3[678]),
   .I0(level4_in[4068]),
   .I1(level4_in[4069]),
   .I2(level4_in[4070]),
   .I3(level4_in[4071]),
   .I4(level4_in[4072]),
   .I5(level4_in[4073])
);

LUT6 #(
   .INIT(64'hd40b0c1fd40b0c1f)  
) LUT6_inst8455 (
   .O(to_level3[679]),
   .I0(level4_in[4074]),
   .I1(level4_in[4075]),
   .I2(level4_in[4076]),
   .I3(level4_in[4077]),
   .I4(level4_in[4078]),
   .I5(level4_in[4079])
);

LUT6 #(
   .INIT(64'h3b9e15363b9e1536)  
) LUT6_inst8456 (
   .O(to_level3[680]),
   .I0(level4_in[4080]),
   .I1(level4_in[4081]),
   .I2(level4_in[4082]),
   .I3(level4_in[4083]),
   .I4(level4_in[4084]),
   .I5(level4_in[4085])
);

LUT6 #(
   .INIT(64'h720e4c6a720e4c6a)  
) LUT6_inst8457 (
   .O(to_level3[681]),
   .I0(level4_in[4086]),
   .I1(level4_in[4087]),
   .I2(level4_in[4088]),
   .I3(level4_in[4089]),
   .I4(level4_in[4090]),
   .I5(level4_in[4091])
);

LUT6 #(
   .INIT(64'h5854cb655854cb65)  
) LUT6_inst8458 (
   .O(to_level3[682]),
   .I0(level4_in[4092]),
   .I1(level4_in[4093]),
   .I2(level4_in[4094]),
   .I3(level4_in[4095]),
   .I4(level4_in[4096]),
   .I5(level4_in[4097])
);

LUT6 #(
   .INIT(64'h5bdb08385bdb0838)  
) LUT6_inst8459 (
   .O(to_level3[683]),
   .I0(level4_in[4098]),
   .I1(level4_in[4099]),
   .I2(level4_in[4100]),
   .I3(level4_in[4101]),
   .I4(level4_in[4102]),
   .I5(level4_in[4103])
);

LUT6 #(
   .INIT(64'h5b313eee5b313eee)  
) LUT6_inst8460 (
   .O(to_level3[684]),
   .I0(level4_in[4104]),
   .I1(level4_in[4105]),
   .I2(level4_in[4106]),
   .I3(level4_in[4107]),
   .I4(level4_in[4108]),
   .I5(level4_in[4109])
);

LUT6 #(
   .INIT(64'h04a76af904a76af9)  
) LUT6_inst8461 (
   .O(to_level3[685]),
   .I0(level4_in[4110]),
   .I1(level4_in[4111]),
   .I2(level4_in[4112]),
   .I3(level4_in[4113]),
   .I4(level4_in[4114]),
   .I5(level4_in[4115])
);

LUT6 #(
   .INIT(64'ha091ff14a091ff14)  
) LUT6_inst8462 (
   .O(to_level3[686]),
   .I0(level4_in[4116]),
   .I1(level4_in[4117]),
   .I2(level4_in[4118]),
   .I3(level4_in[4119]),
   .I4(level4_in[4120]),
   .I5(level4_in[4121])
);

LUT6 #(
   .INIT(64'h719938ff719938ff)  
) LUT6_inst8463 (
   .O(to_level3[687]),
   .I0(level4_in[4122]),
   .I1(level4_in[4123]),
   .I2(level4_in[4124]),
   .I3(level4_in[4125]),
   .I4(level4_in[4126]),
   .I5(level4_in[4127])
);

LUT6 #(
   .INIT(64'hcfd8e94dcfd8e94d)  
) LUT6_inst8464 (
   .O(to_level3[688]),
   .I0(level4_in[4128]),
   .I1(level4_in[4129]),
   .I2(level4_in[4130]),
   .I3(level4_in[4131]),
   .I4(level4_in[4132]),
   .I5(level4_in[4133])
);

LUT6 #(
   .INIT(64'ha50b2892a50b2892)  
) LUT6_inst8465 (
   .O(to_level3[689]),
   .I0(level4_in[4134]),
   .I1(level4_in[4135]),
   .I2(level4_in[4136]),
   .I3(level4_in[4137]),
   .I4(level4_in[4138]),
   .I5(level4_in[4139])
);

LUT6 #(
   .INIT(64'hadee33ccadee33cc)  
) LUT6_inst8466 (
   .O(to_level3[690]),
   .I0(level4_in[4140]),
   .I1(level4_in[4141]),
   .I2(level4_in[4142]),
   .I3(level4_in[4143]),
   .I4(level4_in[4144]),
   .I5(level4_in[4145])
);

LUT6 #(
   .INIT(64'h15a8af2115a8af21)  
) LUT6_inst8467 (
   .O(to_level3[691]),
   .I0(level4_in[4146]),
   .I1(level4_in[4147]),
   .I2(level4_in[4148]),
   .I3(level4_in[4149]),
   .I4(level4_in[4150]),
   .I5(level4_in[4151])
);

LUT6 #(
   .INIT(64'h50c9701d50c9701d)  
) LUT6_inst8468 (
   .O(to_level3[692]),
   .I0(level4_in[4152]),
   .I1(level4_in[4153]),
   .I2(level4_in[4154]),
   .I3(level4_in[4155]),
   .I4(level4_in[4156]),
   .I5(level4_in[4157])
);

LUT6 #(
   .INIT(64'had974652ad974652)  
) LUT6_inst8469 (
   .O(to_level3[693]),
   .I0(level4_in[4158]),
   .I1(level4_in[4159]),
   .I2(level4_in[4160]),
   .I3(level4_in[4161]),
   .I4(level4_in[4162]),
   .I5(level4_in[4163])
);

LUT6 #(
   .INIT(64'h0d35e41e0d35e41e)  
) LUT6_inst8470 (
   .O(to_level3[694]),
   .I0(level4_in[4164]),
   .I1(level4_in[4165]),
   .I2(level4_in[4166]),
   .I3(level4_in[4167]),
   .I4(level4_in[4168]),
   .I5(level4_in[4169])
);

LUT6 #(
   .INIT(64'hdc91bc3bdc91bc3b)  
) LUT6_inst8471 (
   .O(to_level3[695]),
   .I0(level4_in[4170]),
   .I1(level4_in[4171]),
   .I2(level4_in[4172]),
   .I3(level4_in[4173]),
   .I4(level4_in[4174]),
   .I5(level4_in[4175])
);

LUT6 #(
   .INIT(64'hee7085e9ee7085e9)  
) LUT6_inst8472 (
   .O(to_level3[696]),
   .I0(level4_in[4176]),
   .I1(level4_in[4177]),
   .I2(level4_in[4178]),
   .I3(level4_in[4179]),
   .I4(level4_in[4180]),
   .I5(level4_in[4181])
);

LUT6 #(
   .INIT(64'h0cf1f3280cf1f328)  
) LUT6_inst8473 (
   .O(to_level3[697]),
   .I0(level4_in[4182]),
   .I1(level4_in[4183]),
   .I2(level4_in[4184]),
   .I3(level4_in[4185]),
   .I4(level4_in[4186]),
   .I5(level4_in[4187])
);

LUT6 #(
   .INIT(64'h9196fd5e9196fd5e)  
) LUT6_inst8474 (
   .O(to_level3[698]),
   .I0(level4_in[4188]),
   .I1(level4_in[4189]),
   .I2(level4_in[4190]),
   .I3(level4_in[4191]),
   .I4(level4_in[4192]),
   .I5(level4_in[4193])
);

LUT6 #(
   .INIT(64'h5e075a4a5e075a4a)  
) LUT6_inst8475 (
   .O(to_level3[699]),
   .I0(level4_in[4194]),
   .I1(level4_in[4195]),
   .I2(level4_in[4196]),
   .I3(level4_in[4197]),
   .I4(level4_in[4198]),
   .I5(level4_in[4199])
);

LUT6 #(
   .INIT(64'h1c7619de1c7619de)  
) LUT6_inst8476 (
   .O(to_level3[700]),
   .I0(level4_in[4200]),
   .I1(level4_in[4201]),
   .I2(level4_in[4202]),
   .I3(level4_in[4203]),
   .I4(level4_in[4204]),
   .I5(level4_in[4205])
);

LUT6 #(
   .INIT(64'he3e7c660e3e7c660)  
) LUT6_inst8477 (
   .O(to_level3[701]),
   .I0(level4_in[4206]),
   .I1(level4_in[4207]),
   .I2(level4_in[4208]),
   .I3(level4_in[4209]),
   .I4(level4_in[4210]),
   .I5(level4_in[4211])
);

LUT6 #(
   .INIT(64'hfe2eb4a1fe2eb4a1)  
) LUT6_inst8478 (
   .O(to_level3[702]),
   .I0(level4_in[4212]),
   .I1(level4_in[4213]),
   .I2(level4_in[4214]),
   .I3(level4_in[4215]),
   .I4(level4_in[4216]),
   .I5(level4_in[4217])
);

LUT6 #(
   .INIT(64'h07d3b03e07d3b03e)  
) LUT6_inst8479 (
   .O(to_level3[703]),
   .I0(level4_in[4218]),
   .I1(level4_in[4219]),
   .I2(level4_in[4220]),
   .I3(level4_in[4221]),
   .I4(level4_in[4222]),
   .I5(level4_in[4223])
);

LUT6 #(
   .INIT(64'h81b7cad781b7cad7)  
) LUT6_inst8480 (
   .O(to_level3[704]),
   .I0(level4_in[4224]),
   .I1(level4_in[4225]),
   .I2(level4_in[4226]),
   .I3(level4_in[4227]),
   .I4(level4_in[4228]),
   .I5(level4_in[4229])
);

LUT6 #(
   .INIT(64'h3951974939519749)  
) LUT6_inst8481 (
   .O(to_level3[705]),
   .I0(level4_in[4230]),
   .I1(level4_in[4231]),
   .I2(level4_in[4232]),
   .I3(level4_in[4233]),
   .I4(level4_in[4234]),
   .I5(level4_in[4235])
);

LUT6 #(
   .INIT(64'hbe6ebb9bbe6ebb9b)  
) LUT6_inst8482 (
   .O(to_level3[706]),
   .I0(level4_in[4236]),
   .I1(level4_in[4237]),
   .I2(level4_in[4238]),
   .I3(level4_in[4239]),
   .I4(level4_in[4240]),
   .I5(level4_in[4241])
);

LUT6 #(
   .INIT(64'h5819835458198354)  
) LUT6_inst8483 (
   .O(to_level3[707]),
   .I0(level4_in[4242]),
   .I1(level4_in[4243]),
   .I2(level4_in[4244]),
   .I3(level4_in[4245]),
   .I4(level4_in[4246]),
   .I5(level4_in[4247])
);

LUT6 #(
   .INIT(64'h9bfd60419bfd6041)  
) LUT6_inst8484 (
   .O(to_level3[708]),
   .I0(level4_in[4248]),
   .I1(level4_in[4249]),
   .I2(level4_in[4250]),
   .I3(level4_in[4251]),
   .I4(level4_in[4252]),
   .I5(level4_in[4253])
);

LUT6 #(
   .INIT(64'hca6dd873ca6dd873)  
) LUT6_inst8485 (
   .O(to_level3[709]),
   .I0(level4_in[4254]),
   .I1(level4_in[4255]),
   .I2(level4_in[4256]),
   .I3(level4_in[4257]),
   .I4(level4_in[4258]),
   .I5(level4_in[4259])
);

LUT6 #(
   .INIT(64'h40a3247040a32470)  
) LUT6_inst8486 (
   .O(to_level3[710]),
   .I0(level4_in[4260]),
   .I1(level4_in[4261]),
   .I2(level4_in[4262]),
   .I3(level4_in[4263]),
   .I4(level4_in[4264]),
   .I5(level4_in[4265])
);

LUT6 #(
   .INIT(64'h88f4d4dc88f4d4dc)  
) LUT6_inst8487 (
   .O(to_level3[711]),
   .I0(level4_in[4266]),
   .I1(level4_in[4267]),
   .I2(level4_in[4268]),
   .I3(level4_in[4269]),
   .I4(level4_in[4270]),
   .I5(level4_in[4271])
);

LUT6 #(
   .INIT(64'hda65314ada65314a)  
) LUT6_inst8488 (
   .O(to_level3[712]),
   .I0(level4_in[4272]),
   .I1(level4_in[4273]),
   .I2(level4_in[4274]),
   .I3(level4_in[4275]),
   .I4(level4_in[4276]),
   .I5(level4_in[4277])
);

LUT6 #(
   .INIT(64'h4654476c4654476c)  
) LUT6_inst8489 (
   .O(to_level3[713]),
   .I0(level4_in[4278]),
   .I1(level4_in[4279]),
   .I2(level4_in[4280]),
   .I3(level4_in[4281]),
   .I4(level4_in[4282]),
   .I5(level4_in[4283])
);

LUT6 #(
   .INIT(64'he7c18a47e7c18a47)  
) LUT6_inst8490 (
   .O(to_level3[714]),
   .I0(level4_in[4284]),
   .I1(level4_in[4285]),
   .I2(level4_in[4286]),
   .I3(level4_in[4287]),
   .I4(level4_in[4288]),
   .I5(level4_in[4289])
);

LUT6 #(
   .INIT(64'hc0ca1075c0ca1075)  
) LUT6_inst8491 (
   .O(to_level3[715]),
   .I0(level4_in[4290]),
   .I1(level4_in[4291]),
   .I2(level4_in[4292]),
   .I3(level4_in[4293]),
   .I4(level4_in[4294]),
   .I5(level4_in[4295])
);

LUT6 #(
   .INIT(64'h724901b0724901b0)  
) LUT6_inst8492 (
   .O(to_level3[716]),
   .I0(level4_in[4296]),
   .I1(level4_in[4297]),
   .I2(level4_in[4298]),
   .I3(level4_in[4299]),
   .I4(level4_in[4300]),
   .I5(level4_in[4301])
);

LUT6 #(
   .INIT(64'h8196013581960135)  
) LUT6_inst8493 (
   .O(to_level3[717]),
   .I0(level4_in[4302]),
   .I1(level4_in[4303]),
   .I2(level4_in[4304]),
   .I3(level4_in[4305]),
   .I4(level4_in[4306]),
   .I5(level4_in[4307])
);

LUT6 #(
   .INIT(64'h0b63b5a60b63b5a6)  
) LUT6_inst8494 (
   .O(to_level3[718]),
   .I0(level4_in[4308]),
   .I1(level4_in[4309]),
   .I2(level4_in[4310]),
   .I3(level4_in[4311]),
   .I4(level4_in[4312]),
   .I5(level4_in[4313])
);

LUT6 #(
   .INIT(64'h4005419040054190)  
) LUT6_inst8495 (
   .O(to_level3[719]),
   .I0(level4_in[4314]),
   .I1(level4_in[4315]),
   .I2(level4_in[4316]),
   .I3(level4_in[4317]),
   .I4(level4_in[4318]),
   .I5(level4_in[4319])
);

LUT6 #(
   .INIT(64'hbfeadd00bfeadd00)  
) LUT6_inst8496 (
   .O(to_level3[720]),
   .I0(level4_in[4320]),
   .I1(level4_in[4321]),
   .I2(level4_in[4322]),
   .I3(level4_in[4323]),
   .I4(level4_in[4324]),
   .I5(level4_in[4325])
);

LUT6 #(
   .INIT(64'hf5acceaef5acceae)  
) LUT6_inst8497 (
   .O(to_level3[721]),
   .I0(level4_in[4326]),
   .I1(level4_in[4327]),
   .I2(level4_in[4328]),
   .I3(level4_in[4329]),
   .I4(level4_in[4330]),
   .I5(level4_in[4331])
);

LUT6 #(
   .INIT(64'ha8affcd3a8affcd3)  
) LUT6_inst8498 (
   .O(to_level3[722]),
   .I0(level4_in[4332]),
   .I1(level4_in[4333]),
   .I2(level4_in[4334]),
   .I3(level4_in[4335]),
   .I4(level4_in[4336]),
   .I5(level4_in[4337])
);

LUT6 #(
   .INIT(64'hfa4d8d5efa4d8d5e)  
) LUT6_inst8499 (
   .O(to_level3[723]),
   .I0(level4_in[4338]),
   .I1(level4_in[4339]),
   .I2(level4_in[4340]),
   .I3(level4_in[4341]),
   .I4(level4_in[4342]),
   .I5(level4_in[4343])
);

LUT6 #(
   .INIT(64'hcff0214bcff0214b)  
) LUT6_inst8500 (
   .O(to_level3[724]),
   .I0(level4_in[4344]),
   .I1(level4_in[4345]),
   .I2(level4_in[4346]),
   .I3(level4_in[4347]),
   .I4(level4_in[4348]),
   .I5(level4_in[4349])
);

LUT6 #(
   .INIT(64'h1f4761071f476107)  
) LUT6_inst8501 (
   .O(to_level3[725]),
   .I0(level4_in[4350]),
   .I1(level4_in[4351]),
   .I2(level4_in[4352]),
   .I3(level4_in[4353]),
   .I4(level4_in[4354]),
   .I5(level4_in[4355])
);

LUT6 #(
   .INIT(64'hfe931fc6fe931fc6)  
) LUT6_inst8502 (
   .O(to_level3[726]),
   .I0(level4_in[4356]),
   .I1(level4_in[4357]),
   .I2(level4_in[4358]),
   .I3(level4_in[4359]),
   .I4(level4_in[4360]),
   .I5(level4_in[4361])
);

LUT6 #(
   .INIT(64'hc66d976fc66d976f)  
) LUT6_inst8503 (
   .O(to_level3[727]),
   .I0(level4_in[4362]),
   .I1(level4_in[4363]),
   .I2(level4_in[4364]),
   .I3(level4_in[4365]),
   .I4(level4_in[4366]),
   .I5(level4_in[4367])
);

LUT6 #(
   .INIT(64'h841e063e841e063e)  
) LUT6_inst8504 (
   .O(to_level3[728]),
   .I0(level4_in[4368]),
   .I1(level4_in[4369]),
   .I2(level4_in[4370]),
   .I3(level4_in[4371]),
   .I4(level4_in[4372]),
   .I5(level4_in[4373])
);

LUT6 #(
   .INIT(64'h40516d8440516d84)  
) LUT6_inst8505 (
   .O(to_level3[729]),
   .I0(level4_in[4374]),
   .I1(level4_in[4375]),
   .I2(level4_in[4376]),
   .I3(level4_in[4377]),
   .I4(level4_in[4378]),
   .I5(level4_in[4379])
);

LUT6 #(
   .INIT(64'he2842d15e2842d15)  
) LUT6_inst8506 (
   .O(to_level3[730]),
   .I0(level4_in[4380]),
   .I1(level4_in[4381]),
   .I2(level4_in[4382]),
   .I3(level4_in[4383]),
   .I4(level4_in[4384]),
   .I5(level4_in[4385])
);

LUT6 #(
   .INIT(64'h916d9e26916d9e26)  
) LUT6_inst8507 (
   .O(to_level3[731]),
   .I0(level4_in[4386]),
   .I1(level4_in[4387]),
   .I2(level4_in[4388]),
   .I3(level4_in[4389]),
   .I4(level4_in[4390]),
   .I5(level4_in[4391])
);

LUT6 #(
   .INIT(64'hf52daf5af52daf5a)  
) LUT6_inst8508 (
   .O(to_level3[732]),
   .I0(level4_in[4392]),
   .I1(level4_in[4393]),
   .I2(level4_in[4394]),
   .I3(level4_in[4395]),
   .I4(level4_in[4396]),
   .I5(level4_in[4397])
);

LUT6 #(
   .INIT(64'hd0ed8ec5d0ed8ec5)  
) LUT6_inst8509 (
   .O(to_level3[733]),
   .I0(level4_in[4398]),
   .I1(level4_in[4399]),
   .I2(level4_in[4400]),
   .I3(level4_in[4401]),
   .I4(level4_in[4402]),
   .I5(level4_in[4403])
);

LUT6 #(
   .INIT(64'h4ff1b0f94ff1b0f9)  
) LUT6_inst8510 (
   .O(to_level3[734]),
   .I0(level4_in[4404]),
   .I1(level4_in[4405]),
   .I2(level4_in[4406]),
   .I3(level4_in[4407]),
   .I4(level4_in[4408]),
   .I5(level4_in[4409])
);

LUT6 #(
   .INIT(64'h2b4b0fa42b4b0fa4)  
) LUT6_inst8511 (
   .O(to_level3[735]),
   .I0(level4_in[4410]),
   .I1(level4_in[4411]),
   .I2(level4_in[4412]),
   .I3(level4_in[4413]),
   .I4(level4_in[4414]),
   .I5(level4_in[4415])
);

LUT6 #(
   .INIT(64'hf031cdb0f031cdb0)  
) LUT6_inst8512 (
   .O(to_level3[736]),
   .I0(level4_in[4416]),
   .I1(level4_in[4417]),
   .I2(level4_in[4418]),
   .I3(level4_in[4419]),
   .I4(level4_in[4420]),
   .I5(level4_in[4421])
);

LUT6 #(
   .INIT(64'hf916ff1cf916ff1c)  
) LUT6_inst8513 (
   .O(to_level3[737]),
   .I0(level4_in[4422]),
   .I1(level4_in[4423]),
   .I2(level4_in[4424]),
   .I3(level4_in[4425]),
   .I4(level4_in[4426]),
   .I5(level4_in[4427])
);

LUT6 #(
   .INIT(64'h0261a06b0261a06b)  
) LUT6_inst8514 (
   .O(to_level3[738]),
   .I0(level4_in[4428]),
   .I1(level4_in[4429]),
   .I2(level4_in[4430]),
   .I3(level4_in[4431]),
   .I4(level4_in[4432]),
   .I5(level4_in[4433])
);

LUT6 #(
   .INIT(64'h0a5ed19d0a5ed19d)  
) LUT6_inst8515 (
   .O(to_level3[739]),
   .I0(level4_in[4434]),
   .I1(level4_in[4435]),
   .I2(level4_in[4436]),
   .I3(level4_in[4437]),
   .I4(level4_in[4438]),
   .I5(level4_in[4439])
);

LUT6 #(
   .INIT(64'h43659f0043659f00)  
) LUT6_inst8516 (
   .O(to_level3[740]),
   .I0(level4_in[4440]),
   .I1(level4_in[4441]),
   .I2(level4_in[4442]),
   .I3(level4_in[4443]),
   .I4(level4_in[4444]),
   .I5(level4_in[4445])
);

LUT6 #(
   .INIT(64'haa5e569eaa5e569e)  
) LUT6_inst8517 (
   .O(to_level3[741]),
   .I0(level4_in[4446]),
   .I1(level4_in[4447]),
   .I2(level4_in[4448]),
   .I3(level4_in[4449]),
   .I4(level4_in[4450]),
   .I5(level4_in[4451])
);

LUT6 #(
   .INIT(64'hbea461d4bea461d4)  
) LUT6_inst8518 (
   .O(to_level3[742]),
   .I0(level4_in[4452]),
   .I1(level4_in[4453]),
   .I2(level4_in[4454]),
   .I3(level4_in[4455]),
   .I4(level4_in[4456]),
   .I5(level4_in[4457])
);

LUT6 #(
   .INIT(64'hc7064943c7064943)  
) LUT6_inst8519 (
   .O(to_level3[743]),
   .I0(level4_in[4458]),
   .I1(level4_in[4459]),
   .I2(level4_in[4460]),
   .I3(level4_in[4461]),
   .I4(level4_in[4462]),
   .I5(level4_in[4463])
);

LUT6 #(
   .INIT(64'h741c9daa741c9daa)  
) LUT6_inst8520 (
   .O(to_level3[744]),
   .I0(level4_in[4464]),
   .I1(level4_in[4465]),
   .I2(level4_in[4466]),
   .I3(level4_in[4467]),
   .I4(level4_in[4468]),
   .I5(level4_in[4469])
);

LUT6 #(
   .INIT(64'h0902b6fc0902b6fc)  
) LUT6_inst8521 (
   .O(to_level3[745]),
   .I0(level4_in[4470]),
   .I1(level4_in[4471]),
   .I2(level4_in[4472]),
   .I3(level4_in[4473]),
   .I4(level4_in[4474]),
   .I5(level4_in[4475])
);

LUT6 #(
   .INIT(64'hfa92a19dfa92a19d)  
) LUT6_inst8522 (
   .O(to_level3[746]),
   .I0(level4_in[4476]),
   .I1(level4_in[4477]),
   .I2(level4_in[4478]),
   .I3(level4_in[4479]),
   .I4(level4_in[4480]),
   .I5(level4_in[4481])
);

LUT6 #(
   .INIT(64'he0ea18bbe0ea18bb)  
) LUT6_inst8523 (
   .O(to_level3[747]),
   .I0(level4_in[4482]),
   .I1(level4_in[4483]),
   .I2(level4_in[4484]),
   .I3(level4_in[4485]),
   .I4(level4_in[4486]),
   .I5(level4_in[4487])
);

LUT6 #(
   .INIT(64'h1dc2cea31dc2cea3)  
) LUT6_inst8524 (
   .O(to_level3[748]),
   .I0(level4_in[4488]),
   .I1(level4_in[4489]),
   .I2(level4_in[4490]),
   .I3(level4_in[4491]),
   .I4(level4_in[4492]),
   .I5(level4_in[4493])
);

LUT6 #(
   .INIT(64'hecf67f6cecf67f6c)  
) LUT6_inst8525 (
   .O(to_level3[749]),
   .I0(level4_in[4494]),
   .I1(level4_in[4495]),
   .I2(level4_in[4496]),
   .I3(level4_in[4497]),
   .I4(level4_in[4498]),
   .I5(level4_in[4499])
);

LUT6 #(
   .INIT(64'h516a8f80516a8f80)  
) LUT6_inst8526 (
   .O(to_level3[750]),
   .I0(level4_in[4500]),
   .I1(level4_in[4501]),
   .I2(level4_in[4502]),
   .I3(level4_in[4503]),
   .I4(level4_in[4504]),
   .I5(level4_in[4505])
);

LUT6 #(
   .INIT(64'hb8bc6da7b8bc6da7)  
) LUT6_inst8527 (
   .O(to_level3[751]),
   .I0(level4_in[4506]),
   .I1(level4_in[4507]),
   .I2(level4_in[4508]),
   .I3(level4_in[4509]),
   .I4(level4_in[4510]),
   .I5(level4_in[4511])
);

LUT6 #(
   .INIT(64'hba2e76caba2e76ca)  
) LUT6_inst8528 (
   .O(to_level3[752]),
   .I0(level4_in[4512]),
   .I1(level4_in[4513]),
   .I2(level4_in[4514]),
   .I3(level4_in[4515]),
   .I4(level4_in[4516]),
   .I5(level4_in[4517])
);

LUT6 #(
   .INIT(64'h23d86d1223d86d12)  
) LUT6_inst8529 (
   .O(to_level3[753]),
   .I0(level4_in[4518]),
   .I1(level4_in[4519]),
   .I2(level4_in[4520]),
   .I3(level4_in[4521]),
   .I4(level4_in[4522]),
   .I5(level4_in[4523])
);

LUT6 #(
   .INIT(64'h3427942834279428)  
) LUT6_inst8530 (
   .O(to_level3[754]),
   .I0(level4_in[4524]),
   .I1(level4_in[4525]),
   .I2(level4_in[4526]),
   .I3(level4_in[4527]),
   .I4(level4_in[4528]),
   .I5(level4_in[4529])
);

LUT6 #(
   .INIT(64'h8755c25e8755c25e)  
) LUT6_inst8531 (
   .O(to_level3[755]),
   .I0(level4_in[4530]),
   .I1(level4_in[4531]),
   .I2(level4_in[4532]),
   .I3(level4_in[4533]),
   .I4(level4_in[4534]),
   .I5(level4_in[4535])
);

LUT6 #(
   .INIT(64'haffb6364affb6364)  
) LUT6_inst8532 (
   .O(to_level3[756]),
   .I0(level4_in[4536]),
   .I1(level4_in[4537]),
   .I2(level4_in[4538]),
   .I3(level4_in[4539]),
   .I4(level4_in[4540]),
   .I5(level4_in[4541])
);

LUT6 #(
   .INIT(64'h7cbcd9837cbcd983)  
) LUT6_inst8533 (
   .O(to_level3[757]),
   .I0(level4_in[4542]),
   .I1(level4_in[4543]),
   .I2(level4_in[4544]),
   .I3(level4_in[4545]),
   .I4(level4_in[4546]),
   .I5(level4_in[4547])
);

LUT6 #(
   .INIT(64'he769e4a0e769e4a0)  
) LUT6_inst8534 (
   .O(to_level3[758]),
   .I0(level4_in[4548]),
   .I1(level4_in[4549]),
   .I2(level4_in[4550]),
   .I3(level4_in[4551]),
   .I4(level4_in[4552]),
   .I5(level4_in[4553])
);

LUT6 #(
   .INIT(64'h78e62cc578e62cc5)  
) LUT6_inst8535 (
   .O(to_level3[759]),
   .I0(level4_in[4554]),
   .I1(level4_in[4555]),
   .I2(level4_in[4556]),
   .I3(level4_in[4557]),
   .I4(level4_in[4558]),
   .I5(level4_in[4559])
);

LUT6 #(
   .INIT(64'h2220c2642220c264)  
) LUT6_inst8536 (
   .O(to_level3[760]),
   .I0(level4_in[4560]),
   .I1(level4_in[4561]),
   .I2(level4_in[4562]),
   .I3(level4_in[4563]),
   .I4(level4_in[4564]),
   .I5(level4_in[4565])
);

LUT6 #(
   .INIT(64'h80a0670380a06703)  
) LUT6_inst8537 (
   .O(to_level3[761]),
   .I0(level4_in[4566]),
   .I1(level4_in[4567]),
   .I2(level4_in[4568]),
   .I3(level4_in[4569]),
   .I4(level4_in[4570]),
   .I5(level4_in[4571])
);

LUT6 #(
   .INIT(64'hb48bb3d3b48bb3d3)  
) LUT6_inst8538 (
   .O(to_level3[762]),
   .I0(level4_in[4572]),
   .I1(level4_in[4573]),
   .I2(level4_in[4574]),
   .I3(level4_in[4575]),
   .I4(level4_in[4576]),
   .I5(level4_in[4577])
);

LUT6 #(
   .INIT(64'h9c7ad1909c7ad190)  
) LUT6_inst8539 (
   .O(to_level3[763]),
   .I0(level4_in[4578]),
   .I1(level4_in[4579]),
   .I2(level4_in[4580]),
   .I3(level4_in[4581]),
   .I4(level4_in[4582]),
   .I5(level4_in[4583])
);

LUT6 #(
   .INIT(64'h6fea3b9e6fea3b9e)  
) LUT6_inst8540 (
   .O(to_level3[764]),
   .I0(level4_in[4584]),
   .I1(level4_in[4585]),
   .I2(level4_in[4586]),
   .I3(level4_in[4587]),
   .I4(level4_in[4588]),
   .I5(level4_in[4589])
);

LUT6 #(
   .INIT(64'hb7fb19aab7fb19aa)  
) LUT6_inst8541 (
   .O(to_level3[765]),
   .I0(level4_in[4590]),
   .I1(level4_in[4591]),
   .I2(level4_in[4592]),
   .I3(level4_in[4593]),
   .I4(level4_in[4594]),
   .I5(level4_in[4595])
);

LUT6 #(
   .INIT(64'ha86fee3ea86fee3e)  
) LUT6_inst8542 (
   .O(to_level3[766]),
   .I0(level4_in[4596]),
   .I1(level4_in[4597]),
   .I2(level4_in[4598]),
   .I3(level4_in[4599]),
   .I4(level4_in[4600]),
   .I5(level4_in[4601])
);

LUT6 #(
   .INIT(64'hf7839f16f7839f16)  
) LUT6_inst8543 (
   .O(to_level3[767]),
   .I0(level4_in[4602]),
   .I1(level4_in[4603]),
   .I2(level4_in[4604]),
   .I3(level4_in[4605]),
   .I4(level4_in[4606]),
   .I5(level4_in[4607])
);

LUT6 #(
   .INIT(64'h8562933585629335)  
) LUT6_inst8544 (
   .O(to_level3[768]),
   .I0(level4_in[4608]),
   .I1(level4_in[4609]),
   .I2(level4_in[4610]),
   .I3(level4_in[4611]),
   .I4(level4_in[4612]),
   .I5(level4_in[4613])
);

LUT6 #(
   .INIT(64'ha20b6deda20b6ded)  
) LUT6_inst8545 (
   .O(to_level3[769]),
   .I0(level4_in[4614]),
   .I1(level4_in[4615]),
   .I2(level4_in[4616]),
   .I3(level4_in[4617]),
   .I4(level4_in[4618]),
   .I5(level4_in[4619])
);

LUT6 #(
   .INIT(64'hd5b0920ed5b0920e)  
) LUT6_inst8546 (
   .O(to_level3[770]),
   .I0(level4_in[4620]),
   .I1(level4_in[4621]),
   .I2(level4_in[4622]),
   .I3(level4_in[4623]),
   .I4(level4_in[4624]),
   .I5(level4_in[4625])
);

LUT6 #(
   .INIT(64'h728c932f728c932f)  
) LUT6_inst8547 (
   .O(to_level3[771]),
   .I0(level4_in[4626]),
   .I1(level4_in[4627]),
   .I2(level4_in[4628]),
   .I3(level4_in[4629]),
   .I4(level4_in[4630]),
   .I5(level4_in[4631])
);

LUT6 #(
   .INIT(64'h7a356b4f7a356b4f)  
) LUT6_inst8548 (
   .O(to_level3[772]),
   .I0(level4_in[4632]),
   .I1(level4_in[4633]),
   .I2(level4_in[4634]),
   .I3(level4_in[4635]),
   .I4(level4_in[4636]),
   .I5(level4_in[4637])
);

LUT6 #(
   .INIT(64'h94993e1494993e14)  
) LUT6_inst8549 (
   .O(to_level3[773]),
   .I0(level4_in[4638]),
   .I1(level4_in[4639]),
   .I2(level4_in[4640]),
   .I3(level4_in[4641]),
   .I4(level4_in[4642]),
   .I5(level4_in[4643])
);

LUT6 #(
   .INIT(64'h328255ff328255ff)  
) LUT6_inst8550 (
   .O(to_level3[774]),
   .I0(level4_in[4644]),
   .I1(level4_in[4645]),
   .I2(level4_in[4646]),
   .I3(level4_in[4647]),
   .I4(level4_in[4648]),
   .I5(level4_in[4649])
);

LUT6 #(
   .INIT(64'hdb396561db396561)  
) LUT6_inst8551 (
   .O(to_level3[775]),
   .I0(level4_in[4650]),
   .I1(level4_in[4651]),
   .I2(level4_in[4652]),
   .I3(level4_in[4653]),
   .I4(level4_in[4654]),
   .I5(level4_in[4655])
);

LUT6 #(
   .INIT(64'h25db516125db5161)  
) LUT6_inst8552 (
   .O(to_level3[776]),
   .I0(level4_in[4656]),
   .I1(level4_in[4657]),
   .I2(level4_in[4658]),
   .I3(level4_in[4659]),
   .I4(level4_in[4660]),
   .I5(level4_in[4661])
);

LUT6 #(
   .INIT(64'hc433c235c433c235)  
) LUT6_inst8553 (
   .O(to_level3[777]),
   .I0(level4_in[4662]),
   .I1(level4_in[4663]),
   .I2(level4_in[4664]),
   .I3(level4_in[4665]),
   .I4(level4_in[4666]),
   .I5(level4_in[4667])
);

LUT6 #(
   .INIT(64'h9a013c9e9a013c9e)  
) LUT6_inst8554 (
   .O(to_level3[778]),
   .I0(level4_in[4668]),
   .I1(level4_in[4669]),
   .I2(level4_in[4670]),
   .I3(level4_in[4671]),
   .I4(level4_in[4672]),
   .I5(level4_in[4673])
);

LUT6 #(
   .INIT(64'hc4560b23c4560b23)  
) LUT6_inst8555 (
   .O(to_level3[779]),
   .I0(level4_in[4674]),
   .I1(level4_in[4675]),
   .I2(level4_in[4676]),
   .I3(level4_in[4677]),
   .I4(level4_in[4678]),
   .I5(level4_in[4679])
);

LUT6 #(
   .INIT(64'h5406b0f05406b0f0)  
) LUT6_inst8556 (
   .O(to_level3[780]),
   .I0(level4_in[4680]),
   .I1(level4_in[4681]),
   .I2(level4_in[4682]),
   .I3(level4_in[4683]),
   .I4(level4_in[4684]),
   .I5(level4_in[4685])
);

LUT6 #(
   .INIT(64'h50f3beba50f3beba)  
) LUT6_inst8557 (
   .O(to_level3[781]),
   .I0(level4_in[4686]),
   .I1(level4_in[4687]),
   .I2(level4_in[4688]),
   .I3(level4_in[4689]),
   .I4(level4_in[4690]),
   .I5(level4_in[4691])
);

LUT6 #(
   .INIT(64'hcc9197fbcc9197fb)  
) LUT6_inst8558 (
   .O(to_level3[782]),
   .I0(level4_in[4692]),
   .I1(level4_in[4693]),
   .I2(level4_in[4694]),
   .I3(level4_in[4695]),
   .I4(level4_in[4696]),
   .I5(level4_in[4697])
);

LUT6 #(
   .INIT(64'hf5e8d74ff5e8d74f)  
) LUT6_inst8559 (
   .O(to_level3[783]),
   .I0(level4_in[4698]),
   .I1(level4_in[4699]),
   .I2(level4_in[4700]),
   .I3(level4_in[4701]),
   .I4(level4_in[4702]),
   .I5(level4_in[4703])
);

LUT6 #(
   .INIT(64'hd9ae0fd5d9ae0fd5)  
) LUT6_inst8560 (
   .O(to_level3[784]),
   .I0(level4_in[4704]),
   .I1(level4_in[4705]),
   .I2(level4_in[4706]),
   .I3(level4_in[4707]),
   .I4(level4_in[4708]),
   .I5(level4_in[4709])
);

LUT6 #(
   .INIT(64'h67d930f967d930f9)  
) LUT6_inst8561 (
   .O(to_level3[785]),
   .I0(level4_in[4710]),
   .I1(level4_in[4711]),
   .I2(level4_in[4712]),
   .I3(level4_in[4713]),
   .I4(level4_in[4714]),
   .I5(level4_in[4715])
);

LUT6 #(
   .INIT(64'h6d9f45d36d9f45d3)  
) LUT6_inst8562 (
   .O(to_level3[786]),
   .I0(level4_in[4716]),
   .I1(level4_in[4717]),
   .I2(level4_in[4718]),
   .I3(level4_in[4719]),
   .I4(level4_in[4720]),
   .I5(level4_in[4721])
);

LUT6 #(
   .INIT(64'he80c974ce80c974c)  
) LUT6_inst8563 (
   .O(to_level3[787]),
   .I0(level4_in[4722]),
   .I1(level4_in[4723]),
   .I2(level4_in[4724]),
   .I3(level4_in[4725]),
   .I4(level4_in[4726]),
   .I5(level4_in[4727])
);

LUT6 #(
   .INIT(64'h2bd341942bd34194)  
) LUT6_inst8564 (
   .O(to_level3[788]),
   .I0(level4_in[4728]),
   .I1(level4_in[4729]),
   .I2(level4_in[4730]),
   .I3(level4_in[4731]),
   .I4(level4_in[4732]),
   .I5(level4_in[4733])
);

LUT6 #(
   .INIT(64'hf00fa7def00fa7de)  
) LUT6_inst8565 (
   .O(to_level3[789]),
   .I0(level4_in[4734]),
   .I1(level4_in[4735]),
   .I2(level4_in[4736]),
   .I3(level4_in[4737]),
   .I4(level4_in[4738]),
   .I5(level4_in[4739])
);

LUT6 #(
   .INIT(64'h05a18ec605a18ec6)  
) LUT6_inst8566 (
   .O(to_level3[790]),
   .I0(level4_in[4740]),
   .I1(level4_in[4741]),
   .I2(level4_in[4742]),
   .I3(level4_in[4743]),
   .I4(level4_in[4744]),
   .I5(level4_in[4745])
);

LUT6 #(
   .INIT(64'hed177684ed177684)  
) LUT6_inst8567 (
   .O(to_level3[791]),
   .I0(level4_in[4746]),
   .I1(level4_in[4747]),
   .I2(level4_in[4748]),
   .I3(level4_in[4749]),
   .I4(level4_in[4750]),
   .I5(level4_in[4751])
);

LUT6 #(
   .INIT(64'he3c00595e3c00595)  
) LUT6_inst8568 (
   .O(to_level3[792]),
   .I0(level4_in[4752]),
   .I1(level4_in[4753]),
   .I2(level4_in[4754]),
   .I3(level4_in[4755]),
   .I4(level4_in[4756]),
   .I5(level4_in[4757])
);

LUT6 #(
   .INIT(64'hc5f60bd0c5f60bd0)  
) LUT6_inst8569 (
   .O(to_level3[793]),
   .I0(level4_in[4758]),
   .I1(level4_in[4759]),
   .I2(level4_in[4760]),
   .I3(level4_in[4761]),
   .I4(level4_in[4762]),
   .I5(level4_in[4763])
);

LUT6 #(
   .INIT(64'h21b4d8c321b4d8c3)  
) LUT6_inst8570 (
   .O(to_level3[794]),
   .I0(level4_in[4764]),
   .I1(level4_in[4765]),
   .I2(level4_in[4766]),
   .I3(level4_in[4767]),
   .I4(level4_in[4768]),
   .I5(level4_in[4769])
);

LUT6 #(
   .INIT(64'h78771bc178771bc1)  
) LUT6_inst8571 (
   .O(to_level3[795]),
   .I0(level4_in[4770]),
   .I1(level4_in[4771]),
   .I2(level4_in[4772]),
   .I3(level4_in[4773]),
   .I4(level4_in[4774]),
   .I5(level4_in[4775])
);

LUT6 #(
   .INIT(64'h73d7f9b173d7f9b1)  
) LUT6_inst8572 (
   .O(to_level3[796]),
   .I0(level4_in[4776]),
   .I1(level4_in[4777]),
   .I2(level4_in[4778]),
   .I3(level4_in[4779]),
   .I4(level4_in[4780]),
   .I5(level4_in[4781])
);

LUT6 #(
   .INIT(64'hc4399129c4399129)  
) LUT6_inst8573 (
   .O(to_level3[797]),
   .I0(level4_in[4782]),
   .I1(level4_in[4783]),
   .I2(level4_in[4784]),
   .I3(level4_in[4785]),
   .I4(level4_in[4786]),
   .I5(level4_in[4787])
);

LUT6 #(
   .INIT(64'h2391679a2391679a)  
) LUT6_inst8574 (
   .O(to_level3[798]),
   .I0(level4_in[4788]),
   .I1(level4_in[4789]),
   .I2(level4_in[4790]),
   .I3(level4_in[4791]),
   .I4(level4_in[4792]),
   .I5(level4_in[4793])
);

LUT6 #(
   .INIT(64'hb3d4699db3d4699d)  
) LUT6_inst8575 (
   .O(to_level3[799]),
   .I0(level4_in[4794]),
   .I1(level4_in[4795]),
   .I2(level4_in[4796]),
   .I3(level4_in[4797]),
   .I4(level4_in[4798]),
   .I5(level4_in[4799])
);

LUT6 #(
   .INIT(64'h3d83657f3d83657f)  
) LUT6_inst8576 (
   .O(to_level3[800]),
   .I0(level4_in[4800]),
   .I1(level4_in[4801]),
   .I2(level4_in[4802]),
   .I3(level4_in[4803]),
   .I4(level4_in[4804]),
   .I5(level4_in[4805])
);

LUT6 #(
   .INIT(64'h705b1bb5705b1bb5)  
) LUT6_inst8577 (
   .O(to_level3[801]),
   .I0(level4_in[4806]),
   .I1(level4_in[4807]),
   .I2(level4_in[4808]),
   .I3(level4_in[4809]),
   .I4(level4_in[4810]),
   .I5(level4_in[4811])
);

LUT6 #(
   .INIT(64'h5264899c5264899c)  
) LUT6_inst8578 (
   .O(to_level3[802]),
   .I0(level4_in[4812]),
   .I1(level4_in[4813]),
   .I2(level4_in[4814]),
   .I3(level4_in[4815]),
   .I4(level4_in[4816]),
   .I5(level4_in[4817])
);

LUT6 #(
   .INIT(64'hc9edf233c9edf233)  
) LUT6_inst8579 (
   .O(to_level3[803]),
   .I0(level4_in[4818]),
   .I1(level4_in[4819]),
   .I2(level4_in[4820]),
   .I3(level4_in[4821]),
   .I4(level4_in[4822]),
   .I5(level4_in[4823])
);

LUT6 #(
   .INIT(64'h5987ef385987ef38)  
) LUT6_inst8580 (
   .O(to_level3[804]),
   .I0(level4_in[4824]),
   .I1(level4_in[4825]),
   .I2(level4_in[4826]),
   .I3(level4_in[4827]),
   .I4(level4_in[4828]),
   .I5(level4_in[4829])
);

LUT6 #(
   .INIT(64'ha147890ea147890e)  
) LUT6_inst8581 (
   .O(to_level3[805]),
   .I0(level4_in[4830]),
   .I1(level4_in[4831]),
   .I2(level4_in[4832]),
   .I3(level4_in[4833]),
   .I4(level4_in[4834]),
   .I5(level4_in[4835])
);

LUT6 #(
   .INIT(64'he7762aebe7762aeb)  
) LUT6_inst8582 (
   .O(to_level3[806]),
   .I0(level4_in[4836]),
   .I1(level4_in[4837]),
   .I2(level4_in[4838]),
   .I3(level4_in[4839]),
   .I4(level4_in[4840]),
   .I5(level4_in[4841])
);

LUT6 #(
   .INIT(64'hcea9727dcea9727d)  
) LUT6_inst8583 (
   .O(to_level3[807]),
   .I0(level4_in[4842]),
   .I1(level4_in[4843]),
   .I2(level4_in[4844]),
   .I3(level4_in[4845]),
   .I4(level4_in[4846]),
   .I5(level4_in[4847])
);

LUT6 #(
   .INIT(64'h05af99c705af99c7)  
) LUT6_inst8584 (
   .O(to_level3[808]),
   .I0(level4_in[4848]),
   .I1(level4_in[4849]),
   .I2(level4_in[4850]),
   .I3(level4_in[4851]),
   .I4(level4_in[4852]),
   .I5(level4_in[4853])
);

LUT6 #(
   .INIT(64'ha2018540a2018540)  
) LUT6_inst8585 (
   .O(to_level3[809]),
   .I0(level4_in[4854]),
   .I1(level4_in[4855]),
   .I2(level4_in[4856]),
   .I3(level4_in[4857]),
   .I4(level4_in[4858]),
   .I5(level4_in[4859])
);

LUT6 #(
   .INIT(64'hf1286346f1286346)  
) LUT6_inst8586 (
   .O(to_level3[810]),
   .I0(level4_in[4860]),
   .I1(level4_in[4861]),
   .I2(level4_in[4862]),
   .I3(level4_in[4863]),
   .I4(level4_in[4864]),
   .I5(level4_in[4865])
);

LUT6 #(
   .INIT(64'h972723d8972723d8)  
) LUT6_inst8587 (
   .O(to_level3[811]),
   .I0(level4_in[4866]),
   .I1(level4_in[4867]),
   .I2(level4_in[4868]),
   .I3(level4_in[4869]),
   .I4(level4_in[4870]),
   .I5(level4_in[4871])
);

LUT6 #(
   .INIT(64'h53ffd1a353ffd1a3)  
) LUT6_inst8588 (
   .O(to_level3[812]),
   .I0(level4_in[4872]),
   .I1(level4_in[4873]),
   .I2(level4_in[4874]),
   .I3(level4_in[4875]),
   .I4(level4_in[4876]),
   .I5(level4_in[4877])
);

LUT6 #(
   .INIT(64'hf5b60646f5b60646)  
) LUT6_inst8589 (
   .O(to_level3[813]),
   .I0(level4_in[4878]),
   .I1(level4_in[4879]),
   .I2(level4_in[4880]),
   .I3(level4_in[4881]),
   .I4(level4_in[4882]),
   .I5(level4_in[4883])
);

LUT6 #(
   .INIT(64'h661007f2661007f2)  
) LUT6_inst8590 (
   .O(to_level3[814]),
   .I0(level4_in[4884]),
   .I1(level4_in[4885]),
   .I2(level4_in[4886]),
   .I3(level4_in[4887]),
   .I4(level4_in[4888]),
   .I5(level4_in[4889])
);

LUT6 #(
   .INIT(64'h2f92a9802f92a980)  
) LUT6_inst8591 (
   .O(to_level3[815]),
   .I0(level4_in[4890]),
   .I1(level4_in[4891]),
   .I2(level4_in[4892]),
   .I3(level4_in[4893]),
   .I4(level4_in[4894]),
   .I5(level4_in[4895])
);

LUT6 #(
   .INIT(64'h2793812927938129)  
) LUT6_inst8592 (
   .O(to_level3[816]),
   .I0(level4_in[4896]),
   .I1(level4_in[4897]),
   .I2(level4_in[4898]),
   .I3(level4_in[4899]),
   .I4(level4_in[4900]),
   .I5(level4_in[4901])
);

LUT6 #(
   .INIT(64'hedba418dedba418d)  
) LUT6_inst8593 (
   .O(to_level3[817]),
   .I0(level4_in[4902]),
   .I1(level4_in[4903]),
   .I2(level4_in[4904]),
   .I3(level4_in[4905]),
   .I4(level4_in[4906]),
   .I5(level4_in[4907])
);

LUT6 #(
   .INIT(64'h4be1191f4be1191f)  
) LUT6_inst8594 (
   .O(to_level3[818]),
   .I0(level4_in[4908]),
   .I1(level4_in[4909]),
   .I2(level4_in[4910]),
   .I3(level4_in[4911]),
   .I4(level4_in[4912]),
   .I5(level4_in[4913])
);

LUT6 #(
   .INIT(64'h256a0841256a0841)  
) LUT6_inst8595 (
   .O(to_level3[819]),
   .I0(level4_in[4914]),
   .I1(level4_in[4915]),
   .I2(level4_in[4916]),
   .I3(level4_in[4917]),
   .I4(level4_in[4918]),
   .I5(level4_in[4919])
);

LUT6 #(
   .INIT(64'h7cd2f3027cd2f302)  
) LUT6_inst8596 (
   .O(to_level3[820]),
   .I0(level4_in[4920]),
   .I1(level4_in[4921]),
   .I2(level4_in[4922]),
   .I3(level4_in[4923]),
   .I4(level4_in[4924]),
   .I5(level4_in[4925])
);

LUT6 #(
   .INIT(64'h956a0623956a0623)  
) LUT6_inst8597 (
   .O(to_level3[821]),
   .I0(level4_in[4926]),
   .I1(level4_in[4927]),
   .I2(level4_in[4928]),
   .I3(level4_in[4929]),
   .I4(level4_in[4930]),
   .I5(level4_in[4931])
);

LUT6 #(
   .INIT(64'h6f9406526f940652)  
) LUT6_inst8598 (
   .O(to_level3[822]),
   .I0(level4_in[4932]),
   .I1(level4_in[4933]),
   .I2(level4_in[4934]),
   .I3(level4_in[4935]),
   .I4(level4_in[4936]),
   .I5(level4_in[4937])
);

LUT6 #(
   .INIT(64'h5d28aea95d28aea9)  
) LUT6_inst8599 (
   .O(to_level3[823]),
   .I0(level4_in[4938]),
   .I1(level4_in[4939]),
   .I2(level4_in[4940]),
   .I3(level4_in[4941]),
   .I4(level4_in[4942]),
   .I5(level4_in[4943])
);

LUT6 #(
   .INIT(64'hf229c8dbf229c8db)  
) LUT6_inst8600 (
   .O(to_level3[824]),
   .I0(level4_in[4944]),
   .I1(level4_in[4945]),
   .I2(level4_in[4946]),
   .I3(level4_in[4947]),
   .I4(level4_in[4948]),
   .I5(level4_in[4949])
);

LUT6 #(
   .INIT(64'h5b8e73f35b8e73f3)  
) LUT6_inst8601 (
   .O(to_level3[825]),
   .I0(level4_in[4950]),
   .I1(level4_in[4951]),
   .I2(level4_in[4952]),
   .I3(level4_in[4953]),
   .I4(level4_in[4954]),
   .I5(level4_in[4955])
);

LUT6 #(
   .INIT(64'h621ba7fe621ba7fe)  
) LUT6_inst8602 (
   .O(to_level3[826]),
   .I0(level4_in[4956]),
   .I1(level4_in[4957]),
   .I2(level4_in[4958]),
   .I3(level4_in[4959]),
   .I4(level4_in[4960]),
   .I5(level4_in[4961])
);

LUT6 #(
   .INIT(64'h407f76c5407f76c5)  
) LUT6_inst8603 (
   .O(to_level3[827]),
   .I0(level4_in[4962]),
   .I1(level4_in[4963]),
   .I2(level4_in[4964]),
   .I3(level4_in[4965]),
   .I4(level4_in[4966]),
   .I5(level4_in[4967])
);

LUT6 #(
   .INIT(64'h5b1e02ce5b1e02ce)  
) LUT6_inst8604 (
   .O(to_level3[828]),
   .I0(level4_in[4968]),
   .I1(level4_in[4969]),
   .I2(level4_in[4970]),
   .I3(level4_in[4971]),
   .I4(level4_in[4972]),
   .I5(level4_in[4973])
);

LUT6 #(
   .INIT(64'hf0c2207df0c2207d)  
) LUT6_inst8605 (
   .O(to_level3[829]),
   .I0(level4_in[4974]),
   .I1(level4_in[4975]),
   .I2(level4_in[4976]),
   .I3(level4_in[4977]),
   .I4(level4_in[4978]),
   .I5(level4_in[4979])
);

LUT6 #(
   .INIT(64'h0ab154170ab15417)  
) LUT6_inst8606 (
   .O(to_level3[830]),
   .I0(level4_in[4980]),
   .I1(level4_in[4981]),
   .I2(level4_in[4982]),
   .I3(level4_in[4983]),
   .I4(level4_in[4984]),
   .I5(level4_in[4985])
);

LUT6 #(
   .INIT(64'h694ab953694ab953)  
) LUT6_inst8607 (
   .O(to_level3[831]),
   .I0(level4_in[4986]),
   .I1(level4_in[4987]),
   .I2(level4_in[4988]),
   .I3(level4_in[4989]),
   .I4(level4_in[4990]),
   .I5(level4_in[4991])
);

LUT6 #(
   .INIT(64'h3f9f3ea83f9f3ea8)  
) LUT6_inst8608 (
   .O(to_level3[832]),
   .I0(level4_in[4992]),
   .I1(level4_in[4993]),
   .I2(level4_in[4994]),
   .I3(level4_in[4995]),
   .I4(level4_in[4996]),
   .I5(level4_in[4997])
);

LUT6 #(
   .INIT(64'h9d1f04bf9d1f04bf)  
) LUT6_inst8609 (
   .O(to_level3[833]),
   .I0(level4_in[4998]),
   .I1(level4_in[4999]),
   .I2(level4_in[5000]),
   .I3(level4_in[5001]),
   .I4(level4_in[5002]),
   .I5(level4_in[5003])
);

LUT6 #(
   .INIT(64'hb1b8b141b1b8b141)  
) LUT6_inst8610 (
   .O(to_level3[834]),
   .I0(level4_in[5004]),
   .I1(level4_in[5005]),
   .I2(level4_in[5006]),
   .I3(level4_in[5007]),
   .I4(level4_in[5008]),
   .I5(level4_in[5009])
);

LUT6 #(
   .INIT(64'h1b9b0ae31b9b0ae3)  
) LUT6_inst8611 (
   .O(to_level3[835]),
   .I0(level4_in[5010]),
   .I1(level4_in[5011]),
   .I2(level4_in[5012]),
   .I3(level4_in[5013]),
   .I4(level4_in[5014]),
   .I5(level4_in[5015])
);

LUT6 #(
   .INIT(64'h1b7545e71b7545e7)  
) LUT6_inst8612 (
   .O(to_level3[836]),
   .I0(level4_in[5016]),
   .I1(level4_in[5017]),
   .I2(level4_in[5018]),
   .I3(level4_in[5019]),
   .I4(level4_in[5020]),
   .I5(level4_in[5021])
);

LUT6 #(
   .INIT(64'hfc927288fc927288)  
) LUT6_inst8613 (
   .O(to_level3[837]),
   .I0(level4_in[5022]),
   .I1(level4_in[5023]),
   .I2(level4_in[5024]),
   .I3(level4_in[5025]),
   .I4(level4_in[5026]),
   .I5(level4_in[5027])
);

LUT6 #(
   .INIT(64'hf6acebd2f6acebd2)  
) LUT6_inst8614 (
   .O(to_level3[838]),
   .I0(level4_in[5028]),
   .I1(level4_in[5029]),
   .I2(level4_in[5030]),
   .I3(level4_in[5031]),
   .I4(level4_in[5032]),
   .I5(level4_in[5033])
);

LUT6 #(
   .INIT(64'hba9e6b84ba9e6b84)  
) LUT6_inst8615 (
   .O(to_level3[839]),
   .I0(level4_in[5034]),
   .I1(level4_in[5035]),
   .I2(level4_in[5036]),
   .I3(level4_in[5037]),
   .I4(level4_in[5038]),
   .I5(level4_in[5039])
);

LUT6 #(
   .INIT(64'h40cf6ec740cf6ec7)  
) LUT6_inst8616 (
   .O(to_level3[840]),
   .I0(level4_in[5040]),
   .I1(level4_in[5041]),
   .I2(level4_in[5042]),
   .I3(level4_in[5043]),
   .I4(level4_in[5044]),
   .I5(level4_in[5045])
);

LUT6 #(
   .INIT(64'hdd962857dd962857)  
) LUT6_inst8617 (
   .O(to_level3[841]),
   .I0(level4_in[5046]),
   .I1(level4_in[5047]),
   .I2(level4_in[5048]),
   .I3(level4_in[5049]),
   .I4(level4_in[5050]),
   .I5(level4_in[5051])
);

LUT6 #(
   .INIT(64'h1b2151df1b2151df)  
) LUT6_inst8618 (
   .O(to_level3[842]),
   .I0(level4_in[5052]),
   .I1(level4_in[5053]),
   .I2(level4_in[5054]),
   .I3(level4_in[5055]),
   .I4(level4_in[5056]),
   .I5(level4_in[5057])
);

LUT6 #(
   .INIT(64'h728878e4728878e4)  
) LUT6_inst8619 (
   .O(to_level3[843]),
   .I0(level4_in[5058]),
   .I1(level4_in[5059]),
   .I2(level4_in[5060]),
   .I3(level4_in[5061]),
   .I4(level4_in[5062]),
   .I5(level4_in[5063])
);

LUT6 #(
   .INIT(64'h22d659f622d659f6)  
) LUT6_inst8620 (
   .O(to_level3[844]),
   .I0(level4_in[5064]),
   .I1(level4_in[5065]),
   .I2(level4_in[5066]),
   .I3(level4_in[5067]),
   .I4(level4_in[5068]),
   .I5(level4_in[5069])
);

LUT6 #(
   .INIT(64'hd668622cd668622c)  
) LUT6_inst8621 (
   .O(to_level3[845]),
   .I0(level4_in[5070]),
   .I1(level4_in[5071]),
   .I2(level4_in[5072]),
   .I3(level4_in[5073]),
   .I4(level4_in[5074]),
   .I5(level4_in[5075])
);

LUT6 #(
   .INIT(64'h781309ce781309ce)  
) LUT6_inst8622 (
   .O(to_level3[846]),
   .I0(level4_in[5076]),
   .I1(level4_in[5077]),
   .I2(level4_in[5078]),
   .I3(level4_in[5079]),
   .I4(level4_in[5080]),
   .I5(level4_in[5081])
);

LUT6 #(
   .INIT(64'h6105fc956105fc95)  
) LUT6_inst8623 (
   .O(to_level3[847]),
   .I0(level4_in[5082]),
   .I1(level4_in[5083]),
   .I2(level4_in[5084]),
   .I3(level4_in[5085]),
   .I4(level4_in[5086]),
   .I5(level4_in[5087])
);

LUT6 #(
   .INIT(64'hed1937e2ed1937e2)  
) LUT6_inst8624 (
   .O(to_level3[848]),
   .I0(level4_in[5088]),
   .I1(level4_in[5089]),
   .I2(level4_in[5090]),
   .I3(level4_in[5091]),
   .I4(level4_in[5092]),
   .I5(level4_in[5093])
);

LUT6 #(
   .INIT(64'hae93b9c8ae93b9c8)  
) LUT6_inst8625 (
   .O(to_level3[849]),
   .I0(level4_in[5094]),
   .I1(level4_in[5095]),
   .I2(level4_in[5096]),
   .I3(level4_in[5097]),
   .I4(level4_in[5098]),
   .I5(level4_in[5099])
);

LUT6 #(
   .INIT(64'h1a692b071a692b07)  
) LUT6_inst8626 (
   .O(to_level3[850]),
   .I0(level4_in[5100]),
   .I1(level4_in[5101]),
   .I2(level4_in[5102]),
   .I3(level4_in[5103]),
   .I4(level4_in[5104]),
   .I5(level4_in[5105])
);

LUT6 #(
   .INIT(64'h899a3d77899a3d77)  
) LUT6_inst8627 (
   .O(to_level3[851]),
   .I0(level4_in[5106]),
   .I1(level4_in[5107]),
   .I2(level4_in[5108]),
   .I3(level4_in[5109]),
   .I4(level4_in[5110]),
   .I5(level4_in[5111])
);

LUT6 #(
   .INIT(64'hadf283cbadf283cb)  
) LUT6_inst8628 (
   .O(to_level3[852]),
   .I0(level4_in[5112]),
   .I1(level4_in[5113]),
   .I2(level4_in[5114]),
   .I3(level4_in[5115]),
   .I4(level4_in[5116]),
   .I5(level4_in[5117])
);

LUT6 #(
   .INIT(64'h94f9009b94f9009b)  
) LUT6_inst8629 (
   .O(to_level3[853]),
   .I0(level4_in[5118]),
   .I1(level4_in[5119]),
   .I2(level4_in[5120]),
   .I3(level4_in[5121]),
   .I4(level4_in[5122]),
   .I5(level4_in[5123])
);

LUT6 #(
   .INIT(64'h214e866f214e866f)  
) LUT6_inst8630 (
   .O(to_level3[854]),
   .I0(level4_in[5124]),
   .I1(level4_in[5125]),
   .I2(level4_in[5126]),
   .I3(level4_in[5127]),
   .I4(level4_in[5128]),
   .I5(level4_in[5129])
);

LUT6 #(
   .INIT(64'hd425fe6cd425fe6c)  
) LUT6_inst8631 (
   .O(to_level3[855]),
   .I0(level4_in[5130]),
   .I1(level4_in[5131]),
   .I2(level4_in[5132]),
   .I3(level4_in[5133]),
   .I4(level4_in[5134]),
   .I5(level4_in[5135])
);

LUT6 #(
   .INIT(64'h6744355f6744355f)  
) LUT6_inst8632 (
   .O(to_level3[856]),
   .I0(level4_in[5136]),
   .I1(level4_in[5137]),
   .I2(level4_in[5138]),
   .I3(level4_in[5139]),
   .I4(level4_in[5140]),
   .I5(level4_in[5141])
);

LUT6 #(
   .INIT(64'h2a51d8a82a51d8a8)  
) LUT6_inst8633 (
   .O(to_level3[857]),
   .I0(level4_in[5142]),
   .I1(level4_in[5143]),
   .I2(level4_in[5144]),
   .I3(level4_in[5145]),
   .I4(level4_in[5146]),
   .I5(level4_in[5147])
);

LUT6 #(
   .INIT(64'h92e94aaf92e94aaf)  
) LUT6_inst8634 (
   .O(to_level3[858]),
   .I0(level4_in[5148]),
   .I1(level4_in[5149]),
   .I2(level4_in[5150]),
   .I3(level4_in[5151]),
   .I4(level4_in[5152]),
   .I5(level4_in[5153])
);

LUT6 #(
   .INIT(64'h2d8b3db42d8b3db4)  
) LUT6_inst8635 (
   .O(to_level3[859]),
   .I0(level4_in[5154]),
   .I1(level4_in[5155]),
   .I2(level4_in[5156]),
   .I3(level4_in[5157]),
   .I4(level4_in[5158]),
   .I5(level4_in[5159])
);

LUT6 #(
   .INIT(64'h21e8810f21e8810f)  
) LUT6_inst8636 (
   .O(to_level3[860]),
   .I0(level4_in[5160]),
   .I1(level4_in[5161]),
   .I2(level4_in[5162]),
   .I3(level4_in[5163]),
   .I4(level4_in[5164]),
   .I5(level4_in[5165])
);

LUT6 #(
   .INIT(64'h95c1e0b095c1e0b0)  
) LUT6_inst8637 (
   .O(to_level3[861]),
   .I0(level4_in[5166]),
   .I1(level4_in[5167]),
   .I2(level4_in[5168]),
   .I3(level4_in[5169]),
   .I4(level4_in[5170]),
   .I5(level4_in[5171])
);

LUT6 #(
   .INIT(64'h47d9d1ee47d9d1ee)  
) LUT6_inst8638 (
   .O(to_level3[862]),
   .I0(level4_in[5172]),
   .I1(level4_in[5173]),
   .I2(level4_in[5174]),
   .I3(level4_in[5175]),
   .I4(level4_in[5176]),
   .I5(level4_in[5177])
);

LUT6 #(
   .INIT(64'h24fd977324fd9773)  
) LUT6_inst8639 (
   .O(to_level3[863]),
   .I0(level4_in[5178]),
   .I1(level4_in[5179]),
   .I2(level4_in[5180]),
   .I3(level4_in[5181]),
   .I4(level4_in[5182]),
   .I5(level4_in[5183])
);

LUT6 #(
   .INIT(64'ha7c148dba7c148db)  
) LUT6_inst8640 (
   .O(to_level3[864]),
   .I0(level4_in[5184]),
   .I1(level4_in[5185]),
   .I2(level4_in[5186]),
   .I3(level4_in[5187]),
   .I4(level4_in[5188]),
   .I5(level4_in[5189])
);

LUT6 #(
   .INIT(64'h0161710501617105)  
) LUT6_inst8641 (
   .O(to_level3[865]),
   .I0(level4_in[5190]),
   .I1(level4_in[5191]),
   .I2(level4_in[5192]),
   .I3(level4_in[5193]),
   .I4(level4_in[5194]),
   .I5(level4_in[5195])
);

LUT6 #(
   .INIT(64'hfea53226fea53226)  
) LUT6_inst8642 (
   .O(to_level3[866]),
   .I0(level4_in[5196]),
   .I1(level4_in[5197]),
   .I2(level4_in[5198]),
   .I3(level4_in[5199]),
   .I4(level4_in[5200]),
   .I5(level4_in[5201])
);

LUT6 #(
   .INIT(64'h80a0e45a80a0e45a)  
) LUT6_inst8643 (
   .O(to_level3[867]),
   .I0(level4_in[5202]),
   .I1(level4_in[5203]),
   .I2(level4_in[5204]),
   .I3(level4_in[5205]),
   .I4(level4_in[5206]),
   .I5(level4_in[5207])
);

LUT6 #(
   .INIT(64'hba1a9784ba1a9784)  
) LUT6_inst8644 (
   .O(to_level3[868]),
   .I0(level4_in[5208]),
   .I1(level4_in[5209]),
   .I2(level4_in[5210]),
   .I3(level4_in[5211]),
   .I4(level4_in[5212]),
   .I5(level4_in[5213])
);

LUT6 #(
   .INIT(64'haea613bbaea613bb)  
) LUT6_inst8645 (
   .O(to_level3[869]),
   .I0(level4_in[5214]),
   .I1(level4_in[5215]),
   .I2(level4_in[5216]),
   .I3(level4_in[5217]),
   .I4(level4_in[5218]),
   .I5(level4_in[5219])
);

LUT6 #(
   .INIT(64'h791cb2ee791cb2ee)  
) LUT6_inst8646 (
   .O(to_level3[870]),
   .I0(level4_in[5220]),
   .I1(level4_in[5221]),
   .I2(level4_in[5222]),
   .I3(level4_in[5223]),
   .I4(level4_in[5224]),
   .I5(level4_in[5225])
);

LUT6 #(
   .INIT(64'hdaf479bedaf479be)  
) LUT6_inst8647 (
   .O(to_level3[871]),
   .I0(level4_in[5226]),
   .I1(level4_in[5227]),
   .I2(level4_in[5228]),
   .I3(level4_in[5229]),
   .I4(level4_in[5230]),
   .I5(level4_in[5231])
);

LUT6 #(
   .INIT(64'hfe48f98afe48f98a)  
) LUT6_inst8648 (
   .O(to_level3[872]),
   .I0(level4_in[5232]),
   .I1(level4_in[5233]),
   .I2(level4_in[5234]),
   .I3(level4_in[5235]),
   .I4(level4_in[5236]),
   .I5(level4_in[5237])
);

LUT6 #(
   .INIT(64'h6ffbc7646ffbc764)  
) LUT6_inst8649 (
   .O(to_level3[873]),
   .I0(level4_in[5238]),
   .I1(level4_in[5239]),
   .I2(level4_in[5240]),
   .I3(level4_in[5241]),
   .I4(level4_in[5242]),
   .I5(level4_in[5243])
);

LUT6 #(
   .INIT(64'h40162f6240162f62)  
) LUT6_inst8650 (
   .O(to_level3[874]),
   .I0(level4_in[5244]),
   .I1(level4_in[5245]),
   .I2(level4_in[5246]),
   .I3(level4_in[5247]),
   .I4(level4_in[5248]),
   .I5(level4_in[5249])
);

LUT6 #(
   .INIT(64'h7fa217817fa21781)  
) LUT6_inst8651 (
   .O(to_level3[875]),
   .I0(level4_in[5250]),
   .I1(level4_in[5251]),
   .I2(level4_in[5252]),
   .I3(level4_in[5253]),
   .I4(level4_in[5254]),
   .I5(level4_in[5255])
);

LUT6 #(
   .INIT(64'hedc654e1edc654e1)  
) LUT6_inst8652 (
   .O(to_level3[876]),
   .I0(level4_in[5256]),
   .I1(level4_in[5257]),
   .I2(level4_in[5258]),
   .I3(level4_in[5259]),
   .I4(level4_in[5260]),
   .I5(level4_in[5261])
);

LUT6 #(
   .INIT(64'h2d050d752d050d75)  
) LUT6_inst8653 (
   .O(to_level3[877]),
   .I0(level4_in[5262]),
   .I1(level4_in[5263]),
   .I2(level4_in[5264]),
   .I3(level4_in[5265]),
   .I4(level4_in[5266]),
   .I5(level4_in[5267])
);

LUT6 #(
   .INIT(64'hfea4977bfea4977b)  
) LUT6_inst8654 (
   .O(to_level3[878]),
   .I0(level4_in[5268]),
   .I1(level4_in[5269]),
   .I2(level4_in[5270]),
   .I3(level4_in[5271]),
   .I4(level4_in[5272]),
   .I5(level4_in[5273])
);

LUT6 #(
   .INIT(64'hc44aec89c44aec89)  
) LUT6_inst8655 (
   .O(to_level3[879]),
   .I0(level4_in[5274]),
   .I1(level4_in[5275]),
   .I2(level4_in[5276]),
   .I3(level4_in[5277]),
   .I4(level4_in[5278]),
   .I5(level4_in[5279])
);

LUT6 #(
   .INIT(64'h15392b4915392b49)  
) LUT6_inst8656 (
   .O(to_level3[880]),
   .I0(level4_in[5280]),
   .I1(level4_in[5281]),
   .I2(level4_in[5282]),
   .I3(level4_in[5283]),
   .I4(level4_in[5284]),
   .I5(level4_in[5285])
);

LUT6 #(
   .INIT(64'hd5a0a2e3d5a0a2e3)  
) LUT6_inst8657 (
   .O(to_level3[881]),
   .I0(level4_in[5286]),
   .I1(level4_in[5287]),
   .I2(level4_in[5288]),
   .I3(level4_in[5289]),
   .I4(level4_in[5290]),
   .I5(level4_in[5291])
);

LUT6 #(
   .INIT(64'he32ea3a3e32ea3a3)  
) LUT6_inst8658 (
   .O(to_level3[882]),
   .I0(level4_in[5292]),
   .I1(level4_in[5293]),
   .I2(level4_in[5294]),
   .I3(level4_in[5295]),
   .I4(level4_in[5296]),
   .I5(level4_in[5297])
);

LUT6 #(
   .INIT(64'h1ec642f91ec642f9)  
) LUT6_inst8659 (
   .O(to_level3[883]),
   .I0(level4_in[5298]),
   .I1(level4_in[5299]),
   .I2(level4_in[5300]),
   .I3(level4_in[5301]),
   .I4(level4_in[5302]),
   .I5(level4_in[5303])
);

LUT6 #(
   .INIT(64'hd87e1d07d87e1d07)  
) LUT6_inst8660 (
   .O(to_level3[884]),
   .I0(level4_in[5304]),
   .I1(level4_in[5305]),
   .I2(level4_in[5306]),
   .I3(level4_in[5307]),
   .I4(level4_in[5308]),
   .I5(level4_in[5309])
);

LUT6 #(
   .INIT(64'h08c3de4208c3de42)  
) LUT6_inst8661 (
   .O(to_level3[885]),
   .I0(level4_in[5310]),
   .I1(level4_in[5311]),
   .I2(level4_in[5312]),
   .I3(level4_in[5313]),
   .I4(level4_in[5314]),
   .I5(level4_in[5315])
);

LUT6 #(
   .INIT(64'h64c7392664c73926)  
) LUT6_inst8662 (
   .O(to_level3[886]),
   .I0(level4_in[5316]),
   .I1(level4_in[5317]),
   .I2(level4_in[5318]),
   .I3(level4_in[5319]),
   .I4(level4_in[5320]),
   .I5(level4_in[5321])
);

LUT6 #(
   .INIT(64'h9b4650d79b4650d7)  
) LUT6_inst8663 (
   .O(to_level3[887]),
   .I0(level4_in[5322]),
   .I1(level4_in[5323]),
   .I2(level4_in[5324]),
   .I3(level4_in[5325]),
   .I4(level4_in[5326]),
   .I5(level4_in[5327])
);

LUT6 #(
   .INIT(64'h6d6c663d6d6c663d)  
) LUT6_inst8664 (
   .O(to_level3[888]),
   .I0(level4_in[5328]),
   .I1(level4_in[5329]),
   .I2(level4_in[5330]),
   .I3(level4_in[5331]),
   .I4(level4_in[5332]),
   .I5(level4_in[5333])
);

LUT6 #(
   .INIT(64'h7c9b46f87c9b46f8)  
) LUT6_inst8665 (
   .O(to_level3[889]),
   .I0(level4_in[5334]),
   .I1(level4_in[5335]),
   .I2(level4_in[5336]),
   .I3(level4_in[5337]),
   .I4(level4_in[5338]),
   .I5(level4_in[5339])
);

LUT6 #(
   .INIT(64'hca48cbdfca48cbdf)  
) LUT6_inst8666 (
   .O(to_level3[890]),
   .I0(level4_in[5340]),
   .I1(level4_in[5341]),
   .I2(level4_in[5342]),
   .I3(level4_in[5343]),
   .I4(level4_in[5344]),
   .I5(level4_in[5345])
);

LUT6 #(
   .INIT(64'h49e66ac949e66ac9)  
) LUT6_inst8667 (
   .O(to_level3[891]),
   .I0(level4_in[5346]),
   .I1(level4_in[5347]),
   .I2(level4_in[5348]),
   .I3(level4_in[5349]),
   .I4(level4_in[5350]),
   .I5(level4_in[5351])
);

LUT6 #(
   .INIT(64'hff309f7fff309f7f)  
) LUT6_inst8668 (
   .O(to_level3[892]),
   .I0(level4_in[5352]),
   .I1(level4_in[5353]),
   .I2(level4_in[5354]),
   .I3(level4_in[5355]),
   .I4(level4_in[5356]),
   .I5(level4_in[5357])
);

LUT6 #(
   .INIT(64'had5e0cfbad5e0cfb)  
) LUT6_inst8669 (
   .O(to_level3[893]),
   .I0(level4_in[5358]),
   .I1(level4_in[5359]),
   .I2(level4_in[5360]),
   .I3(level4_in[5361]),
   .I4(level4_in[5362]),
   .I5(level4_in[5363])
);

LUT6 #(
   .INIT(64'h0324073a0324073a)  
) LUT6_inst8670 (
   .O(to_level3[894]),
   .I0(level4_in[5364]),
   .I1(level4_in[5365]),
   .I2(level4_in[5366]),
   .I3(level4_in[5367]),
   .I4(level4_in[5368]),
   .I5(level4_in[5369])
);

LUT6 #(
   .INIT(64'h3e071e153e071e15)  
) LUT6_inst8671 (
   .O(to_level3[895]),
   .I0(level4_in[5370]),
   .I1(level4_in[5371]),
   .I2(level4_in[5372]),
   .I3(level4_in[5373]),
   .I4(level4_in[5374]),
   .I5(level4_in[5375])
);

LUT6 #(
   .INIT(64'haf21ac21af21ac21)  
) LUT6_inst8672 (
   .O(to_level3[896]),
   .I0(level4_in[5376]),
   .I1(level4_in[5377]),
   .I2(level4_in[5378]),
   .I3(level4_in[5379]),
   .I4(level4_in[5380]),
   .I5(level4_in[5381])
);

LUT6 #(
   .INIT(64'hf86b7dc0f86b7dc0)  
) LUT6_inst8673 (
   .O(to_level3[897]),
   .I0(level4_in[5382]),
   .I1(level4_in[5383]),
   .I2(level4_in[5384]),
   .I3(level4_in[5385]),
   .I4(level4_in[5386]),
   .I5(level4_in[5387])
);

LUT6 #(
   .INIT(64'h5166286451662864)  
) LUT6_inst8674 (
   .O(to_level3[898]),
   .I0(level4_in[5388]),
   .I1(level4_in[5389]),
   .I2(level4_in[5390]),
   .I3(level4_in[5391]),
   .I4(level4_in[5392]),
   .I5(level4_in[5393])
);

LUT6 #(
   .INIT(64'h4335baa14335baa1)  
) LUT6_inst8675 (
   .O(to_level3[899]),
   .I0(level4_in[5394]),
   .I1(level4_in[5395]),
   .I2(level4_in[5396]),
   .I3(level4_in[5397]),
   .I4(level4_in[5398]),
   .I5(level4_in[5399])
);

LUT6 #(
   .INIT(64'h7fafff397fafff39)  
) LUT6_inst8676 (
   .O(to_level3[900]),
   .I0(level4_in[5400]),
   .I1(level4_in[5401]),
   .I2(level4_in[5402]),
   .I3(level4_in[5403]),
   .I4(level4_in[5404]),
   .I5(level4_in[5405])
);

LUT6 #(
   .INIT(64'hd28a95b0d28a95b0)  
) LUT6_inst8677 (
   .O(to_level3[901]),
   .I0(level4_in[5406]),
   .I1(level4_in[5407]),
   .I2(level4_in[5408]),
   .I3(level4_in[5409]),
   .I4(level4_in[5410]),
   .I5(level4_in[5411])
);

LUT6 #(
   .INIT(64'h8a01d82a8a01d82a)  
) LUT6_inst8678 (
   .O(to_level3[902]),
   .I0(level4_in[5412]),
   .I1(level4_in[5413]),
   .I2(level4_in[5414]),
   .I3(level4_in[5415]),
   .I4(level4_in[5416]),
   .I5(level4_in[5417])
);

LUT6 #(
   .INIT(64'h3614c6253614c625)  
) LUT6_inst8679 (
   .O(to_level3[903]),
   .I0(level4_in[5418]),
   .I1(level4_in[5419]),
   .I2(level4_in[5420]),
   .I3(level4_in[5421]),
   .I4(level4_in[5422]),
   .I5(level4_in[5423])
);

LUT6 #(
   .INIT(64'h3b41564c3b41564c)  
) LUT6_inst8680 (
   .O(to_level3[904]),
   .I0(level4_in[5424]),
   .I1(level4_in[5425]),
   .I2(level4_in[5426]),
   .I3(level4_in[5427]),
   .I4(level4_in[5428]),
   .I5(level4_in[5429])
);

LUT6 #(
   .INIT(64'h715b8ac1715b8ac1)  
) LUT6_inst8681 (
   .O(to_level3[905]),
   .I0(level4_in[5430]),
   .I1(level4_in[5431]),
   .I2(level4_in[5432]),
   .I3(level4_in[5433]),
   .I4(level4_in[5434]),
   .I5(level4_in[5435])
);

LUT6 #(
   .INIT(64'h8a11e80a8a11e80a)  
) LUT6_inst8682 (
   .O(to_level3[906]),
   .I0(level4_in[5436]),
   .I1(level4_in[5437]),
   .I2(level4_in[5438]),
   .I3(level4_in[5439]),
   .I4(level4_in[5440]),
   .I5(level4_in[5441])
);

LUT6 #(
   .INIT(64'hb98048d9b98048d9)  
) LUT6_inst8683 (
   .O(to_level3[907]),
   .I0(level4_in[5442]),
   .I1(level4_in[5443]),
   .I2(level4_in[5444]),
   .I3(level4_in[5445]),
   .I4(level4_in[5446]),
   .I5(level4_in[5447])
);

LUT6 #(
   .INIT(64'hded8fcafded8fcaf)  
) LUT6_inst8684 (
   .O(to_level3[908]),
   .I0(level4_in[5448]),
   .I1(level4_in[5449]),
   .I2(level4_in[5450]),
   .I3(level4_in[5451]),
   .I4(level4_in[5452]),
   .I5(level4_in[5453])
);

LUT6 #(
   .INIT(64'h04c5106c04c5106c)  
) LUT6_inst8685 (
   .O(to_level3[909]),
   .I0(level4_in[5454]),
   .I1(level4_in[5455]),
   .I2(level4_in[5456]),
   .I3(level4_in[5457]),
   .I4(level4_in[5458]),
   .I5(level4_in[5459])
);

LUT6 #(
   .INIT(64'h000ceb21000ceb21)  
) LUT6_inst8686 (
   .O(to_level3[910]),
   .I0(level4_in[5460]),
   .I1(level4_in[5461]),
   .I2(level4_in[5462]),
   .I3(level4_in[5463]),
   .I4(level4_in[5464]),
   .I5(level4_in[5465])
);

LUT6 #(
   .INIT(64'h737c9184737c9184)  
) LUT6_inst8687 (
   .O(to_level3[911]),
   .I0(level4_in[5466]),
   .I1(level4_in[5467]),
   .I2(level4_in[5468]),
   .I3(level4_in[5469]),
   .I4(level4_in[5470]),
   .I5(level4_in[5471])
);

LUT6 #(
   .INIT(64'hea2c7659ea2c7659)  
) LUT6_inst8688 (
   .O(to_level3[912]),
   .I0(level4_in[5472]),
   .I1(level4_in[5473]),
   .I2(level4_in[5474]),
   .I3(level4_in[5475]),
   .I4(level4_in[5476]),
   .I5(level4_in[5477])
);

LUT6 #(
   .INIT(64'h8aeb36098aeb3609)  
) LUT6_inst8689 (
   .O(to_level3[913]),
   .I0(level4_in[5478]),
   .I1(level4_in[5479]),
   .I2(level4_in[5480]),
   .I3(level4_in[5481]),
   .I4(level4_in[5482]),
   .I5(level4_in[5483])
);

LUT6 #(
   .INIT(64'hc03d9d3ec03d9d3e)  
) LUT6_inst8690 (
   .O(to_level3[914]),
   .I0(level4_in[5484]),
   .I1(level4_in[5485]),
   .I2(level4_in[5486]),
   .I3(level4_in[5487]),
   .I4(level4_in[5488]),
   .I5(level4_in[5489])
);

LUT6 #(
   .INIT(64'hfe0860e0fe0860e0)  
) LUT6_inst8691 (
   .O(to_level3[915]),
   .I0(level4_in[5490]),
   .I1(level4_in[5491]),
   .I2(level4_in[5492]),
   .I3(level4_in[5493]),
   .I4(level4_in[5494]),
   .I5(level4_in[5495])
);

LUT6 #(
   .INIT(64'h275fd9e1275fd9e1)  
) LUT6_inst8692 (
   .O(to_level3[916]),
   .I0(level4_in[5496]),
   .I1(level4_in[5497]),
   .I2(level4_in[5498]),
   .I3(level4_in[5499]),
   .I4(level4_in[5500]),
   .I5(level4_in[5501])
);

LUT6 #(
   .INIT(64'h0a048b610a048b61)  
) LUT6_inst8693 (
   .O(to_level3[917]),
   .I0(level4_in[5502]),
   .I1(level4_in[5503]),
   .I2(level4_in[5504]),
   .I3(level4_in[5505]),
   .I4(level4_in[5506]),
   .I5(level4_in[5507])
);

LUT6 #(
   .INIT(64'h535a38b1535a38b1)  
) LUT6_inst8694 (
   .O(to_level3[918]),
   .I0(level4_in[5508]),
   .I1(level4_in[5509]),
   .I2(level4_in[5510]),
   .I3(level4_in[5511]),
   .I4(level4_in[5512]),
   .I5(level4_in[5513])
);

LUT6 #(
   .INIT(64'hac971f15ac971f15)  
) LUT6_inst8695 (
   .O(to_level3[919]),
   .I0(level4_in[5514]),
   .I1(level4_in[5515]),
   .I2(level4_in[5516]),
   .I3(level4_in[5517]),
   .I4(level4_in[5518]),
   .I5(level4_in[5519])
);

LUT6 #(
   .INIT(64'h0e9a859d0e9a859d)  
) LUT6_inst8696 (
   .O(to_level3[920]),
   .I0(level4_in[5520]),
   .I1(level4_in[5521]),
   .I2(level4_in[5522]),
   .I3(level4_in[5523]),
   .I4(level4_in[5524]),
   .I5(level4_in[5525])
);

LUT6 #(
   .INIT(64'h6d54d51d6d54d51d)  
) LUT6_inst8697 (
   .O(to_level3[921]),
   .I0(level4_in[5526]),
   .I1(level4_in[5527]),
   .I2(level4_in[5528]),
   .I3(level4_in[5529]),
   .I4(level4_in[5530]),
   .I5(level4_in[5531])
);

LUT6 #(
   .INIT(64'h153253c8153253c8)  
) LUT6_inst8698 (
   .O(to_level3[922]),
   .I0(level4_in[5532]),
   .I1(level4_in[5533]),
   .I2(level4_in[5534]),
   .I3(level4_in[5535]),
   .I4(level4_in[5536]),
   .I5(level4_in[5537])
);

LUT6 #(
   .INIT(64'hcf99160ecf99160e)  
) LUT6_inst8699 (
   .O(to_level3[923]),
   .I0(level4_in[5538]),
   .I1(level4_in[5539]),
   .I2(level4_in[5540]),
   .I3(level4_in[5541]),
   .I4(level4_in[5542]),
   .I5(level4_in[5543])
);

LUT6 #(
   .INIT(64'hf04f4657f04f4657)  
) LUT6_inst8700 (
   .O(to_level3[924]),
   .I0(level4_in[5544]),
   .I1(level4_in[5545]),
   .I2(level4_in[5546]),
   .I3(level4_in[5547]),
   .I4(level4_in[5548]),
   .I5(level4_in[5549])
);

LUT6 #(
   .INIT(64'h52948c5852948c58)  
) LUT6_inst8701 (
   .O(to_level3[925]),
   .I0(level4_in[5550]),
   .I1(level4_in[5551]),
   .I2(level4_in[5552]),
   .I3(level4_in[5553]),
   .I4(level4_in[5554]),
   .I5(level4_in[5555])
);

LUT6 #(
   .INIT(64'h8acb0f158acb0f15)  
) LUT6_inst8702 (
   .O(to_level3[926]),
   .I0(level4_in[5556]),
   .I1(level4_in[5557]),
   .I2(level4_in[5558]),
   .I3(level4_in[5559]),
   .I4(level4_in[5560]),
   .I5(level4_in[5561])
);

LUT6 #(
   .INIT(64'ha1937844a1937844)  
) LUT6_inst8703 (
   .O(to_level3[927]),
   .I0(level4_in[5562]),
   .I1(level4_in[5563]),
   .I2(level4_in[5564]),
   .I3(level4_in[5565]),
   .I4(level4_in[5566]),
   .I5(level4_in[5567])
);

LUT6 #(
   .INIT(64'h5feb75b55feb75b5)  
) LUT6_inst8704 (
   .O(to_level3[928]),
   .I0(level4_in[5568]),
   .I1(level4_in[5569]),
   .I2(level4_in[5570]),
   .I3(level4_in[5571]),
   .I4(level4_in[5572]),
   .I5(level4_in[5573])
);

LUT6 #(
   .INIT(64'h8b48210b8b48210b)  
) LUT6_inst8705 (
   .O(to_level3[929]),
   .I0(level4_in[5574]),
   .I1(level4_in[5575]),
   .I2(level4_in[5576]),
   .I3(level4_in[5577]),
   .I4(level4_in[5578]),
   .I5(level4_in[5579])
);

LUT6 #(
   .INIT(64'hd614bd07d614bd07)  
) LUT6_inst8706 (
   .O(to_level3[930]),
   .I0(level4_in[5580]),
   .I1(level4_in[5581]),
   .I2(level4_in[5582]),
   .I3(level4_in[5583]),
   .I4(level4_in[5584]),
   .I5(level4_in[5585])
);

LUT6 #(
   .INIT(64'h5f66a6f25f66a6f2)  
) LUT6_inst8707 (
   .O(to_level3[931]),
   .I0(level4_in[5586]),
   .I1(level4_in[5587]),
   .I2(level4_in[5588]),
   .I3(level4_in[5589]),
   .I4(level4_in[5590]),
   .I5(level4_in[5591])
);

LUT6 #(
   .INIT(64'h553e97f2553e97f2)  
) LUT6_inst8708 (
   .O(to_level3[932]),
   .I0(level4_in[5592]),
   .I1(level4_in[5593]),
   .I2(level4_in[5594]),
   .I3(level4_in[5595]),
   .I4(level4_in[5596]),
   .I5(level4_in[5597])
);

LUT6 #(
   .INIT(64'hb15b03a2b15b03a2)  
) LUT6_inst8709 (
   .O(to_level3[933]),
   .I0(level4_in[5598]),
   .I1(level4_in[5599]),
   .I2(level4_in[5600]),
   .I3(level4_in[5601]),
   .I4(level4_in[5602]),
   .I5(level4_in[5603])
);

LUT6 #(
   .INIT(64'h447537cf447537cf)  
) LUT6_inst8710 (
   .O(to_level3[934]),
   .I0(level4_in[5604]),
   .I1(level4_in[5605]),
   .I2(level4_in[5606]),
   .I3(level4_in[5607]),
   .I4(level4_in[5608]),
   .I5(level4_in[5609])
);

LUT6 #(
   .INIT(64'hfaf87d04faf87d04)  
) LUT6_inst8711 (
   .O(to_level3[935]),
   .I0(level4_in[5610]),
   .I1(level4_in[5611]),
   .I2(level4_in[5612]),
   .I3(level4_in[5613]),
   .I4(level4_in[5614]),
   .I5(level4_in[5615])
);

LUT6 #(
   .INIT(64'h3ff6be053ff6be05)  
) LUT6_inst8712 (
   .O(to_level3[936]),
   .I0(level4_in[5616]),
   .I1(level4_in[5617]),
   .I2(level4_in[5618]),
   .I3(level4_in[5619]),
   .I4(level4_in[5620]),
   .I5(level4_in[5621])
);

LUT6 #(
   .INIT(64'h3fd07c693fd07c69)  
) LUT6_inst8713 (
   .O(to_level3[937]),
   .I0(level4_in[5622]),
   .I1(level4_in[5623]),
   .I2(level4_in[5624]),
   .I3(level4_in[5625]),
   .I4(level4_in[5626]),
   .I5(level4_in[5627])
);

LUT6 #(
   .INIT(64'hf45dd6f0f45dd6f0)  
) LUT6_inst8714 (
   .O(to_level3[938]),
   .I0(level4_in[5628]),
   .I1(level4_in[5629]),
   .I2(level4_in[5630]),
   .I3(level4_in[5631]),
   .I4(level4_in[5632]),
   .I5(level4_in[5633])
);

LUT6 #(
   .INIT(64'h695a05d5695a05d5)  
) LUT6_inst8715 (
   .O(to_level3[939]),
   .I0(level4_in[5634]),
   .I1(level4_in[5635]),
   .I2(level4_in[5636]),
   .I3(level4_in[5637]),
   .I4(level4_in[5638]),
   .I5(level4_in[5639])
);

LUT6 #(
   .INIT(64'hed27595bed27595b)  
) LUT6_inst8716 (
   .O(to_level3[940]),
   .I0(level4_in[5640]),
   .I1(level4_in[5641]),
   .I2(level4_in[5642]),
   .I3(level4_in[5643]),
   .I4(level4_in[5644]),
   .I5(level4_in[5645])
);

LUT6 #(
   .INIT(64'h85c4951b85c4951b)  
) LUT6_inst8717 (
   .O(to_level3[941]),
   .I0(level4_in[5646]),
   .I1(level4_in[5647]),
   .I2(level4_in[5648]),
   .I3(level4_in[5649]),
   .I4(level4_in[5650]),
   .I5(level4_in[5651])
);

LUT6 #(
   .INIT(64'he9252ffbe9252ffb)  
) LUT6_inst8718 (
   .O(to_level3[942]),
   .I0(level4_in[5652]),
   .I1(level4_in[5653]),
   .I2(level4_in[5654]),
   .I3(level4_in[5655]),
   .I4(level4_in[5656]),
   .I5(level4_in[5657])
);

LUT6 #(
   .INIT(64'ha7b526b2a7b526b2)  
) LUT6_inst8719 (
   .O(to_level3[943]),
   .I0(level4_in[5658]),
   .I1(level4_in[5659]),
   .I2(level4_in[5660]),
   .I3(level4_in[5661]),
   .I4(level4_in[5662]),
   .I5(level4_in[5663])
);

LUT6 #(
   .INIT(64'h750e433b750e433b)  
) LUT6_inst8720 (
   .O(to_level3[944]),
   .I0(level4_in[5664]),
   .I1(level4_in[5665]),
   .I2(level4_in[5666]),
   .I3(level4_in[5667]),
   .I4(level4_in[5668]),
   .I5(level4_in[5669])
);

LUT6 #(
   .INIT(64'hf99c9134f99c9134)  
) LUT6_inst8721 (
   .O(to_level3[945]),
   .I0(level4_in[5670]),
   .I1(level4_in[5671]),
   .I2(level4_in[5672]),
   .I3(level4_in[5673]),
   .I4(level4_in[5674]),
   .I5(level4_in[5675])
);

LUT6 #(
   .INIT(64'hfbce32c3fbce32c3)  
) LUT6_inst8722 (
   .O(to_level3[946]),
   .I0(level4_in[5676]),
   .I1(level4_in[5677]),
   .I2(level4_in[5678]),
   .I3(level4_in[5679]),
   .I4(level4_in[5680]),
   .I5(level4_in[5681])
);

LUT6 #(
   .INIT(64'h4389b0564389b056)  
) LUT6_inst8723 (
   .O(to_level3[947]),
   .I0(level4_in[5682]),
   .I1(level4_in[5683]),
   .I2(level4_in[5684]),
   .I3(level4_in[5685]),
   .I4(level4_in[5686]),
   .I5(level4_in[5687])
);

LUT6 #(
   .INIT(64'hb3dfd362b3dfd362)  
) LUT6_inst8724 (
   .O(to_level3[948]),
   .I0(level4_in[5688]),
   .I1(level4_in[5689]),
   .I2(level4_in[5690]),
   .I3(level4_in[5691]),
   .I4(level4_in[5692]),
   .I5(level4_in[5693])
);

LUT6 #(
   .INIT(64'hc5c640f2c5c640f2)  
) LUT6_inst8725 (
   .O(to_level3[949]),
   .I0(level4_in[5694]),
   .I1(level4_in[5695]),
   .I2(level4_in[5696]),
   .I3(level4_in[5697]),
   .I4(level4_in[5698]),
   .I5(level4_in[5699])
);

LUT6 #(
   .INIT(64'hf6019e2af6019e2a)  
) LUT6_inst8726 (
   .O(to_level3[950]),
   .I0(level4_in[5700]),
   .I1(level4_in[5701]),
   .I2(level4_in[5702]),
   .I3(level4_in[5703]),
   .I4(level4_in[5704]),
   .I5(level4_in[5705])
);

LUT6 #(
   .INIT(64'h2141344021413440)  
) LUT6_inst8727 (
   .O(to_level3[951]),
   .I0(level4_in[5706]),
   .I1(level4_in[5707]),
   .I2(level4_in[5708]),
   .I3(level4_in[5709]),
   .I4(level4_in[5710]),
   .I5(level4_in[5711])
);

LUT6 #(
   .INIT(64'h64f8ad8a64f8ad8a)  
) LUT6_inst8728 (
   .O(to_level3[952]),
   .I0(level4_in[5712]),
   .I1(level4_in[5713]),
   .I2(level4_in[5714]),
   .I3(level4_in[5715]),
   .I4(level4_in[5716]),
   .I5(level4_in[5717])
);

LUT6 #(
   .INIT(64'hf5d7b112f5d7b112)  
) LUT6_inst8729 (
   .O(to_level3[953]),
   .I0(level4_in[5718]),
   .I1(level4_in[5719]),
   .I2(level4_in[5720]),
   .I3(level4_in[5721]),
   .I4(level4_in[5722]),
   .I5(level4_in[5723])
);

LUT6 #(
   .INIT(64'hbdf21d76bdf21d76)  
) LUT6_inst8730 (
   .O(to_level3[954]),
   .I0(level4_in[5724]),
   .I1(level4_in[5725]),
   .I2(level4_in[5726]),
   .I3(level4_in[5727]),
   .I4(level4_in[5728]),
   .I5(level4_in[5729])
);

LUT6 #(
   .INIT(64'hb8ce7bacb8ce7bac)  
) LUT6_inst8731 (
   .O(to_level3[955]),
   .I0(level4_in[5730]),
   .I1(level4_in[5731]),
   .I2(level4_in[5732]),
   .I3(level4_in[5733]),
   .I4(level4_in[5734]),
   .I5(level4_in[5735])
);

LUT6 #(
   .INIT(64'h3c21d1a03c21d1a0)  
) LUT6_inst8732 (
   .O(to_level3[956]),
   .I0(level4_in[5736]),
   .I1(level4_in[5737]),
   .I2(level4_in[5738]),
   .I3(level4_in[5739]),
   .I4(level4_in[5740]),
   .I5(level4_in[5741])
);

LUT6 #(
   .INIT(64'hbeae8c02beae8c02)  
) LUT6_inst8733 (
   .O(to_level3[957]),
   .I0(level4_in[5742]),
   .I1(level4_in[5743]),
   .I2(level4_in[5744]),
   .I3(level4_in[5745]),
   .I4(level4_in[5746]),
   .I5(level4_in[5747])
);

LUT6 #(
   .INIT(64'hc4c9f598c4c9f598)  
) LUT6_inst8734 (
   .O(to_level3[958]),
   .I0(level4_in[5748]),
   .I1(level4_in[5749]),
   .I2(level4_in[5750]),
   .I3(level4_in[5751]),
   .I4(level4_in[5752]),
   .I5(level4_in[5753])
);

LUT6 #(
   .INIT(64'h86dbce3a86dbce3a)  
) LUT6_inst8735 (
   .O(to_level3[959]),
   .I0(level4_in[5754]),
   .I1(level4_in[5755]),
   .I2(level4_in[5756]),
   .I3(level4_in[5757]),
   .I4(level4_in[5758]),
   .I5(level4_in[5759])
);

LUT6 #(
   .INIT(64'hc427dcb0c427dcb0)  
) LUT6_inst8736 (
   .O(to_level3[960]),
   .I0(level4_in[5760]),
   .I1(level4_in[5761]),
   .I2(level4_in[5762]),
   .I3(level4_in[5763]),
   .I4(level4_in[5764]),
   .I5(level4_in[5765])
);

LUT6 #(
   .INIT(64'hd411b8f0d411b8f0)  
) LUT6_inst8737 (
   .O(to_level3[961]),
   .I0(level4_in[5766]),
   .I1(level4_in[5767]),
   .I2(level4_in[5768]),
   .I3(level4_in[5769]),
   .I4(level4_in[5770]),
   .I5(level4_in[5771])
);

LUT6 #(
   .INIT(64'ha6daf957a6daf957)  
) LUT6_inst8738 (
   .O(to_level3[962]),
   .I0(level4_in[5772]),
   .I1(level4_in[5773]),
   .I2(level4_in[5774]),
   .I3(level4_in[5775]),
   .I4(level4_in[5776]),
   .I5(level4_in[5777])
);

LUT6 #(
   .INIT(64'hec6bc268ec6bc268)  
) LUT6_inst8739 (
   .O(to_level3[963]),
   .I0(level4_in[5778]),
   .I1(level4_in[5779]),
   .I2(level4_in[5780]),
   .I3(level4_in[5781]),
   .I4(level4_in[5782]),
   .I5(level4_in[5783])
);

LUT6 #(
   .INIT(64'h96d2881696d28816)  
) LUT6_inst8740 (
   .O(to_level3[964]),
   .I0(level4_in[5784]),
   .I1(level4_in[5785]),
   .I2(level4_in[5786]),
   .I3(level4_in[5787]),
   .I4(level4_in[5788]),
   .I5(level4_in[5789])
);

LUT6 #(
   .INIT(64'h454086ac454086ac)  
) LUT6_inst8741 (
   .O(to_level3[965]),
   .I0(level4_in[5790]),
   .I1(level4_in[5791]),
   .I2(level4_in[5792]),
   .I3(level4_in[5793]),
   .I4(level4_in[5794]),
   .I5(level4_in[5795])
);

LUT6 #(
   .INIT(64'he0a21ad8e0a21ad8)  
) LUT6_inst8742 (
   .O(to_level3[966]),
   .I0(level4_in[5796]),
   .I1(level4_in[5797]),
   .I2(level4_in[5798]),
   .I3(level4_in[5799]),
   .I4(level4_in[5800]),
   .I5(level4_in[5801])
);

LUT6 #(
   .INIT(64'h3fcb97553fcb9755)  
) LUT6_inst8743 (
   .O(to_level3[967]),
   .I0(level4_in[5802]),
   .I1(level4_in[5803]),
   .I2(level4_in[5804]),
   .I3(level4_in[5805]),
   .I4(level4_in[5806]),
   .I5(level4_in[5807])
);

LUT6 #(
   .INIT(64'h05513bf105513bf1)  
) LUT6_inst8744 (
   .O(to_level3[968]),
   .I0(level4_in[5808]),
   .I1(level4_in[5809]),
   .I2(level4_in[5810]),
   .I3(level4_in[5811]),
   .I4(level4_in[5812]),
   .I5(level4_in[5813])
);

LUT6 #(
   .INIT(64'hb183c785b183c785)  
) LUT6_inst8745 (
   .O(to_level3[969]),
   .I0(level4_in[5814]),
   .I1(level4_in[5815]),
   .I2(level4_in[5816]),
   .I3(level4_in[5817]),
   .I4(level4_in[5818]),
   .I5(level4_in[5819])
);

LUT6 #(
   .INIT(64'hc7d2f33fc7d2f33f)  
) LUT6_inst8746 (
   .O(to_level3[970]),
   .I0(level4_in[5820]),
   .I1(level4_in[5821]),
   .I2(level4_in[5822]),
   .I3(level4_in[5823]),
   .I4(level4_in[5824]),
   .I5(level4_in[5825])
);

LUT6 #(
   .INIT(64'haa2d9ac0aa2d9ac0)  
) LUT6_inst8747 (
   .O(to_level3[971]),
   .I0(level4_in[5826]),
   .I1(level4_in[5827]),
   .I2(level4_in[5828]),
   .I3(level4_in[5829]),
   .I4(level4_in[5830]),
   .I5(level4_in[5831])
);

LUT6 #(
   .INIT(64'h65ed972d65ed972d)  
) LUT6_inst8748 (
   .O(to_level3[972]),
   .I0(level4_in[5832]),
   .I1(level4_in[5833]),
   .I2(level4_in[5834]),
   .I3(level4_in[5835]),
   .I4(level4_in[5836]),
   .I5(level4_in[5837])
);

LUT6 #(
   .INIT(64'hda2bb69ada2bb69a)  
) LUT6_inst8749 (
   .O(to_level3[973]),
   .I0(level4_in[5838]),
   .I1(level4_in[5839]),
   .I2(level4_in[5840]),
   .I3(level4_in[5841]),
   .I4(level4_in[5842]),
   .I5(level4_in[5843])
);

LUT6 #(
   .INIT(64'h93495d0393495d03)  
) LUT6_inst8750 (
   .O(to_level3[974]),
   .I0(level4_in[5844]),
   .I1(level4_in[5845]),
   .I2(level4_in[5846]),
   .I3(level4_in[5847]),
   .I4(level4_in[5848]),
   .I5(level4_in[5849])
);

LUT6 #(
   .INIT(64'h4c2eb52b4c2eb52b)  
) LUT6_inst8751 (
   .O(to_level3[975]),
   .I0(level4_in[5850]),
   .I1(level4_in[5851]),
   .I2(level4_in[5852]),
   .I3(level4_in[5853]),
   .I4(level4_in[5854]),
   .I5(level4_in[5855])
);

LUT6 #(
   .INIT(64'he1e7cb09e1e7cb09)  
) LUT6_inst8752 (
   .O(to_level3[976]),
   .I0(level4_in[5856]),
   .I1(level4_in[5857]),
   .I2(level4_in[5858]),
   .I3(level4_in[5859]),
   .I4(level4_in[5860]),
   .I5(level4_in[5861])
);

LUT6 #(
   .INIT(64'h3cdfdaad3cdfdaad)  
) LUT6_inst8753 (
   .O(to_level3[977]),
   .I0(level4_in[5862]),
   .I1(level4_in[5863]),
   .I2(level4_in[5864]),
   .I3(level4_in[5865]),
   .I4(level4_in[5866]),
   .I5(level4_in[5867])
);

LUT6 #(
   .INIT(64'h8efbad8a8efbad8a)  
) LUT6_inst8754 (
   .O(to_level3[978]),
   .I0(level4_in[5868]),
   .I1(level4_in[5869]),
   .I2(level4_in[5870]),
   .I3(level4_in[5871]),
   .I4(level4_in[5872]),
   .I5(level4_in[5873])
);

LUT6 #(
   .INIT(64'h37553e8537553e85)  
) LUT6_inst8755 (
   .O(to_level3[979]),
   .I0(level4_in[5874]),
   .I1(level4_in[5875]),
   .I2(level4_in[5876]),
   .I3(level4_in[5877]),
   .I4(level4_in[5878]),
   .I5(level4_in[5879])
);

LUT6 #(
   .INIT(64'ha7f843d5a7f843d5)  
) LUT6_inst8756 (
   .O(to_level3[980]),
   .I0(level4_in[5880]),
   .I1(level4_in[5881]),
   .I2(level4_in[5882]),
   .I3(level4_in[5883]),
   .I4(level4_in[5884]),
   .I5(level4_in[5885])
);

LUT6 #(
   .INIT(64'h4222182e4222182e)  
) LUT6_inst8757 (
   .O(to_level3[981]),
   .I0(level4_in[5886]),
   .I1(level4_in[5887]),
   .I2(level4_in[5888]),
   .I3(level4_in[5889]),
   .I4(level4_in[5890]),
   .I5(level4_in[5891])
);

LUT6 #(
   .INIT(64'h89f685ac89f685ac)  
) LUT6_inst8758 (
   .O(to_level3[982]),
   .I0(level4_in[5892]),
   .I1(level4_in[5893]),
   .I2(level4_in[5894]),
   .I3(level4_in[5895]),
   .I4(level4_in[5896]),
   .I5(level4_in[5897])
);

LUT6 #(
   .INIT(64'h347ed981347ed981)  
) LUT6_inst8759 (
   .O(to_level3[983]),
   .I0(level4_in[5898]),
   .I1(level4_in[5899]),
   .I2(level4_in[5900]),
   .I3(level4_in[5901]),
   .I4(level4_in[5902]),
   .I5(level4_in[5903])
);

LUT6 #(
   .INIT(64'ha9b1063ea9b1063e)  
) LUT6_inst8760 (
   .O(to_level3[984]),
   .I0(level4_in[5904]),
   .I1(level4_in[5905]),
   .I2(level4_in[5906]),
   .I3(level4_in[5907]),
   .I4(level4_in[5908]),
   .I5(level4_in[5909])
);

LUT6 #(
   .INIT(64'h7f1e021f7f1e021f)  
) LUT6_inst8761 (
   .O(to_level3[985]),
   .I0(level4_in[5910]),
   .I1(level4_in[5911]),
   .I2(level4_in[5912]),
   .I3(level4_in[5913]),
   .I4(level4_in[5914]),
   .I5(level4_in[5915])
);

LUT6 #(
   .INIT(64'hbb902310bb902310)  
) LUT6_inst8762 (
   .O(to_level3[986]),
   .I0(level4_in[5916]),
   .I1(level4_in[5917]),
   .I2(level4_in[5918]),
   .I3(level4_in[5919]),
   .I4(level4_in[5920]),
   .I5(level4_in[5921])
);

LUT6 #(
   .INIT(64'h4e90a4bf4e90a4bf)  
) LUT6_inst8763 (
   .O(to_level3[987]),
   .I0(level4_in[5922]),
   .I1(level4_in[5923]),
   .I2(level4_in[5924]),
   .I3(level4_in[5925]),
   .I4(level4_in[5926]),
   .I5(level4_in[5927])
);

LUT6 #(
   .INIT(64'hef0e49a6ef0e49a6)  
) LUT6_inst8764 (
   .O(to_level3[988]),
   .I0(level4_in[5928]),
   .I1(level4_in[5929]),
   .I2(level4_in[5930]),
   .I3(level4_in[5931]),
   .I4(level4_in[5932]),
   .I5(level4_in[5933])
);

LUT6 #(
   .INIT(64'hfa944522fa944522)  
) LUT6_inst8765 (
   .O(to_level3[989]),
   .I0(level4_in[5934]),
   .I1(level4_in[5935]),
   .I2(level4_in[5936]),
   .I3(level4_in[5937]),
   .I4(level4_in[5938]),
   .I5(level4_in[5939])
);

LUT6 #(
   .INIT(64'hfc57f1fffc57f1ff)  
) LUT6_inst8766 (
   .O(to_level3[990]),
   .I0(level4_in[5940]),
   .I1(level4_in[5941]),
   .I2(level4_in[5942]),
   .I3(level4_in[5943]),
   .I4(level4_in[5944]),
   .I5(level4_in[5945])
);

LUT6 #(
   .INIT(64'h08c92cf108c92cf1)  
) LUT6_inst8767 (
   .O(to_level3[991]),
   .I0(level4_in[5946]),
   .I1(level4_in[5947]),
   .I2(level4_in[5948]),
   .I3(level4_in[5949]),
   .I4(level4_in[5950]),
   .I5(level4_in[5951])
);

LUT6 #(
   .INIT(64'h3500ec2c3500ec2c)  
) LUT6_inst8768 (
   .O(to_level3[992]),
   .I0(level4_in[5952]),
   .I1(level4_in[5953]),
   .I2(level4_in[5954]),
   .I3(level4_in[5955]),
   .I4(level4_in[5956]),
   .I5(level4_in[5957])
);

LUT6 #(
   .INIT(64'h0ef02bb80ef02bb8)  
) LUT6_inst8769 (
   .O(to_level3[993]),
   .I0(level4_in[5958]),
   .I1(level4_in[5959]),
   .I2(level4_in[5960]),
   .I3(level4_in[5961]),
   .I4(level4_in[5962]),
   .I5(level4_in[5963])
);

LUT6 #(
   .INIT(64'hfac20840fac20840)  
) LUT6_inst8770 (
   .O(to_level3[994]),
   .I0(level4_in[5964]),
   .I1(level4_in[5965]),
   .I2(level4_in[5966]),
   .I3(level4_in[5967]),
   .I4(level4_in[5968]),
   .I5(level4_in[5969])
);

LUT6 #(
   .INIT(64'h2450481c2450481c)  
) LUT6_inst8771 (
   .O(to_level3[995]),
   .I0(level4_in[5970]),
   .I1(level4_in[5971]),
   .I2(level4_in[5972]),
   .I3(level4_in[5973]),
   .I4(level4_in[5974]),
   .I5(level4_in[5975])
);

LUT6 #(
   .INIT(64'h4cc3ee824cc3ee82)  
) LUT6_inst8772 (
   .O(to_level3[996]),
   .I0(level4_in[5976]),
   .I1(level4_in[5977]),
   .I2(level4_in[5978]),
   .I3(level4_in[5979]),
   .I4(level4_in[5980]),
   .I5(level4_in[5981])
);

LUT6 #(
   .INIT(64'hca764ad6ca764ad6)  
) LUT6_inst8773 (
   .O(to_level3[997]),
   .I0(level4_in[5982]),
   .I1(level4_in[5983]),
   .I2(level4_in[5984]),
   .I3(level4_in[5985]),
   .I4(level4_in[5986]),
   .I5(level4_in[5987])
);

LUT6 #(
   .INIT(64'h79a19a8d79a19a8d)  
) LUT6_inst8774 (
   .O(to_level3[998]),
   .I0(level4_in[5988]),
   .I1(level4_in[5989]),
   .I2(level4_in[5990]),
   .I3(level4_in[5991]),
   .I4(level4_in[5992]),
   .I5(level4_in[5993])
);

LUT6 #(
   .INIT(64'h2f954e512f954e51)  
) LUT6_inst8775 (
   .O(to_level3[999]),
   .I0(level4_in[5994]),
   .I1(level4_in[5995]),
   .I2(level4_in[5996]),
   .I3(level4_in[5997]),
   .I4(level4_in[5998]),
   .I5(level4_in[5999])
);

LUT6 #(
   .INIT(64'hd7abe728d7abe728)  
) LUT6_inst8776 (
   .O(to_level3[1000]),
   .I0(level4_in[6000]),
   .I1(level4_in[6001]),
   .I2(level4_in[6002]),
   .I3(level4_in[6003]),
   .I4(level4_in[6004]),
   .I5(level4_in[6005])
);

LUT6 #(
   .INIT(64'h2190953e2190953e)  
) LUT6_inst8777 (
   .O(to_level3[1001]),
   .I0(level4_in[6006]),
   .I1(level4_in[6007]),
   .I2(level4_in[6008]),
   .I3(level4_in[6009]),
   .I4(level4_in[6010]),
   .I5(level4_in[6011])
);

LUT6 #(
   .INIT(64'h1fdc68f01fdc68f0)  
) LUT6_inst8778 (
   .O(to_level3[1002]),
   .I0(level4_in[6012]),
   .I1(level4_in[6013]),
   .I2(level4_in[6014]),
   .I3(level4_in[6015]),
   .I4(level4_in[6016]),
   .I5(level4_in[6017])
);

LUT6 #(
   .INIT(64'h8530fec48530fec4)  
) LUT6_inst8779 (
   .O(to_level3[1003]),
   .I0(level4_in[6018]),
   .I1(level4_in[6019]),
   .I2(level4_in[6020]),
   .I3(level4_in[6021]),
   .I4(level4_in[6022]),
   .I5(level4_in[6023])
);

LUT6 #(
   .INIT(64'h5134c0115134c011)  
) LUT6_inst8780 (
   .O(to_level3[1004]),
   .I0(level4_in[6024]),
   .I1(level4_in[6025]),
   .I2(level4_in[6026]),
   .I3(level4_in[6027]),
   .I4(level4_in[6028]),
   .I5(level4_in[6029])
);

LUT6 #(
   .INIT(64'h1d139d151d139d15)  
) LUT6_inst8781 (
   .O(to_level3[1005]),
   .I0(level4_in[6030]),
   .I1(level4_in[6031]),
   .I2(level4_in[6032]),
   .I3(level4_in[6033]),
   .I4(level4_in[6034]),
   .I5(level4_in[6035])
);

LUT6 #(
   .INIT(64'h4783ae724783ae72)  
) LUT6_inst8782 (
   .O(to_level3[1006]),
   .I0(level4_in[6036]),
   .I1(level4_in[6037]),
   .I2(level4_in[6038]),
   .I3(level4_in[6039]),
   .I4(level4_in[6040]),
   .I5(level4_in[6041])
);

LUT6 #(
   .INIT(64'ha9e2670ba9e2670b)  
) LUT6_inst8783 (
   .O(to_level3[1007]),
   .I0(level4_in[6042]),
   .I1(level4_in[6043]),
   .I2(level4_in[6044]),
   .I3(level4_in[6045]),
   .I4(level4_in[6046]),
   .I5(level4_in[6047])
);

LUT6 #(
   .INIT(64'h4703f9fe4703f9fe)  
) LUT6_inst8784 (
   .O(to_level3[1008]),
   .I0(level4_in[6048]),
   .I1(level4_in[6049]),
   .I2(level4_in[6050]),
   .I3(level4_in[6051]),
   .I4(level4_in[6052]),
   .I5(level4_in[6053])
);

LUT6 #(
   .INIT(64'h6bad1d8f6bad1d8f)  
) LUT6_inst8785 (
   .O(to_level3[1009]),
   .I0(level4_in[6054]),
   .I1(level4_in[6055]),
   .I2(level4_in[6056]),
   .I3(level4_in[6057]),
   .I4(level4_in[6058]),
   .I5(level4_in[6059])
);

LUT6 #(
   .INIT(64'h83e0e68e83e0e68e)  
) LUT6_inst8786 (
   .O(to_level3[1010]),
   .I0(level4_in[6060]),
   .I1(level4_in[6061]),
   .I2(level4_in[6062]),
   .I3(level4_in[6063]),
   .I4(level4_in[6064]),
   .I5(level4_in[6065])
);

LUT6 #(
   .INIT(64'hc3952378c3952378)  
) LUT6_inst8787 (
   .O(to_level3[1011]),
   .I0(level4_in[6066]),
   .I1(level4_in[6067]),
   .I2(level4_in[6068]),
   .I3(level4_in[6069]),
   .I4(level4_in[6070]),
   .I5(level4_in[6071])
);

LUT6 #(
   .INIT(64'h1ce434231ce43423)  
) LUT6_inst8788 (
   .O(to_level3[1012]),
   .I0(level4_in[6072]),
   .I1(level4_in[6073]),
   .I2(level4_in[6074]),
   .I3(level4_in[6075]),
   .I4(level4_in[6076]),
   .I5(level4_in[6077])
);

LUT6 #(
   .INIT(64'hcc534d11cc534d11)  
) LUT6_inst8789 (
   .O(to_level3[1013]),
   .I0(level4_in[6078]),
   .I1(level4_in[6079]),
   .I2(level4_in[6080]),
   .I3(level4_in[6081]),
   .I4(level4_in[6082]),
   .I5(level4_in[6083])
);

LUT6 #(
   .INIT(64'h2643155026431550)  
) LUT6_inst8790 (
   .O(to_level3[1014]),
   .I0(level4_in[6084]),
   .I1(level4_in[6085]),
   .I2(level4_in[6086]),
   .I3(level4_in[6087]),
   .I4(level4_in[6088]),
   .I5(level4_in[6089])
);

LUT6 #(
   .INIT(64'h0f4828020f482802)  
) LUT6_inst8791 (
   .O(to_level3[1015]),
   .I0(level4_in[6090]),
   .I1(level4_in[6091]),
   .I2(level4_in[6092]),
   .I3(level4_in[6093]),
   .I4(level4_in[6094]),
   .I5(level4_in[6095])
);

LUT6 #(
   .INIT(64'hf7df9bc3f7df9bc3)  
) LUT6_inst8792 (
   .O(to_level3[1016]),
   .I0(level4_in[6096]),
   .I1(level4_in[6097]),
   .I2(level4_in[6098]),
   .I3(level4_in[6099]),
   .I4(level4_in[6100]),
   .I5(level4_in[6101])
);

LUT6 #(
   .INIT(64'hd542d430d542d430)  
) LUT6_inst8793 (
   .O(to_level3[1017]),
   .I0(level4_in[6102]),
   .I1(level4_in[6103]),
   .I2(level4_in[6104]),
   .I3(level4_in[6105]),
   .I4(level4_in[6106]),
   .I5(level4_in[6107])
);

LUT6 #(
   .INIT(64'h4a479ec24a479ec2)  
) LUT6_inst8794 (
   .O(to_level3[1018]),
   .I0(level4_in[6108]),
   .I1(level4_in[6109]),
   .I2(level4_in[6110]),
   .I3(level4_in[6111]),
   .I4(level4_in[6112]),
   .I5(level4_in[6113])
);

LUT6 #(
   .INIT(64'h8c28cb5f8c28cb5f)  
) LUT6_inst8795 (
   .O(to_level3[1019]),
   .I0(level4_in[6114]),
   .I1(level4_in[6115]),
   .I2(level4_in[6116]),
   .I3(level4_in[6117]),
   .I4(level4_in[6118]),
   .I5(level4_in[6119])
);

LUT6 #(
   .INIT(64'h22f1d85222f1d852)  
) LUT6_inst8796 (
   .O(to_level3[1020]),
   .I0(level4_in[6120]),
   .I1(level4_in[6121]),
   .I2(level4_in[6122]),
   .I3(level4_in[6123]),
   .I4(level4_in[6124]),
   .I5(level4_in[6125])
);

LUT6 #(
   .INIT(64'h32a2d1c232a2d1c2)  
) LUT6_inst8797 (
   .O(to_level3[1021]),
   .I0(level4_in[6126]),
   .I1(level4_in[6127]),
   .I2(level4_in[6128]),
   .I3(level4_in[6129]),
   .I4(level4_in[6130]),
   .I5(level4_in[6131])
);

LUT6 #(
   .INIT(64'h2c8f3f422c8f3f42)  
) LUT6_inst8798 (
   .O(to_level3[1022]),
   .I0(level4_in[6132]),
   .I1(level4_in[6133]),
   .I2(level4_in[6134]),
   .I3(level4_in[6135]),
   .I4(level4_in[6136]),
   .I5(level4_in[6137])
);

LUT6 #(
   .INIT(64'h40a6bab440a6bab4)  
) LUT6_inst8799 (
   .O(to_level3[1023]),
   .I0(level4_in[6138]),
   .I1(level4_in[6139]),
   .I2(level4_in[6140]),
   .I3(level4_in[6141]),
   .I4(level4_in[6142]),
   .I5(level4_in[6143])
);

LUT6 #(
   .INIT(64'haf90cf44af90cf44)  
) LUT6_inst8800 (
   .O(to_level3[1024]),
   .I0(level4_in[6144]),
   .I1(level4_in[6145]),
   .I2(level4_in[6146]),
   .I3(level4_in[6147]),
   .I4(level4_in[6148]),
   .I5(level4_in[6149])
);

LUT6 #(
   .INIT(64'h3200b46e3200b46e)  
) LUT6_inst8801 (
   .O(to_level3[1025]),
   .I0(level4_in[6150]),
   .I1(level4_in[6151]),
   .I2(level4_in[6152]),
   .I3(level4_in[6153]),
   .I4(level4_in[6154]),
   .I5(level4_in[6155])
);

LUT6 #(
   .INIT(64'hcef5031acef5031a)  
) LUT6_inst8802 (
   .O(to_level3[1026]),
   .I0(level4_in[6156]),
   .I1(level4_in[6157]),
   .I2(level4_in[6158]),
   .I3(level4_in[6159]),
   .I4(level4_in[6160]),
   .I5(level4_in[6161])
);

LUT6 #(
   .INIT(64'h133d2218133d2218)  
) LUT6_inst8803 (
   .O(to_level3[1027]),
   .I0(level4_in[6162]),
   .I1(level4_in[6163]),
   .I2(level4_in[6164]),
   .I3(level4_in[6165]),
   .I4(level4_in[6166]),
   .I5(level4_in[6167])
);

LUT6 #(
   .INIT(64'h800de19e800de19e)  
) LUT6_inst8804 (
   .O(to_level3[1028]),
   .I0(level4_in[6168]),
   .I1(level4_in[6169]),
   .I2(level4_in[6170]),
   .I3(level4_in[6171]),
   .I4(level4_in[6172]),
   .I5(level4_in[6173])
);

LUT6 #(
   .INIT(64'h47f4575b47f4575b)  
) LUT6_inst8805 (
   .O(to_level3[1029]),
   .I0(level4_in[6174]),
   .I1(level4_in[6175]),
   .I2(level4_in[6176]),
   .I3(level4_in[6177]),
   .I4(level4_in[6178]),
   .I5(level4_in[6179])
);

LUT6 #(
   .INIT(64'h188dc2fa188dc2fa)  
) LUT6_inst8806 (
   .O(to_level3[1030]),
   .I0(level4_in[6180]),
   .I1(level4_in[6181]),
   .I2(level4_in[6182]),
   .I3(level4_in[6183]),
   .I4(level4_in[6184]),
   .I5(level4_in[6185])
);

LUT6 #(
   .INIT(64'hd491bc02d491bc02)  
) LUT6_inst8807 (
   .O(to_level3[1031]),
   .I0(level4_in[6186]),
   .I1(level4_in[6187]),
   .I2(level4_in[6188]),
   .I3(level4_in[6189]),
   .I4(level4_in[6190]),
   .I5(level4_in[6191])
);

LUT6 #(
   .INIT(64'haffffdd5affffdd5)  
) LUT6_inst8808 (
   .O(to_level3[1032]),
   .I0(level4_in[6192]),
   .I1(level4_in[6193]),
   .I2(level4_in[6194]),
   .I3(level4_in[6195]),
   .I4(level4_in[6196]),
   .I5(level4_in[6197])
);

LUT6 #(
   .INIT(64'h9b2f00909b2f0090)  
) LUT6_inst8809 (
   .O(to_level3[1033]),
   .I0(level4_in[6198]),
   .I1(level4_in[6199]),
   .I2(level4_in[6200]),
   .I3(level4_in[6201]),
   .I4(level4_in[6202]),
   .I5(level4_in[6203])
);

LUT6 #(
   .INIT(64'he374605de374605d)  
) LUT6_inst8810 (
   .O(to_level3[1034]),
   .I0(level4_in[6204]),
   .I1(level4_in[6205]),
   .I2(level4_in[6206]),
   .I3(level4_in[6207]),
   .I4(level4_in[6208]),
   .I5(level4_in[6209])
);

LUT6 #(
   .INIT(64'h349f5ddb349f5ddb)  
) LUT6_inst8811 (
   .O(to_level3[1035]),
   .I0(level4_in[6210]),
   .I1(level4_in[6211]),
   .I2(level4_in[6212]),
   .I3(level4_in[6213]),
   .I4(level4_in[6214]),
   .I5(level4_in[6215])
);

LUT6 #(
   .INIT(64'hda152c5fda152c5f)  
) LUT6_inst8812 (
   .O(to_level3[1036]),
   .I0(level4_in[6216]),
   .I1(level4_in[6217]),
   .I2(level4_in[6218]),
   .I3(level4_in[6219]),
   .I4(level4_in[6220]),
   .I5(level4_in[6221])
);

LUT6 #(
   .INIT(64'h599854a6599854a6)  
) LUT6_inst8813 (
   .O(to_level3[1037]),
   .I0(level4_in[6222]),
   .I1(level4_in[6223]),
   .I2(level4_in[6224]),
   .I3(level4_in[6225]),
   .I4(level4_in[6226]),
   .I5(level4_in[6227])
);

LUT6 #(
   .INIT(64'h110c4e63110c4e63)  
) LUT6_inst8814 (
   .O(to_level3[1038]),
   .I0(level4_in[6228]),
   .I1(level4_in[6229]),
   .I2(level4_in[6230]),
   .I3(level4_in[6231]),
   .I4(level4_in[6232]),
   .I5(level4_in[6233])
);

LUT6 #(
   .INIT(64'hdb2b577adb2b577a)  
) LUT6_inst8815 (
   .O(to_level3[1039]),
   .I0(level4_in[6234]),
   .I1(level4_in[6235]),
   .I2(level4_in[6236]),
   .I3(level4_in[6237]),
   .I4(level4_in[6238]),
   .I5(level4_in[6239])
);

LUT6 #(
   .INIT(64'hd25a1713d25a1713)  
) LUT6_inst8816 (
   .O(to_level3[1040]),
   .I0(level4_in[6240]),
   .I1(level4_in[6241]),
   .I2(level4_in[6242]),
   .I3(level4_in[6243]),
   .I4(level4_in[6244]),
   .I5(level4_in[6245])
);

LUT6 #(
   .INIT(64'h924173c4924173c4)  
) LUT6_inst8817 (
   .O(to_level3[1041]),
   .I0(level4_in[6246]),
   .I1(level4_in[6247]),
   .I2(level4_in[6248]),
   .I3(level4_in[6249]),
   .I4(level4_in[6250]),
   .I5(level4_in[6251])
);

LUT6 #(
   .INIT(64'h34a439ea34a439ea)  
) LUT6_inst8818 (
   .O(to_level3[1042]),
   .I0(level4_in[6252]),
   .I1(level4_in[6253]),
   .I2(level4_in[6254]),
   .I3(level4_in[6255]),
   .I4(level4_in[6256]),
   .I5(level4_in[6257])
);

LUT6 #(
   .INIT(64'h2362995823629958)  
) LUT6_inst8819 (
   .O(to_level3[1043]),
   .I0(level4_in[6258]),
   .I1(level4_in[6259]),
   .I2(level4_in[6260]),
   .I3(level4_in[6261]),
   .I4(level4_in[6262]),
   .I5(level4_in[6263])
);

LUT6 #(
   .INIT(64'h2ecec0a72ecec0a7)  
) LUT6_inst8820 (
   .O(to_level3[1044]),
   .I0(level4_in[6264]),
   .I1(level4_in[6265]),
   .I2(level4_in[6266]),
   .I3(level4_in[6267]),
   .I4(level4_in[6268]),
   .I5(level4_in[6269])
);

LUT6 #(
   .INIT(64'h5c72d9f35c72d9f3)  
) LUT6_inst8821 (
   .O(to_level3[1045]),
   .I0(level4_in[6270]),
   .I1(level4_in[6271]),
   .I2(level4_in[6272]),
   .I3(level4_in[6273]),
   .I4(level4_in[6274]),
   .I5(level4_in[6275])
);

LUT6 #(
   .INIT(64'hd5127b40d5127b40)  
) LUT6_inst8822 (
   .O(to_level3[1046]),
   .I0(level4_in[6276]),
   .I1(level4_in[6277]),
   .I2(level4_in[6278]),
   .I3(level4_in[6279]),
   .I4(level4_in[6280]),
   .I5(level4_in[6281])
);

LUT6 #(
   .INIT(64'hacca4cdfacca4cdf)  
) LUT6_inst8823 (
   .O(to_level3[1047]),
   .I0(level4_in[6282]),
   .I1(level4_in[6283]),
   .I2(level4_in[6284]),
   .I3(level4_in[6285]),
   .I4(level4_in[6286]),
   .I5(level4_in[6287])
);

LUT6 #(
   .INIT(64'h689ba743689ba743)  
) LUT6_inst8824 (
   .O(to_level3[1048]),
   .I0(level4_in[6288]),
   .I1(level4_in[6289]),
   .I2(level4_in[6290]),
   .I3(level4_in[6291]),
   .I4(level4_in[6292]),
   .I5(level4_in[6293])
);

LUT6 #(
   .INIT(64'h617f5fae617f5fae)  
) LUT6_inst8825 (
   .O(to_level3[1049]),
   .I0(level4_in[6294]),
   .I1(level4_in[6295]),
   .I2(level4_in[6296]),
   .I3(level4_in[6297]),
   .I4(level4_in[6298]),
   .I5(level4_in[6299])
);

LUT6 #(
   .INIT(64'h8312999683129996)  
) LUT6_inst8826 (
   .O(to_level3[1050]),
   .I0(level4_in[6300]),
   .I1(level4_in[6301]),
   .I2(level4_in[6302]),
   .I3(level4_in[6303]),
   .I4(level4_in[6304]),
   .I5(level4_in[6305])
);

LUT6 #(
   .INIT(64'hac90e9b7ac90e9b7)  
) LUT6_inst8827 (
   .O(to_level3[1051]),
   .I0(level4_in[6306]),
   .I1(level4_in[6307]),
   .I2(level4_in[6308]),
   .I3(level4_in[6309]),
   .I4(level4_in[6310]),
   .I5(level4_in[6311])
);

LUT6 #(
   .INIT(64'h002389ee002389ee)  
) LUT6_inst8828 (
   .O(to_level3[1052]),
   .I0(level4_in[6312]),
   .I1(level4_in[6313]),
   .I2(level4_in[6314]),
   .I3(level4_in[6315]),
   .I4(level4_in[6316]),
   .I5(level4_in[6317])
);

LUT6 #(
   .INIT(64'h8fe05a1d8fe05a1d)  
) LUT6_inst8829 (
   .O(to_level3[1053]),
   .I0(level4_in[6318]),
   .I1(level4_in[6319]),
   .I2(level4_in[6320]),
   .I3(level4_in[6321]),
   .I4(level4_in[6322]),
   .I5(level4_in[6323])
);

LUT6 #(
   .INIT(64'h8d8cb7ab8d8cb7ab)  
) LUT6_inst8830 (
   .O(to_level3[1054]),
   .I0(level4_in[6324]),
   .I1(level4_in[6325]),
   .I2(level4_in[6326]),
   .I3(level4_in[6327]),
   .I4(level4_in[6328]),
   .I5(level4_in[6329])
);

LUT6 #(
   .INIT(64'h598c939b598c939b)  
) LUT6_inst8831 (
   .O(to_level3[1055]),
   .I0(level4_in[6330]),
   .I1(level4_in[6331]),
   .I2(level4_in[6332]),
   .I3(level4_in[6333]),
   .I4(level4_in[6334]),
   .I5(level4_in[6335])
);

LUT6 #(
   .INIT(64'h4901ae214901ae21)  
) LUT6_inst8832 (
   .O(to_level3[1056]),
   .I0(level4_in[6336]),
   .I1(level4_in[6337]),
   .I2(level4_in[6338]),
   .I3(level4_in[6339]),
   .I4(level4_in[6340]),
   .I5(level4_in[6341])
);

LUT6 #(
   .INIT(64'h8a7a7e1c8a7a7e1c)  
) LUT6_inst8833 (
   .O(to_level3[1057]),
   .I0(level4_in[6342]),
   .I1(level4_in[6343]),
   .I2(level4_in[6344]),
   .I3(level4_in[6345]),
   .I4(level4_in[6346]),
   .I5(level4_in[6347])
);

LUT6 #(
   .INIT(64'h4b9e24d14b9e24d1)  
) LUT6_inst8834 (
   .O(to_level3[1058]),
   .I0(level4_in[6348]),
   .I1(level4_in[6349]),
   .I2(level4_in[6350]),
   .I3(level4_in[6351]),
   .I4(level4_in[6352]),
   .I5(level4_in[6353])
);

LUT6 #(
   .INIT(64'he24dbaa6e24dbaa6)  
) LUT6_inst8835 (
   .O(to_level3[1059]),
   .I0(level4_in[6354]),
   .I1(level4_in[6355]),
   .I2(level4_in[6356]),
   .I3(level4_in[6357]),
   .I4(level4_in[6358]),
   .I5(level4_in[6359])
);

LUT6 #(
   .INIT(64'h7dc99c357dc99c35)  
) LUT6_inst8836 (
   .O(to_level3[1060]),
   .I0(level4_in[6360]),
   .I1(level4_in[6361]),
   .I2(level4_in[6362]),
   .I3(level4_in[6363]),
   .I4(level4_in[6364]),
   .I5(level4_in[6365])
);

LUT6 #(
   .INIT(64'he9e7e745e9e7e745)  
) LUT6_inst8837 (
   .O(to_level3[1061]),
   .I0(level4_in[6366]),
   .I1(level4_in[6367]),
   .I2(level4_in[6368]),
   .I3(level4_in[6369]),
   .I4(level4_in[6370]),
   .I5(level4_in[6371])
);

LUT6 #(
   .INIT(64'he781db38e781db38)  
) LUT6_inst8838 (
   .O(to_level3[1062]),
   .I0(level4_in[6372]),
   .I1(level4_in[6373]),
   .I2(level4_in[6374]),
   .I3(level4_in[6375]),
   .I4(level4_in[6376]),
   .I5(level4_in[6377])
);

LUT6 #(
   .INIT(64'h68ea0ca468ea0ca4)  
) LUT6_inst8839 (
   .O(to_level3[1063]),
   .I0(level4_in[6378]),
   .I1(level4_in[6379]),
   .I2(level4_in[6380]),
   .I3(level4_in[6381]),
   .I4(level4_in[6382]),
   .I5(level4_in[6383])
);

LUT6 #(
   .INIT(64'hc7657502c7657502)  
) LUT6_inst8840 (
   .O(to_level3[1064]),
   .I0(level4_in[6384]),
   .I1(level4_in[6385]),
   .I2(level4_in[6386]),
   .I3(level4_in[6387]),
   .I4(level4_in[6388]),
   .I5(level4_in[6389])
);

LUT6 #(
   .INIT(64'h375b22c5375b22c5)  
) LUT6_inst8841 (
   .O(to_level3[1065]),
   .I0(level4_in[6390]),
   .I1(level4_in[6391]),
   .I2(level4_in[6392]),
   .I3(level4_in[6393]),
   .I4(level4_in[6394]),
   .I5(level4_in[6395])
);

LUT6 #(
   .INIT(64'h8fc3f5718fc3f571)  
) LUT6_inst8842 (
   .O(to_level3[1066]),
   .I0(level4_in[6396]),
   .I1(level4_in[6397]),
   .I2(level4_in[6398]),
   .I3(level4_in[6399]),
   .I4(level4_in[6400]),
   .I5(level4_in[6401])
);

LUT6 #(
   .INIT(64'hc254d14fc254d14f)  
) LUT6_inst8843 (
   .O(to_level3[1067]),
   .I0(level4_in[6402]),
   .I1(level4_in[6403]),
   .I2(level4_in[6404]),
   .I3(level4_in[6405]),
   .I4(level4_in[6406]),
   .I5(level4_in[6407])
);

LUT6 #(
   .INIT(64'h2acbb8032acbb803)  
) LUT6_inst8844 (
   .O(to_level3[1068]),
   .I0(level4_in[6408]),
   .I1(level4_in[6409]),
   .I2(level4_in[6410]),
   .I3(level4_in[6411]),
   .I4(level4_in[6412]),
   .I5(level4_in[6413])
);

LUT6 #(
   .INIT(64'hc6d31676c6d31676)  
) LUT6_inst8845 (
   .O(to_level3[1069]),
   .I0(level4_in[6414]),
   .I1(level4_in[6415]),
   .I2(level4_in[6416]),
   .I3(level4_in[6417]),
   .I4(level4_in[6418]),
   .I5(level4_in[6419])
);

LUT6 #(
   .INIT(64'h19cf36f019cf36f0)  
) LUT6_inst8846 (
   .O(to_level3[1070]),
   .I0(level4_in[6420]),
   .I1(level4_in[6421]),
   .I2(level4_in[6422]),
   .I3(level4_in[6423]),
   .I4(level4_in[6424]),
   .I5(level4_in[6425])
);

LUT6 #(
   .INIT(64'heae2bf84eae2bf84)  
) LUT6_inst8847 (
   .O(to_level3[1071]),
   .I0(level4_in[6426]),
   .I1(level4_in[6427]),
   .I2(level4_in[6428]),
   .I3(level4_in[6429]),
   .I4(level4_in[6430]),
   .I5(level4_in[6431])
);

LUT6 #(
   .INIT(64'h9b273e839b273e83)  
) LUT6_inst8848 (
   .O(to_level3[1072]),
   .I0(level4_in[6432]),
   .I1(level4_in[6433]),
   .I2(level4_in[6434]),
   .I3(level4_in[6435]),
   .I4(level4_in[6436]),
   .I5(level4_in[6437])
);

LUT6 #(
   .INIT(64'h0ac317b50ac317b5)  
) LUT6_inst8849 (
   .O(to_level3[1073]),
   .I0(level4_in[6438]),
   .I1(level4_in[6439]),
   .I2(level4_in[6440]),
   .I3(level4_in[6441]),
   .I4(level4_in[6442]),
   .I5(level4_in[6443])
);

LUT6 #(
   .INIT(64'h9b74afc69b74afc6)  
) LUT6_inst8850 (
   .O(to_level3[1074]),
   .I0(level4_in[6444]),
   .I1(level4_in[6445]),
   .I2(level4_in[6446]),
   .I3(level4_in[6447]),
   .I4(level4_in[6448]),
   .I5(level4_in[6449])
);

LUT6 #(
   .INIT(64'h7ff7ba407ff7ba40)  
) LUT6_inst8851 (
   .O(to_level3[1075]),
   .I0(level4_in[6450]),
   .I1(level4_in[6451]),
   .I2(level4_in[6452]),
   .I3(level4_in[6453]),
   .I4(level4_in[6454]),
   .I5(level4_in[6455])
);

LUT6 #(
   .INIT(64'h05bf214b05bf214b)  
) LUT6_inst8852 (
   .O(to_level3[1076]),
   .I0(level4_in[6456]),
   .I1(level4_in[6457]),
   .I2(level4_in[6458]),
   .I3(level4_in[6459]),
   .I4(level4_in[6460]),
   .I5(level4_in[6461])
);

LUT6 #(
   .INIT(64'h1d9ae5cf1d9ae5cf)  
) LUT6_inst8853 (
   .O(to_level3[1077]),
   .I0(level4_in[6462]),
   .I1(level4_in[6463]),
   .I2(level4_in[6464]),
   .I3(level4_in[6465]),
   .I4(level4_in[6466]),
   .I5(level4_in[6467])
);

LUT6 #(
   .INIT(64'hd38cbfa6d38cbfa6)  
) LUT6_inst8854 (
   .O(to_level3[1078]),
   .I0(level4_in[6468]),
   .I1(level4_in[6469]),
   .I2(level4_in[6470]),
   .I3(level4_in[6471]),
   .I4(level4_in[6472]),
   .I5(level4_in[6473])
);

LUT6 #(
   .INIT(64'h361c4e0f361c4e0f)  
) LUT6_inst8855 (
   .O(to_level3[1079]),
   .I0(level4_in[6474]),
   .I1(level4_in[6475]),
   .I2(level4_in[6476]),
   .I3(level4_in[6477]),
   .I4(level4_in[6478]),
   .I5(level4_in[6479])
);

LUT6 #(
   .INIT(64'h260f33e8260f33e8)  
) LUT6_inst8856 (
   .O(to_level3[1080]),
   .I0(level4_in[6480]),
   .I1(level4_in[6481]),
   .I2(level4_in[6482]),
   .I3(level4_in[6483]),
   .I4(level4_in[6484]),
   .I5(level4_in[6485])
);

LUT6 #(
   .INIT(64'h1cedae731cedae73)  
) LUT6_inst8857 (
   .O(to_level3[1081]),
   .I0(level4_in[6486]),
   .I1(level4_in[6487]),
   .I2(level4_in[6488]),
   .I3(level4_in[6489]),
   .I4(level4_in[6490]),
   .I5(level4_in[6491])
);

LUT6 #(
   .INIT(64'h71294ec571294ec5)  
) LUT6_inst8858 (
   .O(to_level3[1082]),
   .I0(level4_in[6492]),
   .I1(level4_in[6493]),
   .I2(level4_in[6494]),
   .I3(level4_in[6495]),
   .I4(level4_in[6496]),
   .I5(level4_in[6497])
);

LUT6 #(
   .INIT(64'hb6f349e1b6f349e1)  
) LUT6_inst8859 (
   .O(to_level3[1083]),
   .I0(level4_in[6498]),
   .I1(level4_in[6499]),
   .I2(level4_in[6500]),
   .I3(level4_in[6501]),
   .I4(level4_in[6502]),
   .I5(level4_in[6503])
);

LUT6 #(
   .INIT(64'hb1af8584b1af8584)  
) LUT6_inst8860 (
   .O(to_level3[1084]),
   .I0(level4_in[6504]),
   .I1(level4_in[6505]),
   .I2(level4_in[6506]),
   .I3(level4_in[6507]),
   .I4(level4_in[6508]),
   .I5(level4_in[6509])
);

LUT6 #(
   .INIT(64'h1b7aeb2d1b7aeb2d)  
) LUT6_inst8861 (
   .O(to_level3[1085]),
   .I0(level4_in[6510]),
   .I1(level4_in[6511]),
   .I2(level4_in[6512]),
   .I3(level4_in[6513]),
   .I4(level4_in[6514]),
   .I5(level4_in[6515])
);

LUT6 #(
   .INIT(64'h3b76a5363b76a536)  
) LUT6_inst8862 (
   .O(to_level3[1086]),
   .I0(level4_in[6516]),
   .I1(level4_in[6517]),
   .I2(level4_in[6518]),
   .I3(level4_in[6519]),
   .I4(level4_in[6520]),
   .I5(level4_in[6521])
);

LUT6 #(
   .INIT(64'h7d77e1a27d77e1a2)  
) LUT6_inst8863 (
   .O(to_level3[1087]),
   .I0(level4_in[6522]),
   .I1(level4_in[6523]),
   .I2(level4_in[6524]),
   .I3(level4_in[6525]),
   .I4(level4_in[6526]),
   .I5(level4_in[6527])
);

LUT6 #(
   .INIT(64'h3f6d84fd3f6d84fd)  
) LUT6_inst8864 (
   .O(to_level3[1088]),
   .I0(level4_in[6528]),
   .I1(level4_in[6529]),
   .I2(level4_in[6530]),
   .I3(level4_in[6531]),
   .I4(level4_in[6532]),
   .I5(level4_in[6533])
);

LUT6 #(
   .INIT(64'h1058920b1058920b)  
) LUT6_inst8865 (
   .O(to_level3[1089]),
   .I0(level4_in[6534]),
   .I1(level4_in[6535]),
   .I2(level4_in[6536]),
   .I3(level4_in[6537]),
   .I4(level4_in[6538]),
   .I5(level4_in[6539])
);

LUT6 #(
   .INIT(64'h9bc675bd9bc675bd)  
) LUT6_inst8866 (
   .O(to_level3[1090]),
   .I0(level4_in[6540]),
   .I1(level4_in[6541]),
   .I2(level4_in[6542]),
   .I3(level4_in[6543]),
   .I4(level4_in[6544]),
   .I5(level4_in[6545])
);

LUT6 #(
   .INIT(64'hcaaaeac1caaaeac1)  
) LUT6_inst8867 (
   .O(to_level3[1091]),
   .I0(level4_in[6546]),
   .I1(level4_in[6547]),
   .I2(level4_in[6548]),
   .I3(level4_in[6549]),
   .I4(level4_in[6550]),
   .I5(level4_in[6551])
);

LUT6 #(
   .INIT(64'h4c3129a04c3129a0)  
) LUT6_inst8868 (
   .O(to_level3[1092]),
   .I0(level4_in[6552]),
   .I1(level4_in[6553]),
   .I2(level4_in[6554]),
   .I3(level4_in[6555]),
   .I4(level4_in[6556]),
   .I5(level4_in[6557])
);

LUT6 #(
   .INIT(64'hc77605cfc77605cf)  
) LUT6_inst8869 (
   .O(to_level3[1093]),
   .I0(level4_in[6558]),
   .I1(level4_in[6559]),
   .I2(level4_in[6560]),
   .I3(level4_in[6561]),
   .I4(level4_in[6562]),
   .I5(level4_in[6563])
);

LUT6 #(
   .INIT(64'h10b5d06110b5d061)  
) LUT6_inst8870 (
   .O(to_level3[1094]),
   .I0(level4_in[6564]),
   .I1(level4_in[6565]),
   .I2(level4_in[6566]),
   .I3(level4_in[6567]),
   .I4(level4_in[6568]),
   .I5(level4_in[6569])
);

LUT6 #(
   .INIT(64'h0599475e0599475e)  
) LUT6_inst8871 (
   .O(to_level3[1095]),
   .I0(level4_in[6570]),
   .I1(level4_in[6571]),
   .I2(level4_in[6572]),
   .I3(level4_in[6573]),
   .I4(level4_in[6574]),
   .I5(level4_in[6575])
);

LUT6 #(
   .INIT(64'h291a9bd9291a9bd9)  
) LUT6_inst8872 (
   .O(to_level3[1096]),
   .I0(level4_in[6576]),
   .I1(level4_in[6577]),
   .I2(level4_in[6578]),
   .I3(level4_in[6579]),
   .I4(level4_in[6580]),
   .I5(level4_in[6581])
);

LUT6 #(
   .INIT(64'h103e25f5103e25f5)  
) LUT6_inst8873 (
   .O(to_level3[1097]),
   .I0(level4_in[6582]),
   .I1(level4_in[6583]),
   .I2(level4_in[6584]),
   .I3(level4_in[6585]),
   .I4(level4_in[6586]),
   .I5(level4_in[6587])
);

LUT6 #(
   .INIT(64'hfde54066fde54066)  
) LUT6_inst8874 (
   .O(to_level3[1098]),
   .I0(level4_in[6588]),
   .I1(level4_in[6589]),
   .I2(level4_in[6590]),
   .I3(level4_in[6591]),
   .I4(level4_in[6592]),
   .I5(level4_in[6593])
);

LUT6 #(
   .INIT(64'h68a8830968a88309)  
) LUT6_inst8875 (
   .O(to_level3[1099]),
   .I0(level4_in[6594]),
   .I1(level4_in[6595]),
   .I2(level4_in[6596]),
   .I3(level4_in[6597]),
   .I4(level4_in[6598]),
   .I5(level4_in[6599])
);

LUT6 #(
   .INIT(64'h3c60ab463c60ab46)  
) LUT6_inst8876 (
   .O(to_level3[1100]),
   .I0(level4_in[6600]),
   .I1(level4_in[6601]),
   .I2(level4_in[6602]),
   .I3(level4_in[6603]),
   .I4(level4_in[6604]),
   .I5(level4_in[6605])
);

LUT6 #(
   .INIT(64'h8ffefc9f8ffefc9f)  
) LUT6_inst8877 (
   .O(to_level3[1101]),
   .I0(level4_in[6606]),
   .I1(level4_in[6607]),
   .I2(level4_in[6608]),
   .I3(level4_in[6609]),
   .I4(level4_in[6610]),
   .I5(level4_in[6611])
);

LUT6 #(
   .INIT(64'h7a14bf527a14bf52)  
) LUT6_inst8878 (
   .O(to_level3[1102]),
   .I0(level4_in[6612]),
   .I1(level4_in[6613]),
   .I2(level4_in[6614]),
   .I3(level4_in[6615]),
   .I4(level4_in[6616]),
   .I5(level4_in[6617])
);

LUT6 #(
   .INIT(64'h0062896200628962)  
) LUT6_inst8879 (
   .O(to_level3[1103]),
   .I0(level4_in[6618]),
   .I1(level4_in[6619]),
   .I2(level4_in[6620]),
   .I3(level4_in[6621]),
   .I4(level4_in[6622]),
   .I5(level4_in[6623])
);

LUT6 #(
   .INIT(64'hbd756967bd756967)  
) LUT6_inst8880 (
   .O(to_level3[1104]),
   .I0(level4_in[6624]),
   .I1(level4_in[6625]),
   .I2(level4_in[6626]),
   .I3(level4_in[6627]),
   .I4(level4_in[6628]),
   .I5(level4_in[6629])
);

LUT6 #(
   .INIT(64'hbd4f225dbd4f225d)  
) LUT6_inst8881 (
   .O(to_level3[1105]),
   .I0(level4_in[6630]),
   .I1(level4_in[6631]),
   .I2(level4_in[6632]),
   .I3(level4_in[6633]),
   .I4(level4_in[6634]),
   .I5(level4_in[6635])
);

LUT6 #(
   .INIT(64'he258525de258525d)  
) LUT6_inst8882 (
   .O(to_level3[1106]),
   .I0(level4_in[6636]),
   .I1(level4_in[6637]),
   .I2(level4_in[6638]),
   .I3(level4_in[6639]),
   .I4(level4_in[6640]),
   .I5(level4_in[6641])
);

LUT6 #(
   .INIT(64'hd26f9068d26f9068)  
) LUT6_inst8883 (
   .O(to_level3[1107]),
   .I0(level4_in[6642]),
   .I1(level4_in[6643]),
   .I2(level4_in[6644]),
   .I3(level4_in[6645]),
   .I4(level4_in[6646]),
   .I5(level4_in[6647])
);

LUT6 #(
   .INIT(64'hbbd16048bbd16048)  
) LUT6_inst8884 (
   .O(to_level3[1108]),
   .I0(level4_in[6648]),
   .I1(level4_in[6649]),
   .I2(level4_in[6650]),
   .I3(level4_in[6651]),
   .I4(level4_in[6652]),
   .I5(level4_in[6653])
);

LUT6 #(
   .INIT(64'h28d4acb028d4acb0)  
) LUT6_inst8885 (
   .O(to_level3[1109]),
   .I0(level4_in[6654]),
   .I1(level4_in[6655]),
   .I2(level4_in[6656]),
   .I3(level4_in[6657]),
   .I4(level4_in[6658]),
   .I5(level4_in[6659])
);

LUT6 #(
   .INIT(64'h27bc0b8d27bc0b8d)  
) LUT6_inst8886 (
   .O(to_level3[1110]),
   .I0(level4_in[6660]),
   .I1(level4_in[6661]),
   .I2(level4_in[6662]),
   .I3(level4_in[6663]),
   .I4(level4_in[6664]),
   .I5(level4_in[6665])
);

LUT6 #(
   .INIT(64'he66a59dfe66a59df)  
) LUT6_inst8887 (
   .O(to_level3[1111]),
   .I0(level4_in[6666]),
   .I1(level4_in[6667]),
   .I2(level4_in[6668]),
   .I3(level4_in[6669]),
   .I4(level4_in[6670]),
   .I5(level4_in[6671])
);

LUT6 #(
   .INIT(64'h4a4678cb4a4678cb)  
) LUT6_inst8888 (
   .O(to_level3[1112]),
   .I0(level4_in[6672]),
   .I1(level4_in[6673]),
   .I2(level4_in[6674]),
   .I3(level4_in[6675]),
   .I4(level4_in[6676]),
   .I5(level4_in[6677])
);

LUT6 #(
   .INIT(64'h2197dbc92197dbc9)  
) LUT6_inst8889 (
   .O(to_level3[1113]),
   .I0(level4_in[6678]),
   .I1(level4_in[6679]),
   .I2(level4_in[6680]),
   .I3(level4_in[6681]),
   .I4(level4_in[6682]),
   .I5(level4_in[6683])
);

LUT6 #(
   .INIT(64'h6d98c7596d98c759)  
) LUT6_inst8890 (
   .O(to_level3[1114]),
   .I0(level4_in[6684]),
   .I1(level4_in[6685]),
   .I2(level4_in[6686]),
   .I3(level4_in[6687]),
   .I4(level4_in[6688]),
   .I5(level4_in[6689])
);

LUT6 #(
   .INIT(64'he68ae416e68ae416)  
) LUT6_inst8891 (
   .O(to_level3[1115]),
   .I0(level4_in[6690]),
   .I1(level4_in[6691]),
   .I2(level4_in[6692]),
   .I3(level4_in[6693]),
   .I4(level4_in[6694]),
   .I5(level4_in[6695])
);

LUT6 #(
   .INIT(64'h41aff63f41aff63f)  
) LUT6_inst8892 (
   .O(to_level3[1116]),
   .I0(level4_in[6696]),
   .I1(level4_in[6697]),
   .I2(level4_in[6698]),
   .I3(level4_in[6699]),
   .I4(level4_in[6700]),
   .I5(level4_in[6701])
);

LUT6 #(
   .INIT(64'h00789c2a00789c2a)  
) LUT6_inst8893 (
   .O(to_level3[1117]),
   .I0(level4_in[6702]),
   .I1(level4_in[6703]),
   .I2(level4_in[6704]),
   .I3(level4_in[6705]),
   .I4(level4_in[6706]),
   .I5(level4_in[6707])
);

LUT6 #(
   .INIT(64'h5e6a212b5e6a212b)  
) LUT6_inst8894 (
   .O(to_level3[1118]),
   .I0(level4_in[6708]),
   .I1(level4_in[6709]),
   .I2(level4_in[6710]),
   .I3(level4_in[6711]),
   .I4(level4_in[6712]),
   .I5(level4_in[6713])
);

LUT6 #(
   .INIT(64'ha5bfcd11a5bfcd11)  
) LUT6_inst8895 (
   .O(to_level3[1119]),
   .I0(level4_in[6714]),
   .I1(level4_in[6715]),
   .I2(level4_in[6716]),
   .I3(level4_in[6717]),
   .I4(level4_in[6718]),
   .I5(level4_in[6719])
);

LUT6 #(
   .INIT(64'h9beeaab39beeaab3)  
) LUT6_inst8896 (
   .O(to_level3[1120]),
   .I0(level4_in[6720]),
   .I1(level4_in[6721]),
   .I2(level4_in[6722]),
   .I3(level4_in[6723]),
   .I4(level4_in[6724]),
   .I5(level4_in[6725])
);

LUT6 #(
   .INIT(64'hffc41a37ffc41a37)  
) LUT6_inst8897 (
   .O(to_level3[1121]),
   .I0(level4_in[6726]),
   .I1(level4_in[6727]),
   .I2(level4_in[6728]),
   .I3(level4_in[6729]),
   .I4(level4_in[6730]),
   .I5(level4_in[6731])
);

LUT6 #(
   .INIT(64'he8a811bae8a811ba)  
) LUT6_inst8898 (
   .O(to_level3[1122]),
   .I0(level4_in[6732]),
   .I1(level4_in[6733]),
   .I2(level4_in[6734]),
   .I3(level4_in[6735]),
   .I4(level4_in[6736]),
   .I5(level4_in[6737])
);

LUT6 #(
   .INIT(64'hc75efca2c75efca2)  
) LUT6_inst8899 (
   .O(to_level3[1123]),
   .I0(level4_in[6738]),
   .I1(level4_in[6739]),
   .I2(level4_in[6740]),
   .I3(level4_in[6741]),
   .I4(level4_in[6742]),
   .I5(level4_in[6743])
);

LUT6 #(
   .INIT(64'hf95fa20af95fa20a)  
) LUT6_inst8900 (
   .O(to_level3[1124]),
   .I0(level4_in[6744]),
   .I1(level4_in[6745]),
   .I2(level4_in[6746]),
   .I3(level4_in[6747]),
   .I4(level4_in[6748]),
   .I5(level4_in[6749])
);

LUT6 #(
   .INIT(64'h1dceeb001dceeb00)  
) LUT6_inst8901 (
   .O(to_level3[1125]),
   .I0(level4_in[6750]),
   .I1(level4_in[6751]),
   .I2(level4_in[6752]),
   .I3(level4_in[6753]),
   .I4(level4_in[6754]),
   .I5(level4_in[6755])
);

LUT6 #(
   .INIT(64'hae33facfae33facf)  
) LUT6_inst8902 (
   .O(to_level3[1126]),
   .I0(level4_in[6756]),
   .I1(level4_in[6757]),
   .I2(level4_in[6758]),
   .I3(level4_in[6759]),
   .I4(level4_in[6760]),
   .I5(level4_in[6761])
);

LUT6 #(
   .INIT(64'hc6d8a71dc6d8a71d)  
) LUT6_inst8903 (
   .O(to_level3[1127]),
   .I0(level4_in[6762]),
   .I1(level4_in[6763]),
   .I2(level4_in[6764]),
   .I3(level4_in[6765]),
   .I4(level4_in[6766]),
   .I5(level4_in[6767])
);

LUT6 #(
   .INIT(64'h0f3677840f367784)  
) LUT6_inst8904 (
   .O(to_level3[1128]),
   .I0(level4_in[6768]),
   .I1(level4_in[6769]),
   .I2(level4_in[6770]),
   .I3(level4_in[6771]),
   .I4(level4_in[6772]),
   .I5(level4_in[6773])
);

LUT6 #(
   .INIT(64'h5001133c5001133c)  
) LUT6_inst8905 (
   .O(to_level3[1129]),
   .I0(level4_in[6774]),
   .I1(level4_in[6775]),
   .I2(level4_in[6776]),
   .I3(level4_in[6777]),
   .I4(level4_in[6778]),
   .I5(level4_in[6779])
);

LUT6 #(
   .INIT(64'h57f37d6557f37d65)  
) LUT6_inst8906 (
   .O(to_level3[1130]),
   .I0(level4_in[6780]),
   .I1(level4_in[6781]),
   .I2(level4_in[6782]),
   .I3(level4_in[6783]),
   .I4(level4_in[6784]),
   .I5(level4_in[6785])
);

LUT6 #(
   .INIT(64'h20a5ae5420a5ae54)  
) LUT6_inst8907 (
   .O(to_level3[1131]),
   .I0(level4_in[6786]),
   .I1(level4_in[6787]),
   .I2(level4_in[6788]),
   .I3(level4_in[6789]),
   .I4(level4_in[6790]),
   .I5(level4_in[6791])
);

LUT6 #(
   .INIT(64'h580e2132580e2132)  
) LUT6_inst8908 (
   .O(to_level3[1132]),
   .I0(level4_in[6792]),
   .I1(level4_in[6793]),
   .I2(level4_in[6794]),
   .I3(level4_in[6795]),
   .I4(level4_in[6796]),
   .I5(level4_in[6797])
);

LUT6 #(
   .INIT(64'hae12102cae12102c)  
) LUT6_inst8909 (
   .O(to_level3[1133]),
   .I0(level4_in[6798]),
   .I1(level4_in[6799]),
   .I2(level4_in[6800]),
   .I3(level4_in[6801]),
   .I4(level4_in[6802]),
   .I5(level4_in[6803])
);

LUT6 #(
   .INIT(64'h5ef7c5855ef7c585)  
) LUT6_inst8910 (
   .O(to_level3[1134]),
   .I0(level4_in[6804]),
   .I1(level4_in[6805]),
   .I2(level4_in[6806]),
   .I3(level4_in[6807]),
   .I4(level4_in[6808]),
   .I5(level4_in[6809])
);

LUT6 #(
   .INIT(64'h59a50f3d59a50f3d)  
) LUT6_inst8911 (
   .O(to_level3[1135]),
   .I0(level4_in[6810]),
   .I1(level4_in[6811]),
   .I2(level4_in[6812]),
   .I3(level4_in[6813]),
   .I4(level4_in[6814]),
   .I5(level4_in[6815])
);

LUT6 #(
   .INIT(64'h517cf1d9517cf1d9)  
) LUT6_inst8912 (
   .O(to_level3[1136]),
   .I0(level4_in[6816]),
   .I1(level4_in[6817]),
   .I2(level4_in[6818]),
   .I3(level4_in[6819]),
   .I4(level4_in[6820]),
   .I5(level4_in[6821])
);

LUT6 #(
   .INIT(64'hd5efbee6d5efbee6)  
) LUT6_inst8913 (
   .O(to_level3[1137]),
   .I0(level4_in[6822]),
   .I1(level4_in[6823]),
   .I2(level4_in[6824]),
   .I3(level4_in[6825]),
   .I4(level4_in[6826]),
   .I5(level4_in[6827])
);

LUT6 #(
   .INIT(64'h247a7db9247a7db9)  
) LUT6_inst8914 (
   .O(to_level3[1138]),
   .I0(level4_in[6828]),
   .I1(level4_in[6829]),
   .I2(level4_in[6830]),
   .I3(level4_in[6831]),
   .I4(level4_in[6832]),
   .I5(level4_in[6833])
);

LUT6 #(
   .INIT(64'h77b254dc77b254dc)  
) LUT6_inst8915 (
   .O(to_level3[1139]),
   .I0(level4_in[6834]),
   .I1(level4_in[6835]),
   .I2(level4_in[6836]),
   .I3(level4_in[6837]),
   .I4(level4_in[6838]),
   .I5(level4_in[6839])
);

LUT6 #(
   .INIT(64'h7c4ea9c97c4ea9c9)  
) LUT6_inst8916 (
   .O(to_level3[1140]),
   .I0(level4_in[6840]),
   .I1(level4_in[6841]),
   .I2(level4_in[6842]),
   .I3(level4_in[6843]),
   .I4(level4_in[6844]),
   .I5(level4_in[6845])
);

LUT6 #(
   .INIT(64'ha76b27fea76b27fe)  
) LUT6_inst8917 (
   .O(to_level3[1141]),
   .I0(level4_in[6846]),
   .I1(level4_in[6847]),
   .I2(level4_in[6848]),
   .I3(level4_in[6849]),
   .I4(level4_in[6850]),
   .I5(level4_in[6851])
);

LUT6 #(
   .INIT(64'h1ccc791e1ccc791e)  
) LUT6_inst8918 (
   .O(to_level3[1142]),
   .I0(level4_in[6852]),
   .I1(level4_in[6853]),
   .I2(level4_in[6854]),
   .I3(level4_in[6855]),
   .I4(level4_in[6856]),
   .I5(level4_in[6857])
);

LUT6 #(
   .INIT(64'hb5dd8556b5dd8556)  
) LUT6_inst8919 (
   .O(to_level3[1143]),
   .I0(level4_in[6858]),
   .I1(level4_in[6859]),
   .I2(level4_in[6860]),
   .I3(level4_in[6861]),
   .I4(level4_in[6862]),
   .I5(level4_in[6863])
);

LUT6 #(
   .INIT(64'he07a72f7e07a72f7)  
) LUT6_inst8920 (
   .O(to_level3[1144]),
   .I0(level4_in[6864]),
   .I1(level4_in[6865]),
   .I2(level4_in[6866]),
   .I3(level4_in[6867]),
   .I4(level4_in[6868]),
   .I5(level4_in[6869])
);

LUT6 #(
   .INIT(64'haaa610baaaa610ba)  
) LUT6_inst8921 (
   .O(to_level3[1145]),
   .I0(level4_in[6870]),
   .I1(level4_in[6871]),
   .I2(level4_in[6872]),
   .I3(level4_in[6873]),
   .I4(level4_in[6874]),
   .I5(level4_in[6875])
);

LUT6 #(
   .INIT(64'h42982d7e42982d7e)  
) LUT6_inst8922 (
   .O(to_level3[1146]),
   .I0(level4_in[6876]),
   .I1(level4_in[6877]),
   .I2(level4_in[6878]),
   .I3(level4_in[6879]),
   .I4(level4_in[6880]),
   .I5(level4_in[6881])
);

LUT6 #(
   .INIT(64'h4640f5514640f551)  
) LUT6_inst8923 (
   .O(to_level3[1147]),
   .I0(level4_in[6882]),
   .I1(level4_in[6883]),
   .I2(level4_in[6884]),
   .I3(level4_in[6885]),
   .I4(level4_in[6886]),
   .I5(level4_in[6887])
);

LUT6 #(
   .INIT(64'he93df727e93df727)  
) LUT6_inst8924 (
   .O(to_level3[1148]),
   .I0(level4_in[6888]),
   .I1(level4_in[6889]),
   .I2(level4_in[6890]),
   .I3(level4_in[6891]),
   .I4(level4_in[6892]),
   .I5(level4_in[6893])
);

LUT6 #(
   .INIT(64'h7806a9217806a921)  
) LUT6_inst8925 (
   .O(to_level3[1149]),
   .I0(level4_in[6894]),
   .I1(level4_in[6895]),
   .I2(level4_in[6896]),
   .I3(level4_in[6897]),
   .I4(level4_in[6898]),
   .I5(level4_in[6899])
);

LUT6 #(
   .INIT(64'h017f5775017f5775)  
) LUT6_inst8926 (
   .O(to_level3[1150]),
   .I0(level4_in[6900]),
   .I1(level4_in[6901]),
   .I2(level4_in[6902]),
   .I3(level4_in[6903]),
   .I4(level4_in[6904]),
   .I5(level4_in[6905])
);

LUT6 #(
   .INIT(64'h1c5e62041c5e6204)  
) LUT6_inst8927 (
   .O(to_level3[1151]),
   .I0(level4_in[6906]),
   .I1(level4_in[6907]),
   .I2(level4_in[6908]),
   .I3(level4_in[6909]),
   .I4(level4_in[6910]),
   .I5(level4_in[6911])
);

LUT6 #(
   .INIT(64'h86ae1bac86ae1bac)  
) LUT6_inst8928 (
   .O(to_level3[1152]),
   .I0(level4_in[6912]),
   .I1(level4_in[6913]),
   .I2(level4_in[6914]),
   .I3(level4_in[6915]),
   .I4(level4_in[6916]),
   .I5(level4_in[6917])
);

LUT6 #(
   .INIT(64'h60e931d760e931d7)  
) LUT6_inst8929 (
   .O(to_level3[1153]),
   .I0(level4_in[6918]),
   .I1(level4_in[6919]),
   .I2(level4_in[6920]),
   .I3(level4_in[6921]),
   .I4(level4_in[6922]),
   .I5(level4_in[6923])
);

LUT6 #(
   .INIT(64'h3c5e31203c5e3120)  
) LUT6_inst8930 (
   .O(to_level3[1154]),
   .I0(level4_in[6924]),
   .I1(level4_in[6925]),
   .I2(level4_in[6926]),
   .I3(level4_in[6927]),
   .I4(level4_in[6928]),
   .I5(level4_in[6929])
);

LUT6 #(
   .INIT(64'hf193fb64f193fb64)  
) LUT6_inst8931 (
   .O(to_level3[1155]),
   .I0(level4_in[6930]),
   .I1(level4_in[6931]),
   .I2(level4_in[6932]),
   .I3(level4_in[6933]),
   .I4(level4_in[6934]),
   .I5(level4_in[6935])
);

LUT6 #(
   .INIT(64'hbc5e306cbc5e306c)  
) LUT6_inst8932 (
   .O(to_level3[1156]),
   .I0(level4_in[6936]),
   .I1(level4_in[6937]),
   .I2(level4_in[6938]),
   .I3(level4_in[6939]),
   .I4(level4_in[6940]),
   .I5(level4_in[6941])
);

LUT6 #(
   .INIT(64'he5e69305e5e69305)  
) LUT6_inst8933 (
   .O(to_level3[1157]),
   .I0(level4_in[6942]),
   .I1(level4_in[6943]),
   .I2(level4_in[6944]),
   .I3(level4_in[6945]),
   .I4(level4_in[6946]),
   .I5(level4_in[6947])
);

LUT6 #(
   .INIT(64'hda27445dda27445d)  
) LUT6_inst8934 (
   .O(to_level3[1158]),
   .I0(level4_in[6948]),
   .I1(level4_in[6949]),
   .I2(level4_in[6950]),
   .I3(level4_in[6951]),
   .I4(level4_in[6952]),
   .I5(level4_in[6953])
);

LUT6 #(
   .INIT(64'hc3b13719c3b13719)  
) LUT6_inst8935 (
   .O(to_level3[1159]),
   .I0(level4_in[6954]),
   .I1(level4_in[6955]),
   .I2(level4_in[6956]),
   .I3(level4_in[6957]),
   .I4(level4_in[6958]),
   .I5(level4_in[6959])
);

LUT6 #(
   .INIT(64'h73c3351c73c3351c)  
) LUT6_inst8936 (
   .O(to_level3[1160]),
   .I0(level4_in[6960]),
   .I1(level4_in[6961]),
   .I2(level4_in[6962]),
   .I3(level4_in[6963]),
   .I4(level4_in[6964]),
   .I5(level4_in[6965])
);

LUT6 #(
   .INIT(64'h20cf25a220cf25a2)  
) LUT6_inst8937 (
   .O(to_level3[1161]),
   .I0(level4_in[6966]),
   .I1(level4_in[6967]),
   .I2(level4_in[6968]),
   .I3(level4_in[6969]),
   .I4(level4_in[6970]),
   .I5(level4_in[6971])
);

LUT6 #(
   .INIT(64'hd617a478d617a478)  
) LUT6_inst8938 (
   .O(to_level3[1162]),
   .I0(level4_in[6972]),
   .I1(level4_in[6973]),
   .I2(level4_in[6974]),
   .I3(level4_in[6975]),
   .I4(level4_in[6976]),
   .I5(level4_in[6977])
);

LUT6 #(
   .INIT(64'h35753b5a35753b5a)  
) LUT6_inst8939 (
   .O(to_level3[1163]),
   .I0(level4_in[6978]),
   .I1(level4_in[6979]),
   .I2(level4_in[6980]),
   .I3(level4_in[6981]),
   .I4(level4_in[6982]),
   .I5(level4_in[6983])
);

LUT6 #(
   .INIT(64'h8ace33f28ace33f2)  
) LUT6_inst8940 (
   .O(to_level3[1164]),
   .I0(level4_in[6984]),
   .I1(level4_in[6985]),
   .I2(level4_in[6986]),
   .I3(level4_in[6987]),
   .I4(level4_in[6988]),
   .I5(level4_in[6989])
);

LUT6 #(
   .INIT(64'h5d6b9c665d6b9c66)  
) LUT6_inst8941 (
   .O(to_level3[1165]),
   .I0(level4_in[6990]),
   .I1(level4_in[6991]),
   .I2(level4_in[6992]),
   .I3(level4_in[6993]),
   .I4(level4_in[6994]),
   .I5(level4_in[6995])
);

LUT6 #(
   .INIT(64'hde8291c1de8291c1)  
) LUT6_inst8942 (
   .O(to_level3[1166]),
   .I0(level4_in[6996]),
   .I1(level4_in[6997]),
   .I2(level4_in[6998]),
   .I3(level4_in[6999]),
   .I4(level4_in[7000]),
   .I5(level4_in[7001])
);

LUT6 #(
   .INIT(64'hede43a01ede43a01)  
) LUT6_inst8943 (
   .O(to_level3[1167]),
   .I0(level4_in[7002]),
   .I1(level4_in[7003]),
   .I2(level4_in[7004]),
   .I3(level4_in[7005]),
   .I4(level4_in[7006]),
   .I5(level4_in[7007])
);

LUT6 #(
   .INIT(64'h9137d1039137d103)  
) LUT6_inst8944 (
   .O(to_level3[1168]),
   .I0(level4_in[7008]),
   .I1(level4_in[7009]),
   .I2(level4_in[7010]),
   .I3(level4_in[7011]),
   .I4(level4_in[7012]),
   .I5(level4_in[7013])
);

LUT6 #(
   .INIT(64'h9ddbd6699ddbd669)  
) LUT6_inst8945 (
   .O(to_level3[1169]),
   .I0(level4_in[7014]),
   .I1(level4_in[7015]),
   .I2(level4_in[7016]),
   .I3(level4_in[7017]),
   .I4(level4_in[7018]),
   .I5(level4_in[7019])
);

LUT6 #(
   .INIT(64'h89e519e489e519e4)  
) LUT6_inst8946 (
   .O(to_level3[1170]),
   .I0(level4_in[7020]),
   .I1(level4_in[7021]),
   .I2(level4_in[7022]),
   .I3(level4_in[7023]),
   .I4(level4_in[7024]),
   .I5(level4_in[7025])
);

LUT6 #(
   .INIT(64'h562b12b6562b12b6)  
) LUT6_inst8947 (
   .O(to_level3[1171]),
   .I0(level4_in[7026]),
   .I1(level4_in[7027]),
   .I2(level4_in[7028]),
   .I3(level4_in[7029]),
   .I4(level4_in[7030]),
   .I5(level4_in[7031])
);

LUT6 #(
   .INIT(64'h502014d8502014d8)  
) LUT6_inst8948 (
   .O(to_level3[1172]),
   .I0(level4_in[7032]),
   .I1(level4_in[7033]),
   .I2(level4_in[7034]),
   .I3(level4_in[7035]),
   .I4(level4_in[7036]),
   .I5(level4_in[7037])
);

LUT6 #(
   .INIT(64'hc6699184c6699184)  
) LUT6_inst8949 (
   .O(to_level3[1173]),
   .I0(level4_in[7038]),
   .I1(level4_in[7039]),
   .I2(level4_in[7040]),
   .I3(level4_in[7041]),
   .I4(level4_in[7042]),
   .I5(level4_in[7043])
);

LUT6 #(
   .INIT(64'h9de635639de63563)  
) LUT6_inst8950 (
   .O(to_level3[1174]),
   .I0(level4_in[7044]),
   .I1(level4_in[7045]),
   .I2(level4_in[7046]),
   .I3(level4_in[7047]),
   .I4(level4_in[7048]),
   .I5(level4_in[7049])
);

LUT6 #(
   .INIT(64'hff8f0eb1ff8f0eb1)  
) LUT6_inst8951 (
   .O(to_level3[1175]),
   .I0(level4_in[7050]),
   .I1(level4_in[7051]),
   .I2(level4_in[7052]),
   .I3(level4_in[7053]),
   .I4(level4_in[7054]),
   .I5(level4_in[7055])
);

LUT6 #(
   .INIT(64'h31c36ab731c36ab7)  
) LUT6_inst8952 (
   .O(to_level3[1176]),
   .I0(level4_in[7056]),
   .I1(level4_in[7057]),
   .I2(level4_in[7058]),
   .I3(level4_in[7059]),
   .I4(level4_in[7060]),
   .I5(level4_in[7061])
);

LUT6 #(
   .INIT(64'hc1558671c1558671)  
) LUT6_inst8953 (
   .O(to_level3[1177]),
   .I0(level4_in[7062]),
   .I1(level4_in[7063]),
   .I2(level4_in[7064]),
   .I3(level4_in[7065]),
   .I4(level4_in[7066]),
   .I5(level4_in[7067])
);

LUT6 #(
   .INIT(64'h69329b4b69329b4b)  
) LUT6_inst8954 (
   .O(to_level3[1178]),
   .I0(level4_in[7068]),
   .I1(level4_in[7069]),
   .I2(level4_in[7070]),
   .I3(level4_in[7071]),
   .I4(level4_in[7072]),
   .I5(level4_in[7073])
);

LUT6 #(
   .INIT(64'h0e6e95cd0e6e95cd)  
) LUT6_inst8955 (
   .O(to_level3[1179]),
   .I0(level4_in[7074]),
   .I1(level4_in[7075]),
   .I2(level4_in[7076]),
   .I3(level4_in[7077]),
   .I4(level4_in[7078]),
   .I5(level4_in[7079])
);

LUT6 #(
   .INIT(64'hb372a177b372a177)  
) LUT6_inst8956 (
   .O(to_level3[1180]),
   .I0(level4_in[7080]),
   .I1(level4_in[7081]),
   .I2(level4_in[7082]),
   .I3(level4_in[7083]),
   .I4(level4_in[7084]),
   .I5(level4_in[7085])
);

LUT6 #(
   .INIT(64'h7d4c1b597d4c1b59)  
) LUT6_inst8957 (
   .O(to_level3[1181]),
   .I0(level4_in[7086]),
   .I1(level4_in[7087]),
   .I2(level4_in[7088]),
   .I3(level4_in[7089]),
   .I4(level4_in[7090]),
   .I5(level4_in[7091])
);

LUT6 #(
   .INIT(64'h5ed15f5e5ed15f5e)  
) LUT6_inst8958 (
   .O(to_level3[1182]),
   .I0(level4_in[7092]),
   .I1(level4_in[7093]),
   .I2(level4_in[7094]),
   .I3(level4_in[7095]),
   .I4(level4_in[7096]),
   .I5(level4_in[7097])
);

LUT6 #(
   .INIT(64'hdb80ca83db80ca83)  
) LUT6_inst8959 (
   .O(to_level3[1183]),
   .I0(level4_in[7098]),
   .I1(level4_in[7099]),
   .I2(level4_in[7100]),
   .I3(level4_in[7101]),
   .I4(level4_in[7102]),
   .I5(level4_in[7103])
);

LUT6 #(
   .INIT(64'h1ac7f0d31ac7f0d3)  
) LUT6_inst8960 (
   .O(to_level3[1184]),
   .I0(level4_in[7104]),
   .I1(level4_in[7105]),
   .I2(level4_in[7106]),
   .I3(level4_in[7107]),
   .I4(level4_in[7108]),
   .I5(level4_in[7109])
);

LUT6 #(
   .INIT(64'h6deff0f86deff0f8)  
) LUT6_inst8961 (
   .O(to_level3[1185]),
   .I0(level4_in[7110]),
   .I1(level4_in[7111]),
   .I2(level4_in[7112]),
   .I3(level4_in[7113]),
   .I4(level4_in[7114]),
   .I5(level4_in[7115])
);

LUT6 #(
   .INIT(64'hb1e1dffbb1e1dffb)  
) LUT6_inst8962 (
   .O(to_level3[1186]),
   .I0(level4_in[7116]),
   .I1(level4_in[7117]),
   .I2(level4_in[7118]),
   .I3(level4_in[7119]),
   .I4(level4_in[7120]),
   .I5(level4_in[7121])
);

LUT6 #(
   .INIT(64'h93830f2f93830f2f)  
) LUT6_inst8963 (
   .O(to_level3[1187]),
   .I0(level4_in[7122]),
   .I1(level4_in[7123]),
   .I2(level4_in[7124]),
   .I3(level4_in[7125]),
   .I4(level4_in[7126]),
   .I5(level4_in[7127])
);

LUT6 #(
   .INIT(64'hbf570ff1bf570ff1)  
) LUT6_inst8964 (
   .O(to_level3[1188]),
   .I0(level4_in[7128]),
   .I1(level4_in[7129]),
   .I2(level4_in[7130]),
   .I3(level4_in[7131]),
   .I4(level4_in[7132]),
   .I5(level4_in[7133])
);

LUT6 #(
   .INIT(64'h48fb46f748fb46f7)  
) LUT6_inst8965 (
   .O(to_level3[1189]),
   .I0(level4_in[7134]),
   .I1(level4_in[7135]),
   .I2(level4_in[7136]),
   .I3(level4_in[7137]),
   .I4(level4_in[7138]),
   .I5(level4_in[7139])
);

LUT6 #(
   .INIT(64'hceaaf734ceaaf734)  
) LUT6_inst8966 (
   .O(to_level3[1190]),
   .I0(level4_in[7140]),
   .I1(level4_in[7141]),
   .I2(level4_in[7142]),
   .I3(level4_in[7143]),
   .I4(level4_in[7144]),
   .I5(level4_in[7145])
);

LUT6 #(
   .INIT(64'h386e2f8c386e2f8c)  
) LUT6_inst8967 (
   .O(to_level3[1191]),
   .I0(level4_in[7146]),
   .I1(level4_in[7147]),
   .I2(level4_in[7148]),
   .I3(level4_in[7149]),
   .I4(level4_in[7150]),
   .I5(level4_in[7151])
);

LUT6 #(
   .INIT(64'haf0cedbcaf0cedbc)  
) LUT6_inst8968 (
   .O(to_level3[1192]),
   .I0(level4_in[7152]),
   .I1(level4_in[7153]),
   .I2(level4_in[7154]),
   .I3(level4_in[7155]),
   .I4(level4_in[7156]),
   .I5(level4_in[7157])
);

LUT6 #(
   .INIT(64'h9b9277739b927773)  
) LUT6_inst8969 (
   .O(to_level3[1193]),
   .I0(level4_in[7158]),
   .I1(level4_in[7159]),
   .I2(level4_in[7160]),
   .I3(level4_in[7161]),
   .I4(level4_in[7162]),
   .I5(level4_in[7163])
);

LUT6 #(
   .INIT(64'h847befca847befca)  
) LUT6_inst8970 (
   .O(to_level3[1194]),
   .I0(level4_in[7164]),
   .I1(level4_in[7165]),
   .I2(level4_in[7166]),
   .I3(level4_in[7167]),
   .I4(level4_in[7168]),
   .I5(level4_in[7169])
);

LUT6 #(
   .INIT(64'hb0336515b0336515)  
) LUT6_inst8971 (
   .O(to_level3[1195]),
   .I0(level4_in[7170]),
   .I1(level4_in[7171]),
   .I2(level4_in[7172]),
   .I3(level4_in[7173]),
   .I4(level4_in[7174]),
   .I5(level4_in[7175])
);

LUT6 #(
   .INIT(64'hfbdb0baefbdb0bae)  
) LUT6_inst8972 (
   .O(to_level3[1196]),
   .I0(level4_in[7176]),
   .I1(level4_in[7177]),
   .I2(level4_in[7178]),
   .I3(level4_in[7179]),
   .I4(level4_in[7180]),
   .I5(level4_in[7181])
);

LUT6 #(
   .INIT(64'hb6e28a48b6e28a48)  
) LUT6_inst8973 (
   .O(to_level3[1197]),
   .I0(level4_in[7182]),
   .I1(level4_in[7183]),
   .I2(level4_in[7184]),
   .I3(level4_in[7185]),
   .I4(level4_in[7186]),
   .I5(level4_in[7187])
);

LUT6 #(
   .INIT(64'h060e5c11060e5c11)  
) LUT6_inst8974 (
   .O(to_level3[1198]),
   .I0(level4_in[7188]),
   .I1(level4_in[7189]),
   .I2(level4_in[7190]),
   .I3(level4_in[7191]),
   .I4(level4_in[7192]),
   .I5(level4_in[7193])
);

LUT6 #(
   .INIT(64'hf63a5607f63a5607)  
) LUT6_inst8975 (
   .O(to_level3[1199]),
   .I0(level4_in[7194]),
   .I1(level4_in[7195]),
   .I2(level4_in[7196]),
   .I3(level4_in[7197]),
   .I4(level4_in[7198]),
   .I5(level4_in[7199])
);

LUT6 #(
   .INIT(64'h98e0330098e03300)  
) LUT6_inst8976 (
   .O(to_level3[1200]),
   .I0(level4_in[7200]),
   .I1(level4_in[7201]),
   .I2(level4_in[7202]),
   .I3(level4_in[7203]),
   .I4(level4_in[7204]),
   .I5(level4_in[7205])
);

LUT6 #(
   .INIT(64'hfe2fd3f1fe2fd3f1)  
) LUT6_inst8977 (
   .O(to_level3[1201]),
   .I0(level4_in[7206]),
   .I1(level4_in[7207]),
   .I2(level4_in[7208]),
   .I3(level4_in[7209]),
   .I4(level4_in[7210]),
   .I5(level4_in[7211])
);

LUT6 #(
   .INIT(64'h3ce35f293ce35f29)  
) LUT6_inst8978 (
   .O(to_level3[1202]),
   .I0(level4_in[7212]),
   .I1(level4_in[7213]),
   .I2(level4_in[7214]),
   .I3(level4_in[7215]),
   .I4(level4_in[7216]),
   .I5(level4_in[7217])
);

LUT6 #(
   .INIT(64'ha9d4032ea9d4032e)  
) LUT6_inst8979 (
   .O(to_level3[1203]),
   .I0(level4_in[7218]),
   .I1(level4_in[7219]),
   .I2(level4_in[7220]),
   .I3(level4_in[7221]),
   .I4(level4_in[7222]),
   .I5(level4_in[7223])
);

LUT6 #(
   .INIT(64'h7292cc9e7292cc9e)  
) LUT6_inst8980 (
   .O(to_level3[1204]),
   .I0(level4_in[7224]),
   .I1(level4_in[7225]),
   .I2(level4_in[7226]),
   .I3(level4_in[7227]),
   .I4(level4_in[7228]),
   .I5(level4_in[7229])
);

LUT6 #(
   .INIT(64'h8ce604ac8ce604ac)  
) LUT6_inst8981 (
   .O(to_level3[1205]),
   .I0(level4_in[7230]),
   .I1(level4_in[7231]),
   .I2(level4_in[7232]),
   .I3(level4_in[7233]),
   .I4(level4_in[7234]),
   .I5(level4_in[7235])
);

LUT6 #(
   .INIT(64'hd41356a6d41356a6)  
) LUT6_inst8982 (
   .O(to_level3[1206]),
   .I0(level4_in[7236]),
   .I1(level4_in[7237]),
   .I2(level4_in[7238]),
   .I3(level4_in[7239]),
   .I4(level4_in[7240]),
   .I5(level4_in[7241])
);

LUT6 #(
   .INIT(64'h9d8aedf89d8aedf8)  
) LUT6_inst8983 (
   .O(to_level3[1207]),
   .I0(level4_in[7242]),
   .I1(level4_in[7243]),
   .I2(level4_in[7244]),
   .I3(level4_in[7245]),
   .I4(level4_in[7246]),
   .I5(level4_in[7247])
);

LUT6 #(
   .INIT(64'h464e6af3464e6af3)  
) LUT6_inst8984 (
   .O(to_level3[1208]),
   .I0(level4_in[7248]),
   .I1(level4_in[7249]),
   .I2(level4_in[7250]),
   .I3(level4_in[7251]),
   .I4(level4_in[7252]),
   .I5(level4_in[7253])
);

LUT6 #(
   .INIT(64'h9faf49179faf4917)  
) LUT6_inst8985 (
   .O(to_level3[1209]),
   .I0(level4_in[7254]),
   .I1(level4_in[7255]),
   .I2(level4_in[7256]),
   .I3(level4_in[7257]),
   .I4(level4_in[7258]),
   .I5(level4_in[7259])
);

LUT6 #(
   .INIT(64'hbd923becbd923bec)  
) LUT6_inst8986 (
   .O(to_level3[1210]),
   .I0(level4_in[7260]),
   .I1(level4_in[7261]),
   .I2(level4_in[7262]),
   .I3(level4_in[7263]),
   .I4(level4_in[7264]),
   .I5(level4_in[7265])
);

LUT6 #(
   .INIT(64'h4a0fef924a0fef92)  
) LUT6_inst8987 (
   .O(to_level3[1211]),
   .I0(level4_in[7266]),
   .I1(level4_in[7267]),
   .I2(level4_in[7268]),
   .I3(level4_in[7269]),
   .I4(level4_in[7270]),
   .I5(level4_in[7271])
);

LUT6 #(
   .INIT(64'hc9991e5ac9991e5a)  
) LUT6_inst8988 (
   .O(to_level3[1212]),
   .I0(level4_in[7272]),
   .I1(level4_in[7273]),
   .I2(level4_in[7274]),
   .I3(level4_in[7275]),
   .I4(level4_in[7276]),
   .I5(level4_in[7277])
);

LUT6 #(
   .INIT(64'h29562cce29562cce)  
) LUT6_inst8989 (
   .O(to_level3[1213]),
   .I0(level4_in[7278]),
   .I1(level4_in[7279]),
   .I2(level4_in[7280]),
   .I3(level4_in[7281]),
   .I4(level4_in[7282]),
   .I5(level4_in[7283])
);

LUT6 #(
   .INIT(64'h7ea944ff7ea944ff)  
) LUT6_inst8990 (
   .O(to_level3[1214]),
   .I0(level4_in[7284]),
   .I1(level4_in[7285]),
   .I2(level4_in[7286]),
   .I3(level4_in[7287]),
   .I4(level4_in[7288]),
   .I5(level4_in[7289])
);

LUT6 #(
   .INIT(64'h2d4d2fca2d4d2fca)  
) LUT6_inst8991 (
   .O(to_level3[1215]),
   .I0(level4_in[7290]),
   .I1(level4_in[7291]),
   .I2(level4_in[7292]),
   .I3(level4_in[7293]),
   .I4(level4_in[7294]),
   .I5(level4_in[7295])
);

LUT6 #(
   .INIT(64'h8253646182536461)  
) LUT6_inst8992 (
   .O(to_level3[1216]),
   .I0(level4_in[7296]),
   .I1(level4_in[7297]),
   .I2(level4_in[7298]),
   .I3(level4_in[7299]),
   .I4(level4_in[7300]),
   .I5(level4_in[7301])
);

LUT6 #(
   .INIT(64'h30c392c230c392c2)  
) LUT6_inst8993 (
   .O(to_level3[1217]),
   .I0(level4_in[7302]),
   .I1(level4_in[7303]),
   .I2(level4_in[7304]),
   .I3(level4_in[7305]),
   .I4(level4_in[7306]),
   .I5(level4_in[7307])
);

LUT6 #(
   .INIT(64'h818c3563818c3563)  
) LUT6_inst8994 (
   .O(to_level3[1218]),
   .I0(level4_in[7308]),
   .I1(level4_in[7309]),
   .I2(level4_in[7310]),
   .I3(level4_in[7311]),
   .I4(level4_in[7312]),
   .I5(level4_in[7313])
);

LUT6 #(
   .INIT(64'ha737530fa737530f)  
) LUT6_inst8995 (
   .O(to_level3[1219]),
   .I0(level4_in[7314]),
   .I1(level4_in[7315]),
   .I2(level4_in[7316]),
   .I3(level4_in[7317]),
   .I4(level4_in[7318]),
   .I5(level4_in[7319])
);

LUT6 #(
   .INIT(64'h0e7427c30e7427c3)  
) LUT6_inst8996 (
   .O(to_level3[1220]),
   .I0(level4_in[7320]),
   .I1(level4_in[7321]),
   .I2(level4_in[7322]),
   .I3(level4_in[7323]),
   .I4(level4_in[7324]),
   .I5(level4_in[7325])
);

LUT6 #(
   .INIT(64'h71250ff071250ff0)  
) LUT6_inst8997 (
   .O(to_level3[1221]),
   .I0(level4_in[7326]),
   .I1(level4_in[7327]),
   .I2(level4_in[7328]),
   .I3(level4_in[7329]),
   .I4(level4_in[7330]),
   .I5(level4_in[7331])
);

LUT6 #(
   .INIT(64'h75d51e9e75d51e9e)  
) LUT6_inst8998 (
   .O(to_level3[1222]),
   .I0(level4_in[7332]),
   .I1(level4_in[7333]),
   .I2(level4_in[7334]),
   .I3(level4_in[7335]),
   .I4(level4_in[7336]),
   .I5(level4_in[7337])
);

LUT6 #(
   .INIT(64'h2e0a9b612e0a9b61)  
) LUT6_inst8999 (
   .O(to_level3[1223]),
   .I0(level4_in[7338]),
   .I1(level4_in[7339]),
   .I2(level4_in[7340]),
   .I3(level4_in[7341]),
   .I4(level4_in[7342]),
   .I5(level4_in[7343])
);

LUT6 #(
   .INIT(64'had0abb7fad0abb7f)  
) LUT6_inst9000 (
   .O(to_level3[1224]),
   .I0(level4_in[7344]),
   .I1(level4_in[7345]),
   .I2(level4_in[7346]),
   .I3(level4_in[7347]),
   .I4(level4_in[7348]),
   .I5(level4_in[7349])
);

LUT6 #(
   .INIT(64'hdbb421b8dbb421b8)  
) LUT6_inst9001 (
   .O(to_level3[1225]),
   .I0(level4_in[7350]),
   .I1(level4_in[7351]),
   .I2(level4_in[7352]),
   .I3(level4_in[7353]),
   .I4(level4_in[7354]),
   .I5(level4_in[7355])
);

LUT6 #(
   .INIT(64'h9c396a759c396a75)  
) LUT6_inst9002 (
   .O(to_level3[1226]),
   .I0(level4_in[7356]),
   .I1(level4_in[7357]),
   .I2(level4_in[7358]),
   .I3(level4_in[7359]),
   .I4(level4_in[7360]),
   .I5(level4_in[7361])
);

LUT6 #(
   .INIT(64'hbc0955bfbc0955bf)  
) LUT6_inst9003 (
   .O(to_level3[1227]),
   .I0(level4_in[7362]),
   .I1(level4_in[7363]),
   .I2(level4_in[7364]),
   .I3(level4_in[7365]),
   .I4(level4_in[7366]),
   .I5(level4_in[7367])
);

LUT6 #(
   .INIT(64'hb55ea461b55ea461)  
) LUT6_inst9004 (
   .O(to_level3[1228]),
   .I0(level4_in[7368]),
   .I1(level4_in[7369]),
   .I2(level4_in[7370]),
   .I3(level4_in[7371]),
   .I4(level4_in[7372]),
   .I5(level4_in[7373])
);

LUT6 #(
   .INIT(64'hd3c1241bd3c1241b)  
) LUT6_inst9005 (
   .O(to_level3[1229]),
   .I0(level4_in[7374]),
   .I1(level4_in[7375]),
   .I2(level4_in[7376]),
   .I3(level4_in[7377]),
   .I4(level4_in[7378]),
   .I5(level4_in[7379])
);

LUT6 #(
   .INIT(64'h1e6502be1e6502be)  
) LUT6_inst9006 (
   .O(to_level3[1230]),
   .I0(level4_in[7380]),
   .I1(level4_in[7381]),
   .I2(level4_in[7382]),
   .I3(level4_in[7383]),
   .I4(level4_in[7384]),
   .I5(level4_in[7385])
);

LUT6 #(
   .INIT(64'h8fc17b498fc17b49)  
) LUT6_inst9007 (
   .O(to_level3[1231]),
   .I0(level4_in[7386]),
   .I1(level4_in[7387]),
   .I2(level4_in[7388]),
   .I3(level4_in[7389]),
   .I4(level4_in[7390]),
   .I5(level4_in[7391])
);

LUT6 #(
   .INIT(64'h7fa130f97fa130f9)  
) LUT6_inst9008 (
   .O(to_level3[1232]),
   .I0(level4_in[7392]),
   .I1(level4_in[7393]),
   .I2(level4_in[7394]),
   .I3(level4_in[7395]),
   .I4(level4_in[7396]),
   .I5(level4_in[7397])
);

LUT6 #(
   .INIT(64'h22f4a0d822f4a0d8)  
) LUT6_inst9009 (
   .O(to_level3[1233]),
   .I0(level4_in[7398]),
   .I1(level4_in[7399]),
   .I2(level4_in[7400]),
   .I3(level4_in[7401]),
   .I4(level4_in[7402]),
   .I5(level4_in[7403])
);

LUT6 #(
   .INIT(64'h387d5c80387d5c80)  
) LUT6_inst9010 (
   .O(to_level3[1234]),
   .I0(level4_in[7404]),
   .I1(level4_in[7405]),
   .I2(level4_in[7406]),
   .I3(level4_in[7407]),
   .I4(level4_in[7408]),
   .I5(level4_in[7409])
);

LUT6 #(
   .INIT(64'h9cc631409cc63140)  
) LUT6_inst9011 (
   .O(to_level3[1235]),
   .I0(level4_in[7410]),
   .I1(level4_in[7411]),
   .I2(level4_in[7412]),
   .I3(level4_in[7413]),
   .I4(level4_in[7414]),
   .I5(level4_in[7415])
);

LUT6 #(
   .INIT(64'hfbadeb36fbadeb36)  
) LUT6_inst9012 (
   .O(to_level3[1236]),
   .I0(level4_in[7416]),
   .I1(level4_in[7417]),
   .I2(level4_in[7418]),
   .I3(level4_in[7419]),
   .I4(level4_in[7420]),
   .I5(level4_in[7421])
);

LUT6 #(
   .INIT(64'h260f9a50260f9a50)  
) LUT6_inst9013 (
   .O(to_level3[1237]),
   .I0(level4_in[7422]),
   .I1(level4_in[7423]),
   .I2(level4_in[7424]),
   .I3(level4_in[7425]),
   .I4(level4_in[7426]),
   .I5(level4_in[7427])
);

LUT6 #(
   .INIT(64'h098f08f1098f08f1)  
) LUT6_inst9014 (
   .O(to_level3[1238]),
   .I0(level4_in[7428]),
   .I1(level4_in[7429]),
   .I2(level4_in[7430]),
   .I3(level4_in[7431]),
   .I4(level4_in[7432]),
   .I5(level4_in[7433])
);

LUT6 #(
   .INIT(64'hda086d45da086d45)  
) LUT6_inst9015 (
   .O(to_level3[1239]),
   .I0(level4_in[7434]),
   .I1(level4_in[7435]),
   .I2(level4_in[7436]),
   .I3(level4_in[7437]),
   .I4(level4_in[7438]),
   .I5(level4_in[7439])
);

LUT6 #(
   .INIT(64'h3b028c063b028c06)  
) LUT6_inst9016 (
   .O(to_level3[1240]),
   .I0(level4_in[7440]),
   .I1(level4_in[7441]),
   .I2(level4_in[7442]),
   .I3(level4_in[7443]),
   .I4(level4_in[7444]),
   .I5(level4_in[7445])
);

LUT6 #(
   .INIT(64'h4fcb62b54fcb62b5)  
) LUT6_inst9017 (
   .O(to_level3[1241]),
   .I0(level4_in[7446]),
   .I1(level4_in[7447]),
   .I2(level4_in[7448]),
   .I3(level4_in[7449]),
   .I4(level4_in[7450]),
   .I5(level4_in[7451])
);

LUT6 #(
   .INIT(64'h88e1267b88e1267b)  
) LUT6_inst9018 (
   .O(to_level3[1242]),
   .I0(level4_in[7452]),
   .I1(level4_in[7453]),
   .I2(level4_in[7454]),
   .I3(level4_in[7455]),
   .I4(level4_in[7456]),
   .I5(level4_in[7457])
);

LUT6 #(
   .INIT(64'h144bfcda144bfcda)  
) LUT6_inst9019 (
   .O(to_level3[1243]),
   .I0(level4_in[7458]),
   .I1(level4_in[7459]),
   .I2(level4_in[7460]),
   .I3(level4_in[7461]),
   .I4(level4_in[7462]),
   .I5(level4_in[7463])
);

LUT6 #(
   .INIT(64'h45ac89c945ac89c9)  
) LUT6_inst9020 (
   .O(to_level3[1244]),
   .I0(level4_in[7464]),
   .I1(level4_in[7465]),
   .I2(level4_in[7466]),
   .I3(level4_in[7467]),
   .I4(level4_in[7468]),
   .I5(level4_in[7469])
);

LUT6 #(
   .INIT(64'hc65cd6aac65cd6aa)  
) LUT6_inst9021 (
   .O(to_level3[1245]),
   .I0(level4_in[7470]),
   .I1(level4_in[7471]),
   .I2(level4_in[7472]),
   .I3(level4_in[7473]),
   .I4(level4_in[7474]),
   .I5(level4_in[7475])
);

LUT6 #(
   .INIT(64'h7df251537df25153)  
) LUT6_inst9022 (
   .O(to_level3[1246]),
   .I0(level4_in[7476]),
   .I1(level4_in[7477]),
   .I2(level4_in[7478]),
   .I3(level4_in[7479]),
   .I4(level4_in[7480]),
   .I5(level4_in[7481])
);

LUT6 #(
   .INIT(64'h0ccf8be10ccf8be1)  
) LUT6_inst9023 (
   .O(to_level3[1247]),
   .I0(level4_in[7482]),
   .I1(level4_in[7483]),
   .I2(level4_in[7484]),
   .I3(level4_in[7485]),
   .I4(level4_in[7486]),
   .I5(level4_in[7487])
);

LUT6 #(
   .INIT(64'hd78c8170d78c8170)  
) LUT6_inst9024 (
   .O(to_level3[1248]),
   .I0(level4_in[7488]),
   .I1(level4_in[7489]),
   .I2(level4_in[7490]),
   .I3(level4_in[7491]),
   .I4(level4_in[7492]),
   .I5(level4_in[7493])
);

LUT6 #(
   .INIT(64'hd4cc3070d4cc3070)  
) LUT6_inst9025 (
   .O(to_level3[1249]),
   .I0(level4_in[7494]),
   .I1(level4_in[7495]),
   .I2(level4_in[7496]),
   .I3(level4_in[7497]),
   .I4(level4_in[7498]),
   .I5(level4_in[7499])
);

LUT6 #(
   .INIT(64'hc7586e84c7586e84)  
) LUT6_inst9026 (
   .O(to_level3[1250]),
   .I0(level4_in[7500]),
   .I1(level4_in[7501]),
   .I2(level4_in[7502]),
   .I3(level4_in[7503]),
   .I4(level4_in[7504]),
   .I5(level4_in[7505])
);

LUT6 #(
   .INIT(64'h67cbf12d67cbf12d)  
) LUT6_inst9027 (
   .O(to_level3[1251]),
   .I0(level4_in[7506]),
   .I1(level4_in[7507]),
   .I2(level4_in[7508]),
   .I3(level4_in[7509]),
   .I4(level4_in[7510]),
   .I5(level4_in[7511])
);

LUT6 #(
   .INIT(64'hb1dfc3fbb1dfc3fb)  
) LUT6_inst9028 (
   .O(to_level3[1252]),
   .I0(level4_in[7512]),
   .I1(level4_in[7513]),
   .I2(level4_in[7514]),
   .I3(level4_in[7515]),
   .I4(level4_in[7516]),
   .I5(level4_in[7517])
);

LUT6 #(
   .INIT(64'h999e072a999e072a)  
) LUT6_inst9029 (
   .O(to_level3[1253]),
   .I0(level4_in[7518]),
   .I1(level4_in[7519]),
   .I2(level4_in[7520]),
   .I3(level4_in[7521]),
   .I4(level4_in[7522]),
   .I5(level4_in[7523])
);

LUT6 #(
   .INIT(64'h28d3d29528d3d295)  
) LUT6_inst9030 (
   .O(to_level3[1254]),
   .I0(level4_in[7524]),
   .I1(level4_in[7525]),
   .I2(level4_in[7526]),
   .I3(level4_in[7527]),
   .I4(level4_in[7528]),
   .I5(level4_in[7529])
);

LUT6 #(
   .INIT(64'hbfad95f1bfad95f1)  
) LUT6_inst9031 (
   .O(to_level3[1255]),
   .I0(level4_in[7530]),
   .I1(level4_in[7531]),
   .I2(level4_in[7532]),
   .I3(level4_in[7533]),
   .I4(level4_in[7534]),
   .I5(level4_in[7535])
);

LUT6 #(
   .INIT(64'h97e8b88d97e8b88d)  
) LUT6_inst9032 (
   .O(to_level3[1256]),
   .I0(level4_in[7536]),
   .I1(level4_in[7537]),
   .I2(level4_in[7538]),
   .I3(level4_in[7539]),
   .I4(level4_in[7540]),
   .I5(level4_in[7541])
);

LUT6 #(
   .INIT(64'hfa2e4e8cfa2e4e8c)  
) LUT6_inst9033 (
   .O(to_level3[1257]),
   .I0(level4_in[7542]),
   .I1(level4_in[7543]),
   .I2(level4_in[7544]),
   .I3(level4_in[7545]),
   .I4(level4_in[7546]),
   .I5(level4_in[7547])
);

LUT6 #(
   .INIT(64'h185b4da2185b4da2)  
) LUT6_inst9034 (
   .O(to_level3[1258]),
   .I0(level4_in[7548]),
   .I1(level4_in[7549]),
   .I2(level4_in[7550]),
   .I3(level4_in[7551]),
   .I4(level4_in[7552]),
   .I5(level4_in[7553])
);

LUT6 #(
   .INIT(64'h5200166152001661)  
) LUT6_inst9035 (
   .O(to_level3[1259]),
   .I0(level4_in[7554]),
   .I1(level4_in[7555]),
   .I2(level4_in[7556]),
   .I3(level4_in[7557]),
   .I4(level4_in[7558]),
   .I5(level4_in[7559])
);

LUT6 #(
   .INIT(64'hf2435756f2435756)  
) LUT6_inst9036 (
   .O(to_level3[1260]),
   .I0(level4_in[7560]),
   .I1(level4_in[7561]),
   .I2(level4_in[7562]),
   .I3(level4_in[7563]),
   .I4(level4_in[7564]),
   .I5(level4_in[7565])
);

LUT6 #(
   .INIT(64'hee2285d9ee2285d9)  
) LUT6_inst9037 (
   .O(to_level3[1261]),
   .I0(level4_in[7566]),
   .I1(level4_in[7567]),
   .I2(level4_in[7568]),
   .I3(level4_in[7569]),
   .I4(level4_in[7570]),
   .I5(level4_in[7571])
);

LUT6 #(
   .INIT(64'h21e1ebb321e1ebb3)  
) LUT6_inst9038 (
   .O(to_level3[1262]),
   .I0(level4_in[7572]),
   .I1(level4_in[7573]),
   .I2(level4_in[7574]),
   .I3(level4_in[7575]),
   .I4(level4_in[7576]),
   .I5(level4_in[7577])
);

LUT6 #(
   .INIT(64'hc292a3f1c292a3f1)  
) LUT6_inst9039 (
   .O(to_level3[1263]),
   .I0(level4_in[7578]),
   .I1(level4_in[7579]),
   .I2(level4_in[7580]),
   .I3(level4_in[7581]),
   .I4(level4_in[7582]),
   .I5(level4_in[7583])
);

LUT6 #(
   .INIT(64'h419503f9419503f9)  
) LUT6_inst9040 (
   .O(to_level3[1264]),
   .I0(level4_in[7584]),
   .I1(level4_in[7585]),
   .I2(level4_in[7586]),
   .I3(level4_in[7587]),
   .I4(level4_in[7588]),
   .I5(level4_in[7589])
);

LUT6 #(
   .INIT(64'h4474860744748607)  
) LUT6_inst9041 (
   .O(to_level3[1265]),
   .I0(level4_in[7590]),
   .I1(level4_in[7591]),
   .I2(level4_in[7592]),
   .I3(level4_in[7593]),
   .I4(level4_in[7594]),
   .I5(level4_in[7595])
);

LUT6 #(
   .INIT(64'hc5de4734c5de4734)  
) LUT6_inst9042 (
   .O(to_level3[1266]),
   .I0(level4_in[7596]),
   .I1(level4_in[7597]),
   .I2(level4_in[7598]),
   .I3(level4_in[7599]),
   .I4(level4_in[7600]),
   .I5(level4_in[7601])
);

LUT6 #(
   .INIT(64'h284dd625284dd625)  
) LUT6_inst9043 (
   .O(to_level3[1267]),
   .I0(level4_in[7602]),
   .I1(level4_in[7603]),
   .I2(level4_in[7604]),
   .I3(level4_in[7605]),
   .I4(level4_in[7606]),
   .I5(level4_in[7607])
);

LUT6 #(
   .INIT(64'hf69b8bd9f69b8bd9)  
) LUT6_inst9044 (
   .O(to_level3[1268]),
   .I0(level4_in[7608]),
   .I1(level4_in[7609]),
   .I2(level4_in[7610]),
   .I3(level4_in[7611]),
   .I4(level4_in[7612]),
   .I5(level4_in[7613])
);

LUT6 #(
   .INIT(64'hbbfc7cdabbfc7cda)  
) LUT6_inst9045 (
   .O(to_level3[1269]),
   .I0(level4_in[7614]),
   .I1(level4_in[7615]),
   .I2(level4_in[7616]),
   .I3(level4_in[7617]),
   .I4(level4_in[7618]),
   .I5(level4_in[7619])
);

LUT6 #(
   .INIT(64'h3862556f3862556f)  
) LUT6_inst9046 (
   .O(to_level3[1270]),
   .I0(level4_in[7620]),
   .I1(level4_in[7621]),
   .I2(level4_in[7622]),
   .I3(level4_in[7623]),
   .I4(level4_in[7624]),
   .I5(level4_in[7625])
);

LUT6 #(
   .INIT(64'hce1377d3ce1377d3)  
) LUT6_inst9047 (
   .O(to_level3[1271]),
   .I0(level4_in[7626]),
   .I1(level4_in[7627]),
   .I2(level4_in[7628]),
   .I3(level4_in[7629]),
   .I4(level4_in[7630]),
   .I5(level4_in[7631])
);

LUT6 #(
   .INIT(64'h384bfae9384bfae9)  
) LUT6_inst9048 (
   .O(to_level3[1272]),
   .I0(level4_in[7632]),
   .I1(level4_in[7633]),
   .I2(level4_in[7634]),
   .I3(level4_in[7635]),
   .I4(level4_in[7636]),
   .I5(level4_in[7637])
);

LUT6 #(
   .INIT(64'hebd61a88ebd61a88)  
) LUT6_inst9049 (
   .O(to_level3[1273]),
   .I0(level4_in[7638]),
   .I1(level4_in[7639]),
   .I2(level4_in[7640]),
   .I3(level4_in[7641]),
   .I4(level4_in[7642]),
   .I5(level4_in[7643])
);

LUT6 #(
   .INIT(64'hc3397801c3397801)  
) LUT6_inst9050 (
   .O(to_level3[1274]),
   .I0(level4_in[7644]),
   .I1(level4_in[7645]),
   .I2(level4_in[7646]),
   .I3(level4_in[7647]),
   .I4(level4_in[7648]),
   .I5(level4_in[7649])
);

LUT6 #(
   .INIT(64'h954ff7b1954ff7b1)  
) LUT6_inst9051 (
   .O(to_level3[1275]),
   .I0(level4_in[7650]),
   .I1(level4_in[7651]),
   .I2(level4_in[7652]),
   .I3(level4_in[7653]),
   .I4(level4_in[7654]),
   .I5(level4_in[7655])
);

LUT6 #(
   .INIT(64'h42d4fbfe42d4fbfe)  
) LUT6_inst9052 (
   .O(to_level3[1276]),
   .I0(level4_in[7656]),
   .I1(level4_in[7657]),
   .I2(level4_in[7658]),
   .I3(level4_in[7659]),
   .I4(level4_in[7660]),
   .I5(level4_in[7661])
);

LUT6 #(
   .INIT(64'h5d6a63065d6a6306)  
) LUT6_inst9053 (
   .O(to_level3[1277]),
   .I0(level4_in[7662]),
   .I1(level4_in[7663]),
   .I2(level4_in[7664]),
   .I3(level4_in[7665]),
   .I4(level4_in[7666]),
   .I5(level4_in[7667])
);

LUT6 #(
   .INIT(64'h93f58eb493f58eb4)  
) LUT6_inst9054 (
   .O(to_level3[1278]),
   .I0(level4_in[7668]),
   .I1(level4_in[7669]),
   .I2(level4_in[7670]),
   .I3(level4_in[7671]),
   .I4(level4_in[7672]),
   .I5(level4_in[7673])
);

LUT6 #(
   .INIT(64'ha13127f4a13127f4)  
) LUT6_inst9055 (
   .O(to_level3[1279]),
   .I0(level4_in[7674]),
   .I1(level4_in[7675]),
   .I2(level4_in[7676]),
   .I3(level4_in[7677]),
   .I4(level4_in[7678]),
   .I5(level4_in[7679])
);

LUT6 #(
   .INIT(64'h347c703a347c703a)  
) LUT6_inst9056 (
   .O(to_level3[1280]),
   .I0(level4_in[7680]),
   .I1(level4_in[7681]),
   .I2(level4_in[7682]),
   .I3(level4_in[7683]),
   .I4(level4_in[7684]),
   .I5(level4_in[7685])
);

LUT6 #(
   .INIT(64'h7206d50b7206d50b)  
) LUT6_inst9057 (
   .O(to_level3[1281]),
   .I0(level4_in[7686]),
   .I1(level4_in[7687]),
   .I2(level4_in[7688]),
   .I3(level4_in[7689]),
   .I4(level4_in[7690]),
   .I5(level4_in[7691])
);

LUT6 #(
   .INIT(64'h9b7092869b709286)  
) LUT6_inst9058 (
   .O(to_level3[1282]),
   .I0(level4_in[7692]),
   .I1(level4_in[7693]),
   .I2(level4_in[7694]),
   .I3(level4_in[7695]),
   .I4(level4_in[7696]),
   .I5(level4_in[7697])
);

LUT6 #(
   .INIT(64'hed6704a4ed6704a4)  
) LUT6_inst9059 (
   .O(to_level3[1283]),
   .I0(level4_in[7698]),
   .I1(level4_in[7699]),
   .I2(level4_in[7700]),
   .I3(level4_in[7701]),
   .I4(level4_in[7702]),
   .I5(level4_in[7703])
);

LUT6 #(
   .INIT(64'h0292fdb40292fdb4)  
) LUT6_inst9060 (
   .O(to_level3[1284]),
   .I0(level4_in[7704]),
   .I1(level4_in[7705]),
   .I2(level4_in[7706]),
   .I3(level4_in[7707]),
   .I4(level4_in[7708]),
   .I5(level4_in[7709])
);

LUT6 #(
   .INIT(64'hab514abeab514abe)  
) LUT6_inst9061 (
   .O(to_level3[1285]),
   .I0(level4_in[7710]),
   .I1(level4_in[7711]),
   .I2(level4_in[7712]),
   .I3(level4_in[7713]),
   .I4(level4_in[7714]),
   .I5(level4_in[7715])
);

LUT6 #(
   .INIT(64'hd1ce4d44d1ce4d44)  
) LUT6_inst9062 (
   .O(to_level3[1286]),
   .I0(level4_in[7716]),
   .I1(level4_in[7717]),
   .I2(level4_in[7718]),
   .I3(level4_in[7719]),
   .I4(level4_in[7720]),
   .I5(level4_in[7721])
);

LUT6 #(
   .INIT(64'h0573554805735548)  
) LUT6_inst9063 (
   .O(to_level3[1287]),
   .I0(level4_in[7722]),
   .I1(level4_in[7723]),
   .I2(level4_in[7724]),
   .I3(level4_in[7725]),
   .I4(level4_in[7726]),
   .I5(level4_in[7727])
);

LUT6 #(
   .INIT(64'ha6df1e01a6df1e01)  
) LUT6_inst9064 (
   .O(to_level3[1288]),
   .I0(level4_in[7728]),
   .I1(level4_in[7729]),
   .I2(level4_in[7730]),
   .I3(level4_in[7731]),
   .I4(level4_in[7732]),
   .I5(level4_in[7733])
);

LUT6 #(
   .INIT(64'h111c0907111c0907)  
) LUT6_inst9065 (
   .O(to_level3[1289]),
   .I0(level4_in[7734]),
   .I1(level4_in[7735]),
   .I2(level4_in[7736]),
   .I3(level4_in[7737]),
   .I4(level4_in[7738]),
   .I5(level4_in[7739])
);

LUT6 #(
   .INIT(64'h211c937b211c937b)  
) LUT6_inst9066 (
   .O(to_level3[1290]),
   .I0(level4_in[7740]),
   .I1(level4_in[7741]),
   .I2(level4_in[7742]),
   .I3(level4_in[7743]),
   .I4(level4_in[7744]),
   .I5(level4_in[7745])
);

LUT6 #(
   .INIT(64'hcc42e236cc42e236)  
) LUT6_inst9067 (
   .O(to_level3[1291]),
   .I0(level4_in[7746]),
   .I1(level4_in[7747]),
   .I2(level4_in[7748]),
   .I3(level4_in[7749]),
   .I4(level4_in[7750]),
   .I5(level4_in[7751])
);

LUT6 #(
   .INIT(64'hcce22f96cce22f96)  
) LUT6_inst9068 (
   .O(to_level3[1292]),
   .I0(level4_in[7752]),
   .I1(level4_in[7753]),
   .I2(level4_in[7754]),
   .I3(level4_in[7755]),
   .I4(level4_in[7756]),
   .I5(level4_in[7757])
);

LUT6 #(
   .INIT(64'h022ec5ad022ec5ad)  
) LUT6_inst9069 (
   .O(to_level3[1293]),
   .I0(level4_in[7758]),
   .I1(level4_in[7759]),
   .I2(level4_in[7760]),
   .I3(level4_in[7761]),
   .I4(level4_in[7762]),
   .I5(level4_in[7763])
);

LUT6 #(
   .INIT(64'h49adf33a49adf33a)  
) LUT6_inst9070 (
   .O(to_level3[1294]),
   .I0(level4_in[7764]),
   .I1(level4_in[7765]),
   .I2(level4_in[7766]),
   .I3(level4_in[7767]),
   .I4(level4_in[7768]),
   .I5(level4_in[7769])
);

LUT6 #(
   .INIT(64'hd9d82a39d9d82a39)  
) LUT6_inst9071 (
   .O(to_level3[1295]),
   .I0(level4_in[7770]),
   .I1(level4_in[7771]),
   .I2(level4_in[7772]),
   .I3(level4_in[7773]),
   .I4(level4_in[7774]),
   .I5(level4_in[7775])
);
////////////// level 3 starts below:/n
LUT6 #(
   .INIT(64'h37c4b52937c4b529)  
) LUT6_inst9072 (
   .O(to_level2[0]),
   .I0(level3_in[0]),
   .I1(level3_in[1]),
   .I2(level3_in[2]),
   .I3(level3_in[3]),
   .I4(level3_in[4]),
   .I5(level3_in[5])
);

LUT6 #(
   .INIT(64'h7caa70b97caa70b9)  
) LUT6_inst9073 (
   .O(to_level2[1]),
   .I0(level3_in[6]),
   .I1(level3_in[7]),
   .I2(level3_in[8]),
   .I3(level3_in[9]),
   .I4(level3_in[10]),
   .I5(level3_in[11])
);

LUT6 #(
   .INIT(64'hef0f2b4fef0f2b4f)  
) LUT6_inst9074 (
   .O(to_level2[2]),
   .I0(level3_in[12]),
   .I1(level3_in[13]),
   .I2(level3_in[14]),
   .I3(level3_in[15]),
   .I4(level3_in[16]),
   .I5(level3_in[17])
);

LUT6 #(
   .INIT(64'h9642ed089642ed08)  
) LUT6_inst9075 (
   .O(to_level2[3]),
   .I0(level3_in[18]),
   .I1(level3_in[19]),
   .I2(level3_in[20]),
   .I3(level3_in[21]),
   .I4(level3_in[22]),
   .I5(level3_in[23])
);

LUT6 #(
   .INIT(64'h9d76c5829d76c582)  
) LUT6_inst9076 (
   .O(to_level2[4]),
   .I0(level3_in[24]),
   .I1(level3_in[25]),
   .I2(level3_in[26]),
   .I3(level3_in[27]),
   .I4(level3_in[28]),
   .I5(level3_in[29])
);

LUT6 #(
   .INIT(64'h57c7c52457c7c524)  
) LUT6_inst9077 (
   .O(to_level2[5]),
   .I0(level3_in[30]),
   .I1(level3_in[31]),
   .I2(level3_in[32]),
   .I3(level3_in[33]),
   .I4(level3_in[34]),
   .I5(level3_in[35])
);

LUT6 #(
   .INIT(64'h9ab776199ab77619)  
) LUT6_inst9078 (
   .O(to_level2[6]),
   .I0(level3_in[36]),
   .I1(level3_in[37]),
   .I2(level3_in[38]),
   .I3(level3_in[39]),
   .I4(level3_in[40]),
   .I5(level3_in[41])
);

LUT6 #(
   .INIT(64'h84e655bc84e655bc)  
) LUT6_inst9079 (
   .O(to_level2[7]),
   .I0(level3_in[42]),
   .I1(level3_in[43]),
   .I2(level3_in[44]),
   .I3(level3_in[45]),
   .I4(level3_in[46]),
   .I5(level3_in[47])
);

LUT6 #(
   .INIT(64'h5823dfd85823dfd8)  
) LUT6_inst9080 (
   .O(to_level2[8]),
   .I0(level3_in[48]),
   .I1(level3_in[49]),
   .I2(level3_in[50]),
   .I3(level3_in[51]),
   .I4(level3_in[52]),
   .I5(level3_in[53])
);

LUT6 #(
   .INIT(64'h9df97d879df97d87)  
) LUT6_inst9081 (
   .O(to_level2[9]),
   .I0(level3_in[54]),
   .I1(level3_in[55]),
   .I2(level3_in[56]),
   .I3(level3_in[57]),
   .I4(level3_in[58]),
   .I5(level3_in[59])
);

LUT6 #(
   .INIT(64'hb9a469d8b9a469d8)  
) LUT6_inst9082 (
   .O(to_level2[10]),
   .I0(level3_in[60]),
   .I1(level3_in[61]),
   .I2(level3_in[62]),
   .I3(level3_in[63]),
   .I4(level3_in[64]),
   .I5(level3_in[65])
);

LUT6 #(
   .INIT(64'hf722194ff722194f)  
) LUT6_inst9083 (
   .O(to_level2[11]),
   .I0(level3_in[66]),
   .I1(level3_in[67]),
   .I2(level3_in[68]),
   .I3(level3_in[69]),
   .I4(level3_in[70]),
   .I5(level3_in[71])
);

LUT6 #(
   .INIT(64'hf93c9e03f93c9e03)  
) LUT6_inst9084 (
   .O(to_level2[12]),
   .I0(level3_in[72]),
   .I1(level3_in[73]),
   .I2(level3_in[74]),
   .I3(level3_in[75]),
   .I4(level3_in[76]),
   .I5(level3_in[77])
);

LUT6 #(
   .INIT(64'h0aa8de1c0aa8de1c)  
) LUT6_inst9085 (
   .O(to_level2[13]),
   .I0(level3_in[78]),
   .I1(level3_in[79]),
   .I2(level3_in[80]),
   .I3(level3_in[81]),
   .I4(level3_in[82]),
   .I5(level3_in[83])
);

LUT6 #(
   .INIT(64'hdbbc061cdbbc061c)  
) LUT6_inst9086 (
   .O(to_level2[14]),
   .I0(level3_in[84]),
   .I1(level3_in[85]),
   .I2(level3_in[86]),
   .I3(level3_in[87]),
   .I4(level3_in[88]),
   .I5(level3_in[89])
);

LUT6 #(
   .INIT(64'h27ad0e2c27ad0e2c)  
) LUT6_inst9087 (
   .O(to_level2[15]),
   .I0(level3_in[90]),
   .I1(level3_in[91]),
   .I2(level3_in[92]),
   .I3(level3_in[93]),
   .I4(level3_in[94]),
   .I5(level3_in[95])
);

LUT6 #(
   .INIT(64'hc23d6cbac23d6cba)  
) LUT6_inst9088 (
   .O(to_level2[16]),
   .I0(level3_in[96]),
   .I1(level3_in[97]),
   .I2(level3_in[98]),
   .I3(level3_in[99]),
   .I4(level3_in[100]),
   .I5(level3_in[101])
);

LUT6 #(
   .INIT(64'h348aba9e348aba9e)  
) LUT6_inst9089 (
   .O(to_level2[17]),
   .I0(level3_in[102]),
   .I1(level3_in[103]),
   .I2(level3_in[104]),
   .I3(level3_in[105]),
   .I4(level3_in[106]),
   .I5(level3_in[107])
);

LUT6 #(
   .INIT(64'h290ddd75290ddd75)  
) LUT6_inst9090 (
   .O(to_level2[18]),
   .I0(level3_in[108]),
   .I1(level3_in[109]),
   .I2(level3_in[110]),
   .I3(level3_in[111]),
   .I4(level3_in[112]),
   .I5(level3_in[113])
);

LUT6 #(
   .INIT(64'h4326b4ad4326b4ad)  
) LUT6_inst9091 (
   .O(to_level2[19]),
   .I0(level3_in[114]),
   .I1(level3_in[115]),
   .I2(level3_in[116]),
   .I3(level3_in[117]),
   .I4(level3_in[118]),
   .I5(level3_in[119])
);

LUT6 #(
   .INIT(64'h0dd8df180dd8df18)  
) LUT6_inst9092 (
   .O(to_level2[20]),
   .I0(level3_in[120]),
   .I1(level3_in[121]),
   .I2(level3_in[122]),
   .I3(level3_in[123]),
   .I4(level3_in[124]),
   .I5(level3_in[125])
);

LUT6 #(
   .INIT(64'hd08710a8d08710a8)  
) LUT6_inst9093 (
   .O(to_level2[21]),
   .I0(level3_in[126]),
   .I1(level3_in[127]),
   .I2(level3_in[128]),
   .I3(level3_in[129]),
   .I4(level3_in[130]),
   .I5(level3_in[131])
);

LUT6 #(
   .INIT(64'hdbd09ad4dbd09ad4)  
) LUT6_inst9094 (
   .O(to_level2[22]),
   .I0(level3_in[132]),
   .I1(level3_in[133]),
   .I2(level3_in[134]),
   .I3(level3_in[135]),
   .I4(level3_in[136]),
   .I5(level3_in[137])
);

LUT6 #(
   .INIT(64'h4a85e77d4a85e77d)  
) LUT6_inst9095 (
   .O(to_level2[23]),
   .I0(level3_in[138]),
   .I1(level3_in[139]),
   .I2(level3_in[140]),
   .I3(level3_in[141]),
   .I4(level3_in[142]),
   .I5(level3_in[143])
);

LUT6 #(
   .INIT(64'he6d9e715e6d9e715)  
) LUT6_inst9096 (
   .O(to_level2[24]),
   .I0(level3_in[144]),
   .I1(level3_in[145]),
   .I2(level3_in[146]),
   .I3(level3_in[147]),
   .I4(level3_in[148]),
   .I5(level3_in[149])
);

LUT6 #(
   .INIT(64'h6c968a656c968a65)  
) LUT6_inst9097 (
   .O(to_level2[25]),
   .I0(level3_in[150]),
   .I1(level3_in[151]),
   .I2(level3_in[152]),
   .I3(level3_in[153]),
   .I4(level3_in[154]),
   .I5(level3_in[155])
);

LUT6 #(
   .INIT(64'h028495fb028495fb)  
) LUT6_inst9098 (
   .O(to_level2[26]),
   .I0(level3_in[156]),
   .I1(level3_in[157]),
   .I2(level3_in[158]),
   .I3(level3_in[159]),
   .I4(level3_in[160]),
   .I5(level3_in[161])
);

LUT6 #(
   .INIT(64'h2509c1482509c148)  
) LUT6_inst9099 (
   .O(to_level2[27]),
   .I0(level3_in[162]),
   .I1(level3_in[163]),
   .I2(level3_in[164]),
   .I3(level3_in[165]),
   .I4(level3_in[166]),
   .I5(level3_in[167])
);

LUT6 #(
   .INIT(64'h5e55253a5e55253a)  
) LUT6_inst9100 (
   .O(to_level2[28]),
   .I0(level3_in[168]),
   .I1(level3_in[169]),
   .I2(level3_in[170]),
   .I3(level3_in[171]),
   .I4(level3_in[172]),
   .I5(level3_in[173])
);

LUT6 #(
   .INIT(64'h47e1f0b047e1f0b0)  
) LUT6_inst9101 (
   .O(to_level2[29]),
   .I0(level3_in[174]),
   .I1(level3_in[175]),
   .I2(level3_in[176]),
   .I3(level3_in[177]),
   .I4(level3_in[178]),
   .I5(level3_in[179])
);

LUT6 #(
   .INIT(64'hb0c2725db0c2725d)  
) LUT6_inst9102 (
   .O(to_level2[30]),
   .I0(level3_in[180]),
   .I1(level3_in[181]),
   .I2(level3_in[182]),
   .I3(level3_in[183]),
   .I4(level3_in[184]),
   .I5(level3_in[185])
);

LUT6 #(
   .INIT(64'hcdbc082bcdbc082b)  
) LUT6_inst9103 (
   .O(to_level2[31]),
   .I0(level3_in[186]),
   .I1(level3_in[187]),
   .I2(level3_in[188]),
   .I3(level3_in[189]),
   .I4(level3_in[190]),
   .I5(level3_in[191])
);

LUT6 #(
   .INIT(64'h6c6961b36c6961b3)  
) LUT6_inst9104 (
   .O(to_level2[32]),
   .I0(level3_in[192]),
   .I1(level3_in[193]),
   .I2(level3_in[194]),
   .I3(level3_in[195]),
   .I4(level3_in[196]),
   .I5(level3_in[197])
);

LUT6 #(
   .INIT(64'hd6ceb708d6ceb708)  
) LUT6_inst9105 (
   .O(to_level2[33]),
   .I0(level3_in[198]),
   .I1(level3_in[199]),
   .I2(level3_in[200]),
   .I3(level3_in[201]),
   .I4(level3_in[202]),
   .I5(level3_in[203])
);

LUT6 #(
   .INIT(64'hcf2b43dbcf2b43db)  
) LUT6_inst9106 (
   .O(to_level2[34]),
   .I0(level3_in[204]),
   .I1(level3_in[205]),
   .I2(level3_in[206]),
   .I3(level3_in[207]),
   .I4(level3_in[208]),
   .I5(level3_in[209])
);

LUT6 #(
   .INIT(64'he20ebee1e20ebee1)  
) LUT6_inst9107 (
   .O(to_level2[35]),
   .I0(level3_in[210]),
   .I1(level3_in[211]),
   .I2(level3_in[212]),
   .I3(level3_in[213]),
   .I4(level3_in[214]),
   .I5(level3_in[215])
);

LUT6 #(
   .INIT(64'hf959d56bf959d56b)  
) LUT6_inst9108 (
   .O(to_level2[36]),
   .I0(level3_in[216]),
   .I1(level3_in[217]),
   .I2(level3_in[218]),
   .I3(level3_in[219]),
   .I4(level3_in[220]),
   .I5(level3_in[221])
);

LUT6 #(
   .INIT(64'h34ab8e8834ab8e88)  
) LUT6_inst9109 (
   .O(to_level2[37]),
   .I0(level3_in[222]),
   .I1(level3_in[223]),
   .I2(level3_in[224]),
   .I3(level3_in[225]),
   .I4(level3_in[226]),
   .I5(level3_in[227])
);

LUT6 #(
   .INIT(64'h2ab876492ab87649)  
) LUT6_inst9110 (
   .O(to_level2[38]),
   .I0(level3_in[228]),
   .I1(level3_in[229]),
   .I2(level3_in[230]),
   .I3(level3_in[231]),
   .I4(level3_in[232]),
   .I5(level3_in[233])
);

LUT6 #(
   .INIT(64'h479a2109479a2109)  
) LUT6_inst9111 (
   .O(to_level2[39]),
   .I0(level3_in[234]),
   .I1(level3_in[235]),
   .I2(level3_in[236]),
   .I3(level3_in[237]),
   .I4(level3_in[238]),
   .I5(level3_in[239])
);

LUT6 #(
   .INIT(64'hc6a333ccc6a333cc)  
) LUT6_inst9112 (
   .O(to_level2[40]),
   .I0(level3_in[240]),
   .I1(level3_in[241]),
   .I2(level3_in[242]),
   .I3(level3_in[243]),
   .I4(level3_in[244]),
   .I5(level3_in[245])
);

LUT6 #(
   .INIT(64'h8e3d930d8e3d930d)  
) LUT6_inst9113 (
   .O(to_level2[41]),
   .I0(level3_in[246]),
   .I1(level3_in[247]),
   .I2(level3_in[248]),
   .I3(level3_in[249]),
   .I4(level3_in[250]),
   .I5(level3_in[251])
);

LUT6 #(
   .INIT(64'h736cf3eb736cf3eb)  
) LUT6_inst9114 (
   .O(to_level2[42]),
   .I0(level3_in[252]),
   .I1(level3_in[253]),
   .I2(level3_in[254]),
   .I3(level3_in[255]),
   .I4(level3_in[256]),
   .I5(level3_in[257])
);

LUT6 #(
   .INIT(64'h55f05daf55f05daf)  
) LUT6_inst9115 (
   .O(to_level2[43]),
   .I0(level3_in[258]),
   .I1(level3_in[259]),
   .I2(level3_in[260]),
   .I3(level3_in[261]),
   .I4(level3_in[262]),
   .I5(level3_in[263])
);

LUT6 #(
   .INIT(64'h74fe8d1274fe8d12)  
) LUT6_inst9116 (
   .O(to_level2[44]),
   .I0(level3_in[264]),
   .I1(level3_in[265]),
   .I2(level3_in[266]),
   .I3(level3_in[267]),
   .I4(level3_in[268]),
   .I5(level3_in[269])
);

LUT6 #(
   .INIT(64'he6326fe7e6326fe7)  
) LUT6_inst9117 (
   .O(to_level2[45]),
   .I0(level3_in[270]),
   .I1(level3_in[271]),
   .I2(level3_in[272]),
   .I3(level3_in[273]),
   .I4(level3_in[274]),
   .I5(level3_in[275])
);

LUT6 #(
   .INIT(64'h6f61f3b46f61f3b4)  
) LUT6_inst9118 (
   .O(to_level2[46]),
   .I0(level3_in[276]),
   .I1(level3_in[277]),
   .I2(level3_in[278]),
   .I3(level3_in[279]),
   .I4(level3_in[280]),
   .I5(level3_in[281])
);

LUT6 #(
   .INIT(64'ha82d6a93a82d6a93)  
) LUT6_inst9119 (
   .O(to_level2[47]),
   .I0(level3_in[282]),
   .I1(level3_in[283]),
   .I2(level3_in[284]),
   .I3(level3_in[285]),
   .I4(level3_in[286]),
   .I5(level3_in[287])
);

LUT6 #(
   .INIT(64'hacf86f1aacf86f1a)  
) LUT6_inst9120 (
   .O(to_level2[48]),
   .I0(level3_in[288]),
   .I1(level3_in[289]),
   .I2(level3_in[290]),
   .I3(level3_in[291]),
   .I4(level3_in[292]),
   .I5(level3_in[293])
);

LUT6 #(
   .INIT(64'h3482d9633482d963)  
) LUT6_inst9121 (
   .O(to_level2[49]),
   .I0(level3_in[294]),
   .I1(level3_in[295]),
   .I2(level3_in[296]),
   .I3(level3_in[297]),
   .I4(level3_in[298]),
   .I5(level3_in[299])
);

LUT6 #(
   .INIT(64'h791a4979791a4979)  
) LUT6_inst9122 (
   .O(to_level2[50]),
   .I0(level3_in[300]),
   .I1(level3_in[301]),
   .I2(level3_in[302]),
   .I3(level3_in[303]),
   .I4(level3_in[304]),
   .I5(level3_in[305])
);

LUT6 #(
   .INIT(64'h92231d3292231d32)  
) LUT6_inst9123 (
   .O(to_level2[51]),
   .I0(level3_in[306]),
   .I1(level3_in[307]),
   .I2(level3_in[308]),
   .I3(level3_in[309]),
   .I4(level3_in[310]),
   .I5(level3_in[311])
);

LUT6 #(
   .INIT(64'hdaaa9240daaa9240)  
) LUT6_inst9124 (
   .O(to_level2[52]),
   .I0(level3_in[312]),
   .I1(level3_in[313]),
   .I2(level3_in[314]),
   .I3(level3_in[315]),
   .I4(level3_in[316]),
   .I5(level3_in[317])
);

LUT6 #(
   .INIT(64'h535b7320535b7320)  
) LUT6_inst9125 (
   .O(to_level2[53]),
   .I0(level3_in[318]),
   .I1(level3_in[319]),
   .I2(level3_in[320]),
   .I3(level3_in[321]),
   .I4(level3_in[322]),
   .I5(level3_in[323])
);

LUT6 #(
   .INIT(64'h1f02d35f1f02d35f)  
) LUT6_inst9126 (
   .O(to_level2[54]),
   .I0(level3_in[324]),
   .I1(level3_in[325]),
   .I2(level3_in[326]),
   .I3(level3_in[327]),
   .I4(level3_in[328]),
   .I5(level3_in[329])
);

LUT6 #(
   .INIT(64'h891d75bc891d75bc)  
) LUT6_inst9127 (
   .O(to_level2[55]),
   .I0(level3_in[330]),
   .I1(level3_in[331]),
   .I2(level3_in[332]),
   .I3(level3_in[333]),
   .I4(level3_in[334]),
   .I5(level3_in[335])
);

LUT6 #(
   .INIT(64'h7f216ed27f216ed2)  
) LUT6_inst9128 (
   .O(to_level2[56]),
   .I0(level3_in[336]),
   .I1(level3_in[337]),
   .I2(level3_in[338]),
   .I3(level3_in[339]),
   .I4(level3_in[340]),
   .I5(level3_in[341])
);

LUT6 #(
   .INIT(64'h03e7dcbe03e7dcbe)  
) LUT6_inst9129 (
   .O(to_level2[57]),
   .I0(level3_in[342]),
   .I1(level3_in[343]),
   .I2(level3_in[344]),
   .I3(level3_in[345]),
   .I4(level3_in[346]),
   .I5(level3_in[347])
);

LUT6 #(
   .INIT(64'ha4de4e6ca4de4e6c)  
) LUT6_inst9130 (
   .O(to_level2[58]),
   .I0(level3_in[348]),
   .I1(level3_in[349]),
   .I2(level3_in[350]),
   .I3(level3_in[351]),
   .I4(level3_in[352]),
   .I5(level3_in[353])
);

LUT6 #(
   .INIT(64'h8640e0c18640e0c1)  
) LUT6_inst9131 (
   .O(to_level2[59]),
   .I0(level3_in[354]),
   .I1(level3_in[355]),
   .I2(level3_in[356]),
   .I3(level3_in[357]),
   .I4(level3_in[358]),
   .I5(level3_in[359])
);

LUT6 #(
   .INIT(64'hc1a8937ec1a8937e)  
) LUT6_inst9132 (
   .O(to_level2[60]),
   .I0(level3_in[360]),
   .I1(level3_in[361]),
   .I2(level3_in[362]),
   .I3(level3_in[363]),
   .I4(level3_in[364]),
   .I5(level3_in[365])
);

LUT6 #(
   .INIT(64'hd8845f1dd8845f1d)  
) LUT6_inst9133 (
   .O(to_level2[61]),
   .I0(level3_in[366]),
   .I1(level3_in[367]),
   .I2(level3_in[368]),
   .I3(level3_in[369]),
   .I4(level3_in[370]),
   .I5(level3_in[371])
);

LUT6 #(
   .INIT(64'h704a6435704a6435)  
) LUT6_inst9134 (
   .O(to_level2[62]),
   .I0(level3_in[372]),
   .I1(level3_in[373]),
   .I2(level3_in[374]),
   .I3(level3_in[375]),
   .I4(level3_in[376]),
   .I5(level3_in[377])
);

LUT6 #(
   .INIT(64'hc93968d1c93968d1)  
) LUT6_inst9135 (
   .O(to_level2[63]),
   .I0(level3_in[378]),
   .I1(level3_in[379]),
   .I2(level3_in[380]),
   .I3(level3_in[381]),
   .I4(level3_in[382]),
   .I5(level3_in[383])
);

LUT6 #(
   .INIT(64'hf99e31b2f99e31b2)  
) LUT6_inst9136 (
   .O(to_level2[64]),
   .I0(level3_in[384]),
   .I1(level3_in[385]),
   .I2(level3_in[386]),
   .I3(level3_in[387]),
   .I4(level3_in[388]),
   .I5(level3_in[389])
);

LUT6 #(
   .INIT(64'h7ced551d7ced551d)  
) LUT6_inst9137 (
   .O(to_level2[65]),
   .I0(level3_in[390]),
   .I1(level3_in[391]),
   .I2(level3_in[392]),
   .I3(level3_in[393]),
   .I4(level3_in[394]),
   .I5(level3_in[395])
);

LUT6 #(
   .INIT(64'h9f7c98129f7c9812)  
) LUT6_inst9138 (
   .O(to_level2[66]),
   .I0(level3_in[396]),
   .I1(level3_in[397]),
   .I2(level3_in[398]),
   .I3(level3_in[399]),
   .I4(level3_in[400]),
   .I5(level3_in[401])
);

LUT6 #(
   .INIT(64'h549d34fc549d34fc)  
) LUT6_inst9139 (
   .O(to_level2[67]),
   .I0(level3_in[402]),
   .I1(level3_in[403]),
   .I2(level3_in[404]),
   .I3(level3_in[405]),
   .I4(level3_in[406]),
   .I5(level3_in[407])
);

LUT6 #(
   .INIT(64'h367cc3ad367cc3ad)  
) LUT6_inst9140 (
   .O(to_level2[68]),
   .I0(level3_in[408]),
   .I1(level3_in[409]),
   .I2(level3_in[410]),
   .I3(level3_in[411]),
   .I4(level3_in[412]),
   .I5(level3_in[413])
);

LUT6 #(
   .INIT(64'h5bb1020f5bb1020f)  
) LUT6_inst9141 (
   .O(to_level2[69]),
   .I0(level3_in[414]),
   .I1(level3_in[415]),
   .I2(level3_in[416]),
   .I3(level3_in[417]),
   .I4(level3_in[418]),
   .I5(level3_in[419])
);

LUT6 #(
   .INIT(64'h216f8efa216f8efa)  
) LUT6_inst9142 (
   .O(to_level2[70]),
   .I0(level3_in[420]),
   .I1(level3_in[421]),
   .I2(level3_in[422]),
   .I3(level3_in[423]),
   .I4(level3_in[424]),
   .I5(level3_in[425])
);

LUT6 #(
   .INIT(64'h0f3806e50f3806e5)  
) LUT6_inst9143 (
   .O(to_level2[71]),
   .I0(level3_in[426]),
   .I1(level3_in[427]),
   .I2(level3_in[428]),
   .I3(level3_in[429]),
   .I4(level3_in[430]),
   .I5(level3_in[431])
);

LUT6 #(
   .INIT(64'h8a05420e8a05420e)  
) LUT6_inst9144 (
   .O(to_level2[72]),
   .I0(level3_in[432]),
   .I1(level3_in[433]),
   .I2(level3_in[434]),
   .I3(level3_in[435]),
   .I4(level3_in[436]),
   .I5(level3_in[437])
);

LUT6 #(
   .INIT(64'hc9cda7f5c9cda7f5)  
) LUT6_inst9145 (
   .O(to_level2[73]),
   .I0(level3_in[438]),
   .I1(level3_in[439]),
   .I2(level3_in[440]),
   .I3(level3_in[441]),
   .I4(level3_in[442]),
   .I5(level3_in[443])
);

LUT6 #(
   .INIT(64'h1c8c42631c8c4263)  
) LUT6_inst9146 (
   .O(to_level2[74]),
   .I0(level3_in[444]),
   .I1(level3_in[445]),
   .I2(level3_in[446]),
   .I3(level3_in[447]),
   .I4(level3_in[448]),
   .I5(level3_in[449])
);

LUT6 #(
   .INIT(64'hc8f3dd0bc8f3dd0b)  
) LUT6_inst9147 (
   .O(to_level2[75]),
   .I0(level3_in[450]),
   .I1(level3_in[451]),
   .I2(level3_in[452]),
   .I3(level3_in[453]),
   .I4(level3_in[454]),
   .I5(level3_in[455])
);

LUT6 #(
   .INIT(64'hdd24f145dd24f145)  
) LUT6_inst9148 (
   .O(to_level2[76]),
   .I0(level3_in[456]),
   .I1(level3_in[457]),
   .I2(level3_in[458]),
   .I3(level3_in[459]),
   .I4(level3_in[460]),
   .I5(level3_in[461])
);

LUT6 #(
   .INIT(64'h2b2112a02b2112a0)  
) LUT6_inst9149 (
   .O(to_level2[77]),
   .I0(level3_in[462]),
   .I1(level3_in[463]),
   .I2(level3_in[464]),
   .I3(level3_in[465]),
   .I4(level3_in[466]),
   .I5(level3_in[467])
);

LUT6 #(
   .INIT(64'h591f8fa7591f8fa7)  
) LUT6_inst9150 (
   .O(to_level2[78]),
   .I0(level3_in[468]),
   .I1(level3_in[469]),
   .I2(level3_in[470]),
   .I3(level3_in[471]),
   .I4(level3_in[472]),
   .I5(level3_in[473])
);

LUT6 #(
   .INIT(64'h4dfa55534dfa5553)  
) LUT6_inst9151 (
   .O(to_level2[79]),
   .I0(level3_in[474]),
   .I1(level3_in[475]),
   .I2(level3_in[476]),
   .I3(level3_in[477]),
   .I4(level3_in[478]),
   .I5(level3_in[479])
);

LUT6 #(
   .INIT(64'hfbd98272fbd98272)  
) LUT6_inst9152 (
   .O(to_level2[80]),
   .I0(level3_in[480]),
   .I1(level3_in[481]),
   .I2(level3_in[482]),
   .I3(level3_in[483]),
   .I4(level3_in[484]),
   .I5(level3_in[485])
);

LUT6 #(
   .INIT(64'h9d187d739d187d73)  
) LUT6_inst9153 (
   .O(to_level2[81]),
   .I0(level3_in[486]),
   .I1(level3_in[487]),
   .I2(level3_in[488]),
   .I3(level3_in[489]),
   .I4(level3_in[490]),
   .I5(level3_in[491])
);

LUT6 #(
   .INIT(64'hb7e10eadb7e10ead)  
) LUT6_inst9154 (
   .O(to_level2[82]),
   .I0(level3_in[492]),
   .I1(level3_in[493]),
   .I2(level3_in[494]),
   .I3(level3_in[495]),
   .I4(level3_in[496]),
   .I5(level3_in[497])
);

LUT6 #(
   .INIT(64'h1696479e1696479e)  
) LUT6_inst9155 (
   .O(to_level2[83]),
   .I0(level3_in[498]),
   .I1(level3_in[499]),
   .I2(level3_in[500]),
   .I3(level3_in[501]),
   .I4(level3_in[502]),
   .I5(level3_in[503])
);

LUT6 #(
   .INIT(64'ha4424257a4424257)  
) LUT6_inst9156 (
   .O(to_level2[84]),
   .I0(level3_in[504]),
   .I1(level3_in[505]),
   .I2(level3_in[506]),
   .I3(level3_in[507]),
   .I4(level3_in[508]),
   .I5(level3_in[509])
);

LUT6 #(
   .INIT(64'h3de78e623de78e62)  
) LUT6_inst9157 (
   .O(to_level2[85]),
   .I0(level3_in[510]),
   .I1(level3_in[511]),
   .I2(level3_in[512]),
   .I3(level3_in[513]),
   .I4(level3_in[514]),
   .I5(level3_in[515])
);

LUT6 #(
   .INIT(64'hd78031ffd78031ff)  
) LUT6_inst9158 (
   .O(to_level2[86]),
   .I0(level3_in[516]),
   .I1(level3_in[517]),
   .I2(level3_in[518]),
   .I3(level3_in[519]),
   .I4(level3_in[520]),
   .I5(level3_in[521])
);

LUT6 #(
   .INIT(64'hea15170fea15170f)  
) LUT6_inst9159 (
   .O(to_level2[87]),
   .I0(level3_in[522]),
   .I1(level3_in[523]),
   .I2(level3_in[524]),
   .I3(level3_in[525]),
   .I4(level3_in[526]),
   .I5(level3_in[527])
);

LUT6 #(
   .INIT(64'h8dd19b548dd19b54)  
) LUT6_inst9160 (
   .O(to_level2[88]),
   .I0(level3_in[528]),
   .I1(level3_in[529]),
   .I2(level3_in[530]),
   .I3(level3_in[531]),
   .I4(level3_in[532]),
   .I5(level3_in[533])
);

LUT6 #(
   .INIT(64'hf008391ef008391e)  
) LUT6_inst9161 (
   .O(to_level2[89]),
   .I0(level3_in[534]),
   .I1(level3_in[535]),
   .I2(level3_in[536]),
   .I3(level3_in[537]),
   .I4(level3_in[538]),
   .I5(level3_in[539])
);

LUT6 #(
   .INIT(64'h4205d8c74205d8c7)  
) LUT6_inst9162 (
   .O(to_level2[90]),
   .I0(level3_in[540]),
   .I1(level3_in[541]),
   .I2(level3_in[542]),
   .I3(level3_in[543]),
   .I4(level3_in[544]),
   .I5(level3_in[545])
);

LUT6 #(
   .INIT(64'h193167cb193167cb)  
) LUT6_inst9163 (
   .O(to_level2[91]),
   .I0(level3_in[546]),
   .I1(level3_in[547]),
   .I2(level3_in[548]),
   .I3(level3_in[549]),
   .I4(level3_in[550]),
   .I5(level3_in[551])
);

LUT6 #(
   .INIT(64'h2ff3736b2ff3736b)  
) LUT6_inst9164 (
   .O(to_level2[92]),
   .I0(level3_in[552]),
   .I1(level3_in[553]),
   .I2(level3_in[554]),
   .I3(level3_in[555]),
   .I4(level3_in[556]),
   .I5(level3_in[557])
);

LUT6 #(
   .INIT(64'hdf31ecfddf31ecfd)  
) LUT6_inst9165 (
   .O(to_level2[93]),
   .I0(level3_in[558]),
   .I1(level3_in[559]),
   .I2(level3_in[560]),
   .I3(level3_in[561]),
   .I4(level3_in[562]),
   .I5(level3_in[563])
);

LUT6 #(
   .INIT(64'ha27001fea27001fe)  
) LUT6_inst9166 (
   .O(to_level2[94]),
   .I0(level3_in[564]),
   .I1(level3_in[565]),
   .I2(level3_in[566]),
   .I3(level3_in[567]),
   .I4(level3_in[568]),
   .I5(level3_in[569])
);

LUT6 #(
   .INIT(64'h0699647506996475)  
) LUT6_inst9167 (
   .O(to_level2[95]),
   .I0(level3_in[570]),
   .I1(level3_in[571]),
   .I2(level3_in[572]),
   .I3(level3_in[573]),
   .I4(level3_in[574]),
   .I5(level3_in[575])
);

LUT6 #(
   .INIT(64'h086c4e4f086c4e4f)  
) LUT6_inst9168 (
   .O(to_level2[96]),
   .I0(level3_in[576]),
   .I1(level3_in[577]),
   .I2(level3_in[578]),
   .I3(level3_in[579]),
   .I4(level3_in[580]),
   .I5(level3_in[581])
);

LUT6 #(
   .INIT(64'h963e85f3963e85f3)  
) LUT6_inst9169 (
   .O(to_level2[97]),
   .I0(level3_in[582]),
   .I1(level3_in[583]),
   .I2(level3_in[584]),
   .I3(level3_in[585]),
   .I4(level3_in[586]),
   .I5(level3_in[587])
);

LUT6 #(
   .INIT(64'h58fb551f58fb551f)  
) LUT6_inst9170 (
   .O(to_level2[98]),
   .I0(level3_in[588]),
   .I1(level3_in[589]),
   .I2(level3_in[590]),
   .I3(level3_in[591]),
   .I4(level3_in[592]),
   .I5(level3_in[593])
);

LUT6 #(
   .INIT(64'hf727a953f727a953)  
) LUT6_inst9171 (
   .O(to_level2[99]),
   .I0(level3_in[594]),
   .I1(level3_in[595]),
   .I2(level3_in[596]),
   .I3(level3_in[597]),
   .I4(level3_in[598]),
   .I5(level3_in[599])
);

LUT6 #(
   .INIT(64'h8cdbca538cdbca53)  
) LUT6_inst9172 (
   .O(to_level2[100]),
   .I0(level3_in[600]),
   .I1(level3_in[601]),
   .I2(level3_in[602]),
   .I3(level3_in[603]),
   .I4(level3_in[604]),
   .I5(level3_in[605])
);

LUT6 #(
   .INIT(64'hf7044bb5f7044bb5)  
) LUT6_inst9173 (
   .O(to_level2[101]),
   .I0(level3_in[606]),
   .I1(level3_in[607]),
   .I2(level3_in[608]),
   .I3(level3_in[609]),
   .I4(level3_in[610]),
   .I5(level3_in[611])
);

LUT6 #(
   .INIT(64'ha906b845a906b845)  
) LUT6_inst9174 (
   .O(to_level2[102]),
   .I0(level3_in[612]),
   .I1(level3_in[613]),
   .I2(level3_in[614]),
   .I3(level3_in[615]),
   .I4(level3_in[616]),
   .I5(level3_in[617])
);

LUT6 #(
   .INIT(64'h18fcfc7918fcfc79)  
) LUT6_inst9175 (
   .O(to_level2[103]),
   .I0(level3_in[618]),
   .I1(level3_in[619]),
   .I2(level3_in[620]),
   .I3(level3_in[621]),
   .I4(level3_in[622]),
   .I5(level3_in[623])
);

LUT6 #(
   .INIT(64'hdf441499df441499)  
) LUT6_inst9176 (
   .O(to_level2[104]),
   .I0(level3_in[624]),
   .I1(level3_in[625]),
   .I2(level3_in[626]),
   .I3(level3_in[627]),
   .I4(level3_in[628]),
   .I5(level3_in[629])
);

LUT6 #(
   .INIT(64'h88c2c39888c2c398)  
) LUT6_inst9177 (
   .O(to_level2[105]),
   .I0(level3_in[630]),
   .I1(level3_in[631]),
   .I2(level3_in[632]),
   .I3(level3_in[633]),
   .I4(level3_in[634]),
   .I5(level3_in[635])
);

LUT6 #(
   .INIT(64'hcd2c9e7bcd2c9e7b)  
) LUT6_inst9178 (
   .O(to_level2[106]),
   .I0(level3_in[636]),
   .I1(level3_in[637]),
   .I2(level3_in[638]),
   .I3(level3_in[639]),
   .I4(level3_in[640]),
   .I5(level3_in[641])
);

LUT6 #(
   .INIT(64'h7a23d27d7a23d27d)  
) LUT6_inst9179 (
   .O(to_level2[107]),
   .I0(level3_in[642]),
   .I1(level3_in[643]),
   .I2(level3_in[644]),
   .I3(level3_in[645]),
   .I4(level3_in[646]),
   .I5(level3_in[647])
);

LUT6 #(
   .INIT(64'h4ee7d5b64ee7d5b6)  
) LUT6_inst9180 (
   .O(to_level2[108]),
   .I0(level3_in[648]),
   .I1(level3_in[649]),
   .I2(level3_in[650]),
   .I3(level3_in[651]),
   .I4(level3_in[652]),
   .I5(level3_in[653])
);

LUT6 #(
   .INIT(64'he3be1072e3be1072)  
) LUT6_inst9181 (
   .O(to_level2[109]),
   .I0(level3_in[654]),
   .I1(level3_in[655]),
   .I2(level3_in[656]),
   .I3(level3_in[657]),
   .I4(level3_in[658]),
   .I5(level3_in[659])
);

LUT6 #(
   .INIT(64'he3ffb50fe3ffb50f)  
) LUT6_inst9182 (
   .O(to_level2[110]),
   .I0(level3_in[660]),
   .I1(level3_in[661]),
   .I2(level3_in[662]),
   .I3(level3_in[663]),
   .I4(level3_in[664]),
   .I5(level3_in[665])
);

LUT6 #(
   .INIT(64'h112ff996112ff996)  
) LUT6_inst9183 (
   .O(to_level2[111]),
   .I0(level3_in[666]),
   .I1(level3_in[667]),
   .I2(level3_in[668]),
   .I3(level3_in[669]),
   .I4(level3_in[670]),
   .I5(level3_in[671])
);

LUT6 #(
   .INIT(64'hc9e9000ec9e9000e)  
) LUT6_inst9184 (
   .O(to_level2[112]),
   .I0(level3_in[672]),
   .I1(level3_in[673]),
   .I2(level3_in[674]),
   .I3(level3_in[675]),
   .I4(level3_in[676]),
   .I5(level3_in[677])
);

LUT6 #(
   .INIT(64'h7757bff97757bff9)  
) LUT6_inst9185 (
   .O(to_level2[113]),
   .I0(level3_in[678]),
   .I1(level3_in[679]),
   .I2(level3_in[680]),
   .I3(level3_in[681]),
   .I4(level3_in[682]),
   .I5(level3_in[683])
);

LUT6 #(
   .INIT(64'h0b7b373c0b7b373c)  
) LUT6_inst9186 (
   .O(to_level2[114]),
   .I0(level3_in[684]),
   .I1(level3_in[685]),
   .I2(level3_in[686]),
   .I3(level3_in[687]),
   .I4(level3_in[688]),
   .I5(level3_in[689])
);

LUT6 #(
   .INIT(64'hd78a7dc9d78a7dc9)  
) LUT6_inst9187 (
   .O(to_level2[115]),
   .I0(level3_in[690]),
   .I1(level3_in[691]),
   .I2(level3_in[692]),
   .I3(level3_in[693]),
   .I4(level3_in[694]),
   .I5(level3_in[695])
);

LUT6 #(
   .INIT(64'h74ca077674ca0776)  
) LUT6_inst9188 (
   .O(to_level2[116]),
   .I0(level3_in[696]),
   .I1(level3_in[697]),
   .I2(level3_in[698]),
   .I3(level3_in[699]),
   .I4(level3_in[700]),
   .I5(level3_in[701])
);

LUT6 #(
   .INIT(64'h99447b6699447b66)  
) LUT6_inst9189 (
   .O(to_level2[117]),
   .I0(level3_in[702]),
   .I1(level3_in[703]),
   .I2(level3_in[704]),
   .I3(level3_in[705]),
   .I4(level3_in[706]),
   .I5(level3_in[707])
);

LUT6 #(
   .INIT(64'h1e82cedf1e82cedf)  
) LUT6_inst9190 (
   .O(to_level2[118]),
   .I0(level3_in[708]),
   .I1(level3_in[709]),
   .I2(level3_in[710]),
   .I3(level3_in[711]),
   .I4(level3_in[712]),
   .I5(level3_in[713])
);

LUT6 #(
   .INIT(64'h99d7f9af99d7f9af)  
) LUT6_inst9191 (
   .O(to_level2[119]),
   .I0(level3_in[714]),
   .I1(level3_in[715]),
   .I2(level3_in[716]),
   .I3(level3_in[717]),
   .I4(level3_in[718]),
   .I5(level3_in[719])
);

LUT6 #(
   .INIT(64'h280299b3280299b3)  
) LUT6_inst9192 (
   .O(to_level2[120]),
   .I0(level3_in[720]),
   .I1(level3_in[721]),
   .I2(level3_in[722]),
   .I3(level3_in[723]),
   .I4(level3_in[724]),
   .I5(level3_in[725])
);

LUT6 #(
   .INIT(64'h7f259bbe7f259bbe)  
) LUT6_inst9193 (
   .O(to_level2[121]),
   .I0(level3_in[726]),
   .I1(level3_in[727]),
   .I2(level3_in[728]),
   .I3(level3_in[729]),
   .I4(level3_in[730]),
   .I5(level3_in[731])
);

LUT6 #(
   .INIT(64'h05625d4605625d46)  
) LUT6_inst9194 (
   .O(to_level2[122]),
   .I0(level3_in[732]),
   .I1(level3_in[733]),
   .I2(level3_in[734]),
   .I3(level3_in[735]),
   .I4(level3_in[736]),
   .I5(level3_in[737])
);

LUT6 #(
   .INIT(64'he9f4607fe9f4607f)  
) LUT6_inst9195 (
   .O(to_level2[123]),
   .I0(level3_in[738]),
   .I1(level3_in[739]),
   .I2(level3_in[740]),
   .I3(level3_in[741]),
   .I4(level3_in[742]),
   .I5(level3_in[743])
);

LUT6 #(
   .INIT(64'ha271f01ba271f01b)  
) LUT6_inst9196 (
   .O(to_level2[124]),
   .I0(level3_in[744]),
   .I1(level3_in[745]),
   .I2(level3_in[746]),
   .I3(level3_in[747]),
   .I4(level3_in[748]),
   .I5(level3_in[749])
);

LUT6 #(
   .INIT(64'h56f2e27b56f2e27b)  
) LUT6_inst9197 (
   .O(to_level2[125]),
   .I0(level3_in[750]),
   .I1(level3_in[751]),
   .I2(level3_in[752]),
   .I3(level3_in[753]),
   .I4(level3_in[754]),
   .I5(level3_in[755])
);

LUT6 #(
   .INIT(64'h815d55b0815d55b0)  
) LUT6_inst9198 (
   .O(to_level2[126]),
   .I0(level3_in[756]),
   .I1(level3_in[757]),
   .I2(level3_in[758]),
   .I3(level3_in[759]),
   .I4(level3_in[760]),
   .I5(level3_in[761])
);

LUT6 #(
   .INIT(64'h8fe536118fe53611)  
) LUT6_inst9199 (
   .O(to_level2[127]),
   .I0(level3_in[762]),
   .I1(level3_in[763]),
   .I2(level3_in[764]),
   .I3(level3_in[765]),
   .I4(level3_in[766]),
   .I5(level3_in[767])
);

LUT6 #(
   .INIT(64'hb40fb385b40fb385)  
) LUT6_inst9200 (
   .O(to_level2[128]),
   .I0(level3_in[768]),
   .I1(level3_in[769]),
   .I2(level3_in[770]),
   .I3(level3_in[771]),
   .I4(level3_in[772]),
   .I5(level3_in[773])
);

LUT6 #(
   .INIT(64'h30bd40d430bd40d4)  
) LUT6_inst9201 (
   .O(to_level2[129]),
   .I0(level3_in[774]),
   .I1(level3_in[775]),
   .I2(level3_in[776]),
   .I3(level3_in[777]),
   .I4(level3_in[778]),
   .I5(level3_in[779])
);

LUT6 #(
   .INIT(64'h36e282fa36e282fa)  
) LUT6_inst9202 (
   .O(to_level2[130]),
   .I0(level3_in[780]),
   .I1(level3_in[781]),
   .I2(level3_in[782]),
   .I3(level3_in[783]),
   .I4(level3_in[784]),
   .I5(level3_in[785])
);

LUT6 #(
   .INIT(64'hd5c7172ed5c7172e)  
) LUT6_inst9203 (
   .O(to_level2[131]),
   .I0(level3_in[786]),
   .I1(level3_in[787]),
   .I2(level3_in[788]),
   .I3(level3_in[789]),
   .I4(level3_in[790]),
   .I5(level3_in[791])
);

LUT6 #(
   .INIT(64'hf5afd4a6f5afd4a6)  
) LUT6_inst9204 (
   .O(to_level2[132]),
   .I0(level3_in[792]),
   .I1(level3_in[793]),
   .I2(level3_in[794]),
   .I3(level3_in[795]),
   .I4(level3_in[796]),
   .I5(level3_in[797])
);

LUT6 #(
   .INIT(64'h11be62d211be62d2)  
) LUT6_inst9205 (
   .O(to_level2[133]),
   .I0(level3_in[798]),
   .I1(level3_in[799]),
   .I2(level3_in[800]),
   .I3(level3_in[801]),
   .I4(level3_in[802]),
   .I5(level3_in[803])
);

LUT6 #(
   .INIT(64'hcca63f64cca63f64)  
) LUT6_inst9206 (
   .O(to_level2[134]),
   .I0(level3_in[804]),
   .I1(level3_in[805]),
   .I2(level3_in[806]),
   .I3(level3_in[807]),
   .I4(level3_in[808]),
   .I5(level3_in[809])
);

LUT6 #(
   .INIT(64'h6bef40e06bef40e0)  
) LUT6_inst9207 (
   .O(to_level2[135]),
   .I0(level3_in[810]),
   .I1(level3_in[811]),
   .I2(level3_in[812]),
   .I3(level3_in[813]),
   .I4(level3_in[814]),
   .I5(level3_in[815])
);

LUT6 #(
   .INIT(64'hdfaad5a7dfaad5a7)  
) LUT6_inst9208 (
   .O(to_level2[136]),
   .I0(level3_in[816]),
   .I1(level3_in[817]),
   .I2(level3_in[818]),
   .I3(level3_in[819]),
   .I4(level3_in[820]),
   .I5(level3_in[821])
);

LUT6 #(
   .INIT(64'hd44802e0d44802e0)  
) LUT6_inst9209 (
   .O(to_level2[137]),
   .I0(level3_in[822]),
   .I1(level3_in[823]),
   .I2(level3_in[824]),
   .I3(level3_in[825]),
   .I4(level3_in[826]),
   .I5(level3_in[827])
);

LUT6 #(
   .INIT(64'h9167e22d9167e22d)  
) LUT6_inst9210 (
   .O(to_level2[138]),
   .I0(level3_in[828]),
   .I1(level3_in[829]),
   .I2(level3_in[830]),
   .I3(level3_in[831]),
   .I4(level3_in[832]),
   .I5(level3_in[833])
);

LUT6 #(
   .INIT(64'h76bd662f76bd662f)  
) LUT6_inst9211 (
   .O(to_level2[139]),
   .I0(level3_in[834]),
   .I1(level3_in[835]),
   .I2(level3_in[836]),
   .I3(level3_in[837]),
   .I4(level3_in[838]),
   .I5(level3_in[839])
);

LUT6 #(
   .INIT(64'hd2627180d2627180)  
) LUT6_inst9212 (
   .O(to_level2[140]),
   .I0(level3_in[840]),
   .I1(level3_in[841]),
   .I2(level3_in[842]),
   .I3(level3_in[843]),
   .I4(level3_in[844]),
   .I5(level3_in[845])
);

LUT6 #(
   .INIT(64'h38f5836638f58366)  
) LUT6_inst9213 (
   .O(to_level2[141]),
   .I0(level3_in[846]),
   .I1(level3_in[847]),
   .I2(level3_in[848]),
   .I3(level3_in[849]),
   .I4(level3_in[850]),
   .I5(level3_in[851])
);

LUT6 #(
   .INIT(64'h162cbdf5162cbdf5)  
) LUT6_inst9214 (
   .O(to_level2[142]),
   .I0(level3_in[852]),
   .I1(level3_in[853]),
   .I2(level3_in[854]),
   .I3(level3_in[855]),
   .I4(level3_in[856]),
   .I5(level3_in[857])
);

LUT6 #(
   .INIT(64'h4ee56f664ee56f66)  
) LUT6_inst9215 (
   .O(to_level2[143]),
   .I0(level3_in[858]),
   .I1(level3_in[859]),
   .I2(level3_in[860]),
   .I3(level3_in[861]),
   .I4(level3_in[862]),
   .I5(level3_in[863])
);

LUT6 #(
   .INIT(64'h5151f2c85151f2c8)  
) LUT6_inst9216 (
   .O(to_level2[144]),
   .I0(level3_in[864]),
   .I1(level3_in[865]),
   .I2(level3_in[866]),
   .I3(level3_in[867]),
   .I4(level3_in[868]),
   .I5(level3_in[869])
);

LUT6 #(
   .INIT(64'hff789a0fff789a0f)  
) LUT6_inst9217 (
   .O(to_level2[145]),
   .I0(level3_in[870]),
   .I1(level3_in[871]),
   .I2(level3_in[872]),
   .I3(level3_in[873]),
   .I4(level3_in[874]),
   .I5(level3_in[875])
);

LUT6 #(
   .INIT(64'h81f30f3e81f30f3e)  
) LUT6_inst9218 (
   .O(to_level2[146]),
   .I0(level3_in[876]),
   .I1(level3_in[877]),
   .I2(level3_in[878]),
   .I3(level3_in[879]),
   .I4(level3_in[880]),
   .I5(level3_in[881])
);

LUT6 #(
   .INIT(64'hf018bafff018baff)  
) LUT6_inst9219 (
   .O(to_level2[147]),
   .I0(level3_in[882]),
   .I1(level3_in[883]),
   .I2(level3_in[884]),
   .I3(level3_in[885]),
   .I4(level3_in[886]),
   .I5(level3_in[887])
);

LUT6 #(
   .INIT(64'h753c0db8753c0db8)  
) LUT6_inst9220 (
   .O(to_level2[148]),
   .I0(level3_in[888]),
   .I1(level3_in[889]),
   .I2(level3_in[890]),
   .I3(level3_in[891]),
   .I4(level3_in[892]),
   .I5(level3_in[893])
);

LUT6 #(
   .INIT(64'h909c5467909c5467)  
) LUT6_inst9221 (
   .O(to_level2[149]),
   .I0(level3_in[894]),
   .I1(level3_in[895]),
   .I2(level3_in[896]),
   .I3(level3_in[897]),
   .I4(level3_in[898]),
   .I5(level3_in[899])
);

LUT6 #(
   .INIT(64'h1d03b5081d03b508)  
) LUT6_inst9222 (
   .O(to_level2[150]),
   .I0(level3_in[900]),
   .I1(level3_in[901]),
   .I2(level3_in[902]),
   .I3(level3_in[903]),
   .I4(level3_in[904]),
   .I5(level3_in[905])
);

LUT6 #(
   .INIT(64'h9f5e34a79f5e34a7)  
) LUT6_inst9223 (
   .O(to_level2[151]),
   .I0(level3_in[906]),
   .I1(level3_in[907]),
   .I2(level3_in[908]),
   .I3(level3_in[909]),
   .I4(level3_in[910]),
   .I5(level3_in[911])
);

LUT6 #(
   .INIT(64'h7bde933a7bde933a)  
) LUT6_inst9224 (
   .O(to_level2[152]),
   .I0(level3_in[912]),
   .I1(level3_in[913]),
   .I2(level3_in[914]),
   .I3(level3_in[915]),
   .I4(level3_in[916]),
   .I5(level3_in[917])
);

LUT6 #(
   .INIT(64'ha8564ba9a8564ba9)  
) LUT6_inst9225 (
   .O(to_level2[153]),
   .I0(level3_in[918]),
   .I1(level3_in[919]),
   .I2(level3_in[920]),
   .I3(level3_in[921]),
   .I4(level3_in[922]),
   .I5(level3_in[923])
);

LUT6 #(
   .INIT(64'hf8ee0704f8ee0704)  
) LUT6_inst9226 (
   .O(to_level2[154]),
   .I0(level3_in[924]),
   .I1(level3_in[925]),
   .I2(level3_in[926]),
   .I3(level3_in[927]),
   .I4(level3_in[928]),
   .I5(level3_in[929])
);

LUT6 #(
   .INIT(64'h2fa507e82fa507e8)  
) LUT6_inst9227 (
   .O(to_level2[155]),
   .I0(level3_in[930]),
   .I1(level3_in[931]),
   .I2(level3_in[932]),
   .I3(level3_in[933]),
   .I4(level3_in[934]),
   .I5(level3_in[935])
);

LUT6 #(
   .INIT(64'h654b33c8654b33c8)  
) LUT6_inst9228 (
   .O(to_level2[156]),
   .I0(level3_in[936]),
   .I1(level3_in[937]),
   .I2(level3_in[938]),
   .I3(level3_in[939]),
   .I4(level3_in[940]),
   .I5(level3_in[941])
);

LUT6 #(
   .INIT(64'h87f159a087f159a0)  
) LUT6_inst9229 (
   .O(to_level2[157]),
   .I0(level3_in[942]),
   .I1(level3_in[943]),
   .I2(level3_in[944]),
   .I3(level3_in[945]),
   .I4(level3_in[946]),
   .I5(level3_in[947])
);

LUT6 #(
   .INIT(64'h170c98a5170c98a5)  
) LUT6_inst9230 (
   .O(to_level2[158]),
   .I0(level3_in[948]),
   .I1(level3_in[949]),
   .I2(level3_in[950]),
   .I3(level3_in[951]),
   .I4(level3_in[952]),
   .I5(level3_in[953])
);

LUT6 #(
   .INIT(64'h6d48d7e06d48d7e0)  
) LUT6_inst9231 (
   .O(to_level2[159]),
   .I0(level3_in[954]),
   .I1(level3_in[955]),
   .I2(level3_in[956]),
   .I3(level3_in[957]),
   .I4(level3_in[958]),
   .I5(level3_in[959])
);

LUT6 #(
   .INIT(64'h2780a9ac2780a9ac)  
) LUT6_inst9232 (
   .O(to_level2[160]),
   .I0(level3_in[960]),
   .I1(level3_in[961]),
   .I2(level3_in[962]),
   .I3(level3_in[963]),
   .I4(level3_in[964]),
   .I5(level3_in[965])
);

LUT6 #(
   .INIT(64'h93a2d0d993a2d0d9)  
) LUT6_inst9233 (
   .O(to_level2[161]),
   .I0(level3_in[966]),
   .I1(level3_in[967]),
   .I2(level3_in[968]),
   .I3(level3_in[969]),
   .I4(level3_in[970]),
   .I5(level3_in[971])
);

LUT6 #(
   .INIT(64'h624d7bee624d7bee)  
) LUT6_inst9234 (
   .O(to_level2[162]),
   .I0(level3_in[972]),
   .I1(level3_in[973]),
   .I2(level3_in[974]),
   .I3(level3_in[975]),
   .I4(level3_in[976]),
   .I5(level3_in[977])
);

LUT6 #(
   .INIT(64'h3897a9893897a989)  
) LUT6_inst9235 (
   .O(to_level2[163]),
   .I0(level3_in[978]),
   .I1(level3_in[979]),
   .I2(level3_in[980]),
   .I3(level3_in[981]),
   .I4(level3_in[982]),
   .I5(level3_in[983])
);

LUT6 #(
   .INIT(64'h9c124ba19c124ba1)  
) LUT6_inst9236 (
   .O(to_level2[164]),
   .I0(level3_in[984]),
   .I1(level3_in[985]),
   .I2(level3_in[986]),
   .I3(level3_in[987]),
   .I4(level3_in[988]),
   .I5(level3_in[989])
);

LUT6 #(
   .INIT(64'hf4f88262f4f88262)  
) LUT6_inst9237 (
   .O(to_level2[165]),
   .I0(level3_in[990]),
   .I1(level3_in[991]),
   .I2(level3_in[992]),
   .I3(level3_in[993]),
   .I4(level3_in[994]),
   .I5(level3_in[995])
);

LUT6 #(
   .INIT(64'ha56b1c71a56b1c71)  
) LUT6_inst9238 (
   .O(to_level2[166]),
   .I0(level3_in[996]),
   .I1(level3_in[997]),
   .I2(level3_in[998]),
   .I3(level3_in[999]),
   .I4(level3_in[1000]),
   .I5(level3_in[1001])
);

LUT6 #(
   .INIT(64'h323cf933323cf933)  
) LUT6_inst9239 (
   .O(to_level2[167]),
   .I0(level3_in[1002]),
   .I1(level3_in[1003]),
   .I2(level3_in[1004]),
   .I3(level3_in[1005]),
   .I4(level3_in[1006]),
   .I5(level3_in[1007])
);

LUT6 #(
   .INIT(64'h9430ae529430ae52)  
) LUT6_inst9240 (
   .O(to_level2[168]),
   .I0(level3_in[1008]),
   .I1(level3_in[1009]),
   .I2(level3_in[1010]),
   .I3(level3_in[1011]),
   .I4(level3_in[1012]),
   .I5(level3_in[1013])
);

LUT6 #(
   .INIT(64'he9879b37e9879b37)  
) LUT6_inst9241 (
   .O(to_level2[169]),
   .I0(level3_in[1014]),
   .I1(level3_in[1015]),
   .I2(level3_in[1016]),
   .I3(level3_in[1017]),
   .I4(level3_in[1018]),
   .I5(level3_in[1019])
);

LUT6 #(
   .INIT(64'ha27867b2a27867b2)  
) LUT6_inst9242 (
   .O(to_level2[170]),
   .I0(level3_in[1020]),
   .I1(level3_in[1021]),
   .I2(level3_in[1022]),
   .I3(level3_in[1023]),
   .I4(level3_in[1024]),
   .I5(level3_in[1025])
);

LUT6 #(
   .INIT(64'hf5c8942af5c8942a)  
) LUT6_inst9243 (
   .O(to_level2[171]),
   .I0(level3_in[1026]),
   .I1(level3_in[1027]),
   .I2(level3_in[1028]),
   .I3(level3_in[1029]),
   .I4(level3_in[1030]),
   .I5(level3_in[1031])
);

LUT6 #(
   .INIT(64'hb2bee1dbb2bee1db)  
) LUT6_inst9244 (
   .O(to_level2[172]),
   .I0(level3_in[1032]),
   .I1(level3_in[1033]),
   .I2(level3_in[1034]),
   .I3(level3_in[1035]),
   .I4(level3_in[1036]),
   .I5(level3_in[1037])
);

LUT6 #(
   .INIT(64'h440f8696440f8696)  
) LUT6_inst9245 (
   .O(to_level2[173]),
   .I0(level3_in[1038]),
   .I1(level3_in[1039]),
   .I2(level3_in[1040]),
   .I3(level3_in[1041]),
   .I4(level3_in[1042]),
   .I5(level3_in[1043])
);

LUT6 #(
   .INIT(64'h0dbea2950dbea295)  
) LUT6_inst9246 (
   .O(to_level2[174]),
   .I0(level3_in[1044]),
   .I1(level3_in[1045]),
   .I2(level3_in[1046]),
   .I3(level3_in[1047]),
   .I4(level3_in[1048]),
   .I5(level3_in[1049])
);

LUT6 #(
   .INIT(64'hfd37c20dfd37c20d)  
) LUT6_inst9247 (
   .O(to_level2[175]),
   .I0(level3_in[1050]),
   .I1(level3_in[1051]),
   .I2(level3_in[1052]),
   .I3(level3_in[1053]),
   .I4(level3_in[1054]),
   .I5(level3_in[1055])
);

LUT6 #(
   .INIT(64'hac4d83f8ac4d83f8)  
) LUT6_inst9248 (
   .O(to_level2[176]),
   .I0(level3_in[1056]),
   .I1(level3_in[1057]),
   .I2(level3_in[1058]),
   .I3(level3_in[1059]),
   .I4(level3_in[1060]),
   .I5(level3_in[1061])
);

LUT6 #(
   .INIT(64'h2c8557bf2c8557bf)  
) LUT6_inst9249 (
   .O(to_level2[177]),
   .I0(level3_in[1062]),
   .I1(level3_in[1063]),
   .I2(level3_in[1064]),
   .I3(level3_in[1065]),
   .I4(level3_in[1066]),
   .I5(level3_in[1067])
);

LUT6 #(
   .INIT(64'h52728fde52728fde)  
) LUT6_inst9250 (
   .O(to_level2[178]),
   .I0(level3_in[1068]),
   .I1(level3_in[1069]),
   .I2(level3_in[1070]),
   .I3(level3_in[1071]),
   .I4(level3_in[1072]),
   .I5(level3_in[1073])
);

LUT6 #(
   .INIT(64'h9b7c264a9b7c264a)  
) LUT6_inst9251 (
   .O(to_level2[179]),
   .I0(level3_in[1074]),
   .I1(level3_in[1075]),
   .I2(level3_in[1076]),
   .I3(level3_in[1077]),
   .I4(level3_in[1078]),
   .I5(level3_in[1079])
);

LUT6 #(
   .INIT(64'hd1d35c47d1d35c47)  
) LUT6_inst9252 (
   .O(to_level2[180]),
   .I0(level3_in[1080]),
   .I1(level3_in[1081]),
   .I2(level3_in[1082]),
   .I3(level3_in[1083]),
   .I4(level3_in[1084]),
   .I5(level3_in[1085])
);

LUT6 #(
   .INIT(64'h5d0a526f5d0a526f)  
) LUT6_inst9253 (
   .O(to_level2[181]),
   .I0(level3_in[1086]),
   .I1(level3_in[1087]),
   .I2(level3_in[1088]),
   .I3(level3_in[1089]),
   .I4(level3_in[1090]),
   .I5(level3_in[1091])
);

LUT6 #(
   .INIT(64'hfe4d10a4fe4d10a4)  
) LUT6_inst9254 (
   .O(to_level2[182]),
   .I0(level3_in[1092]),
   .I1(level3_in[1093]),
   .I2(level3_in[1094]),
   .I3(level3_in[1095]),
   .I4(level3_in[1096]),
   .I5(level3_in[1097])
);

LUT6 #(
   .INIT(64'h35b2e21035b2e210)  
) LUT6_inst9255 (
   .O(to_level2[183]),
   .I0(level3_in[1098]),
   .I1(level3_in[1099]),
   .I2(level3_in[1100]),
   .I3(level3_in[1101]),
   .I4(level3_in[1102]),
   .I5(level3_in[1103])
);

LUT6 #(
   .INIT(64'ha170b1d4a170b1d4)  
) LUT6_inst9256 (
   .O(to_level2[184]),
   .I0(level3_in[1104]),
   .I1(level3_in[1105]),
   .I2(level3_in[1106]),
   .I3(level3_in[1107]),
   .I4(level3_in[1108]),
   .I5(level3_in[1109])
);

LUT6 #(
   .INIT(64'h96d6450796d64507)  
) LUT6_inst9257 (
   .O(to_level2[185]),
   .I0(level3_in[1110]),
   .I1(level3_in[1111]),
   .I2(level3_in[1112]),
   .I3(level3_in[1113]),
   .I4(level3_in[1114]),
   .I5(level3_in[1115])
);

LUT6 #(
   .INIT(64'h45c5ef2b45c5ef2b)  
) LUT6_inst9258 (
   .O(to_level2[186]),
   .I0(level3_in[1116]),
   .I1(level3_in[1117]),
   .I2(level3_in[1118]),
   .I3(level3_in[1119]),
   .I4(level3_in[1120]),
   .I5(level3_in[1121])
);

LUT6 #(
   .INIT(64'he65e5330e65e5330)  
) LUT6_inst9259 (
   .O(to_level2[187]),
   .I0(level3_in[1122]),
   .I1(level3_in[1123]),
   .I2(level3_in[1124]),
   .I3(level3_in[1125]),
   .I4(level3_in[1126]),
   .I5(level3_in[1127])
);

LUT6 #(
   .INIT(64'h706c578d706c578d)  
) LUT6_inst9260 (
   .O(to_level2[188]),
   .I0(level3_in[1128]),
   .I1(level3_in[1129]),
   .I2(level3_in[1130]),
   .I3(level3_in[1131]),
   .I4(level3_in[1132]),
   .I5(level3_in[1133])
);

LUT6 #(
   .INIT(64'h8d586da68d586da6)  
) LUT6_inst9261 (
   .O(to_level2[189]),
   .I0(level3_in[1134]),
   .I1(level3_in[1135]),
   .I2(level3_in[1136]),
   .I3(level3_in[1137]),
   .I4(level3_in[1138]),
   .I5(level3_in[1139])
);

LUT6 #(
   .INIT(64'h8ec5c5c98ec5c5c9)  
) LUT6_inst9262 (
   .O(to_level2[190]),
   .I0(level3_in[1140]),
   .I1(level3_in[1141]),
   .I2(level3_in[1142]),
   .I3(level3_in[1143]),
   .I4(level3_in[1144]),
   .I5(level3_in[1145])
);

LUT6 #(
   .INIT(64'hecdc730aecdc730a)  
) LUT6_inst9263 (
   .O(to_level2[191]),
   .I0(level3_in[1146]),
   .I1(level3_in[1147]),
   .I2(level3_in[1148]),
   .I3(level3_in[1149]),
   .I4(level3_in[1150]),
   .I5(level3_in[1151])
);

LUT6 #(
   .INIT(64'h6a294bb16a294bb1)  
) LUT6_inst9264 (
   .O(to_level2[192]),
   .I0(level3_in[1152]),
   .I1(level3_in[1153]),
   .I2(level3_in[1154]),
   .I3(level3_in[1155]),
   .I4(level3_in[1156]),
   .I5(level3_in[1157])
);

LUT6 #(
   .INIT(64'hb91a401db91a401d)  
) LUT6_inst9265 (
   .O(to_level2[193]),
   .I0(level3_in[1158]),
   .I1(level3_in[1159]),
   .I2(level3_in[1160]),
   .I3(level3_in[1161]),
   .I4(level3_in[1162]),
   .I5(level3_in[1163])
);

LUT6 #(
   .INIT(64'he63319f5e63319f5)  
) LUT6_inst9266 (
   .O(to_level2[194]),
   .I0(level3_in[1164]),
   .I1(level3_in[1165]),
   .I2(level3_in[1166]),
   .I3(level3_in[1167]),
   .I4(level3_in[1168]),
   .I5(level3_in[1169])
);

LUT6 #(
   .INIT(64'h29c1879e29c1879e)  
) LUT6_inst9267 (
   .O(to_level2[195]),
   .I0(level3_in[1170]),
   .I1(level3_in[1171]),
   .I2(level3_in[1172]),
   .I3(level3_in[1173]),
   .I4(level3_in[1174]),
   .I5(level3_in[1175])
);

LUT6 #(
   .INIT(64'hab2f098eab2f098e)  
) LUT6_inst9268 (
   .O(to_level2[196]),
   .I0(level3_in[1176]),
   .I1(level3_in[1177]),
   .I2(level3_in[1178]),
   .I3(level3_in[1179]),
   .I4(level3_in[1180]),
   .I5(level3_in[1181])
);

LUT6 #(
   .INIT(64'hb9ece5adb9ece5ad)  
) LUT6_inst9269 (
   .O(to_level2[197]),
   .I0(level3_in[1182]),
   .I1(level3_in[1183]),
   .I2(level3_in[1184]),
   .I3(level3_in[1185]),
   .I4(level3_in[1186]),
   .I5(level3_in[1187])
);

LUT6 #(
   .INIT(64'h7d5d8a867d5d8a86)  
) LUT6_inst9270 (
   .O(to_level2[198]),
   .I0(level3_in[1188]),
   .I1(level3_in[1189]),
   .I2(level3_in[1190]),
   .I3(level3_in[1191]),
   .I4(level3_in[1192]),
   .I5(level3_in[1193])
);

LUT6 #(
   .INIT(64'h970b33ad970b33ad)  
) LUT6_inst9271 (
   .O(to_level2[199]),
   .I0(level3_in[1194]),
   .I1(level3_in[1195]),
   .I2(level3_in[1196]),
   .I3(level3_in[1197]),
   .I4(level3_in[1198]),
   .I5(level3_in[1199])
);

LUT6 #(
   .INIT(64'h382099b4382099b4)  
) LUT6_inst9272 (
   .O(to_level2[200]),
   .I0(level3_in[1200]),
   .I1(level3_in[1201]),
   .I2(level3_in[1202]),
   .I3(level3_in[1203]),
   .I4(level3_in[1204]),
   .I5(level3_in[1205])
);

LUT6 #(
   .INIT(64'hcf8a9b77cf8a9b77)  
) LUT6_inst9273 (
   .O(to_level2[201]),
   .I0(level3_in[1206]),
   .I1(level3_in[1207]),
   .I2(level3_in[1208]),
   .I3(level3_in[1209]),
   .I4(level3_in[1210]),
   .I5(level3_in[1211])
);

LUT6 #(
   .INIT(64'h2967382429673824)  
) LUT6_inst9274 (
   .O(to_level2[202]),
   .I0(level3_in[1212]),
   .I1(level3_in[1213]),
   .I2(level3_in[1214]),
   .I3(level3_in[1215]),
   .I4(level3_in[1216]),
   .I5(level3_in[1217])
);

LUT6 #(
   .INIT(64'h0270969902709699)  
) LUT6_inst9275 (
   .O(to_level2[203]),
   .I0(level3_in[1218]),
   .I1(level3_in[1219]),
   .I2(level3_in[1220]),
   .I3(level3_in[1221]),
   .I4(level3_in[1222]),
   .I5(level3_in[1223])
);

LUT6 #(
   .INIT(64'h08074fb308074fb3)  
) LUT6_inst9276 (
   .O(to_level2[204]),
   .I0(level3_in[1224]),
   .I1(level3_in[1225]),
   .I2(level3_in[1226]),
   .I3(level3_in[1227]),
   .I4(level3_in[1228]),
   .I5(level3_in[1229])
);

LUT6 #(
   .INIT(64'h3105313d3105313d)  
) LUT6_inst9277 (
   .O(to_level2[205]),
   .I0(level3_in[1230]),
   .I1(level3_in[1231]),
   .I2(level3_in[1232]),
   .I3(level3_in[1233]),
   .I4(level3_in[1234]),
   .I5(level3_in[1235])
);

LUT6 #(
   .INIT(64'hf2d2be17f2d2be17)  
) LUT6_inst9278 (
   .O(to_level2[206]),
   .I0(level3_in[1236]),
   .I1(level3_in[1237]),
   .I2(level3_in[1238]),
   .I3(level3_in[1239]),
   .I4(level3_in[1240]),
   .I5(level3_in[1241])
);

LUT6 #(
   .INIT(64'h494f3c65494f3c65)  
) LUT6_inst9279 (
   .O(to_level2[207]),
   .I0(level3_in[1242]),
   .I1(level3_in[1243]),
   .I2(level3_in[1244]),
   .I3(level3_in[1245]),
   .I4(level3_in[1246]),
   .I5(level3_in[1247])
);

LUT6 #(
   .INIT(64'he5c5bcaae5c5bcaa)  
) LUT6_inst9280 (
   .O(to_level2[208]),
   .I0(level3_in[1248]),
   .I1(level3_in[1249]),
   .I2(level3_in[1250]),
   .I3(level3_in[1251]),
   .I4(level3_in[1252]),
   .I5(level3_in[1253])
);

LUT6 #(
   .INIT(64'h4aa9f0424aa9f042)  
) LUT6_inst9281 (
   .O(to_level2[209]),
   .I0(level3_in[1254]),
   .I1(level3_in[1255]),
   .I2(level3_in[1256]),
   .I3(level3_in[1257]),
   .I4(level3_in[1258]),
   .I5(level3_in[1259])
);

LUT6 #(
   .INIT(64'h9733d2279733d227)  
) LUT6_inst9282 (
   .O(to_level2[210]),
   .I0(level3_in[1260]),
   .I1(level3_in[1261]),
   .I2(level3_in[1262]),
   .I3(level3_in[1263]),
   .I4(level3_in[1264]),
   .I5(level3_in[1265])
);

LUT6 #(
   .INIT(64'hd2bffdd2d2bffdd2)  
) LUT6_inst9283 (
   .O(to_level2[211]),
   .I0(level3_in[1266]),
   .I1(level3_in[1267]),
   .I2(level3_in[1268]),
   .I3(level3_in[1269]),
   .I4(level3_in[1270]),
   .I5(level3_in[1271])
);

LUT6 #(
   .INIT(64'h92a82e3c92a82e3c)  
) LUT6_inst9284 (
   .O(to_level2[212]),
   .I0(level3_in[1272]),
   .I1(level3_in[1273]),
   .I2(level3_in[1274]),
   .I3(level3_in[1275]),
   .I4(level3_in[1276]),
   .I5(level3_in[1277])
);

LUT6 #(
   .INIT(64'h09a88f9809a88f98)  
) LUT6_inst9285 (
   .O(to_level2[213]),
   .I0(level3_in[1278]),
   .I1(level3_in[1279]),
   .I2(level3_in[1280]),
   .I3(level3_in[1281]),
   .I4(level3_in[1282]),
   .I5(level3_in[1283])
);

LUT6 #(
   .INIT(64'hbb4a17fdbb4a17fd)  
) LUT6_inst9286 (
   .O(to_level2[214]),
   .I0(level3_in[1284]),
   .I1(level3_in[1285]),
   .I2(level3_in[1286]),
   .I3(level3_in[1287]),
   .I4(level3_in[1288]),
   .I5(level3_in[1289])
);

LUT6 #(
   .INIT(64'h673f2e45673f2e45)  
) LUT6_inst9287 (
   .O(to_level2[215]),
   .I0(level3_in[1290]),
   .I1(level3_in[1291]),
   .I2(level3_in[1292]),
   .I3(level3_in[1293]),
   .I4(level3_in[1294]),
   .I5(level3_in[1295])
);
////////////// level 2 starts below:/n
LUT6 #(
   .INIT(64'hc2e11fc9c2e11fc9)  
) LUT6_inst9288 (
   .O(to_level1[0]),
   .I0(level2_in[0]),
   .I1(level2_in[1]),
   .I2(level2_in[2]),
   .I3(level2_in[3]),
   .I4(level2_in[4]),
   .I5(level2_in[5])
);

LUT6 #(
   .INIT(64'h63aec2f463aec2f4)  
) LUT6_inst9289 (
   .O(to_level1[1]),
   .I0(level2_in[6]),
   .I1(level2_in[7]),
   .I2(level2_in[8]),
   .I3(level2_in[9]),
   .I4(level2_in[10]),
   .I5(level2_in[11])
);

LUT6 #(
   .INIT(64'h051020b3051020b3)  
) LUT6_inst9290 (
   .O(to_level1[2]),
   .I0(level2_in[12]),
   .I1(level2_in[13]),
   .I2(level2_in[14]),
   .I3(level2_in[15]),
   .I4(level2_in[16]),
   .I5(level2_in[17])
);

LUT6 #(
   .INIT(64'h5748809157488091)  
) LUT6_inst9291 (
   .O(to_level1[3]),
   .I0(level2_in[18]),
   .I1(level2_in[19]),
   .I2(level2_in[20]),
   .I3(level2_in[21]),
   .I4(level2_in[22]),
   .I5(level2_in[23])
);

LUT6 #(
   .INIT(64'hff2e7562ff2e7562)  
) LUT6_inst9292 (
   .O(to_level1[4]),
   .I0(level2_in[24]),
   .I1(level2_in[25]),
   .I2(level2_in[26]),
   .I3(level2_in[27]),
   .I4(level2_in[28]),
   .I5(level2_in[29])
);

LUT6 #(
   .INIT(64'h603136a8603136a8)  
) LUT6_inst9293 (
   .O(to_level1[5]),
   .I0(level2_in[30]),
   .I1(level2_in[31]),
   .I2(level2_in[32]),
   .I3(level2_in[33]),
   .I4(level2_in[34]),
   .I5(level2_in[35])
);

LUT6 #(
   .INIT(64'he0842754e0842754)  
) LUT6_inst9294 (
   .O(to_level1[6]),
   .I0(level2_in[36]),
   .I1(level2_in[37]),
   .I2(level2_in[38]),
   .I3(level2_in[39]),
   .I4(level2_in[40]),
   .I5(level2_in[41])
);

LUT6 #(
   .INIT(64'h03ba328a03ba328a)  
) LUT6_inst9295 (
   .O(to_level1[7]),
   .I0(level2_in[42]),
   .I1(level2_in[43]),
   .I2(level2_in[44]),
   .I3(level2_in[45]),
   .I4(level2_in[46]),
   .I5(level2_in[47])
);

LUT6 #(
   .INIT(64'ha7e492dba7e492db)  
) LUT6_inst9296 (
   .O(to_level1[8]),
   .I0(level2_in[48]),
   .I1(level2_in[49]),
   .I2(level2_in[50]),
   .I3(level2_in[51]),
   .I4(level2_in[52]),
   .I5(level2_in[53])
);

LUT6 #(
   .INIT(64'hdd3cbaaadd3cbaaa)  
) LUT6_inst9297 (
   .O(to_level1[9]),
   .I0(level2_in[54]),
   .I1(level2_in[55]),
   .I2(level2_in[56]),
   .I3(level2_in[57]),
   .I4(level2_in[58]),
   .I5(level2_in[59])
);

LUT6 #(
   .INIT(64'hecf1a649ecf1a649)  
) LUT6_inst9298 (
   .O(to_level1[10]),
   .I0(level2_in[60]),
   .I1(level2_in[61]),
   .I2(level2_in[62]),
   .I3(level2_in[63]),
   .I4(level2_in[64]),
   .I5(level2_in[65])
);

LUT6 #(
   .INIT(64'hc46fcc75c46fcc75)  
) LUT6_inst9299 (
   .O(to_level1[11]),
   .I0(level2_in[66]),
   .I1(level2_in[67]),
   .I2(level2_in[68]),
   .I3(level2_in[69]),
   .I4(level2_in[70]),
   .I5(level2_in[71])
);

LUT6 #(
   .INIT(64'h3c0f57563c0f5756)  
) LUT6_inst9300 (
   .O(to_level1[12]),
   .I0(level2_in[72]),
   .I1(level2_in[73]),
   .I2(level2_in[74]),
   .I3(level2_in[75]),
   .I4(level2_in[76]),
   .I5(level2_in[77])
);

LUT6 #(
   .INIT(64'h5b8574ae5b8574ae)  
) LUT6_inst9301 (
   .O(to_level1[13]),
   .I0(level2_in[78]),
   .I1(level2_in[79]),
   .I2(level2_in[80]),
   .I3(level2_in[81]),
   .I4(level2_in[82]),
   .I5(level2_in[83])
);

LUT6 #(
   .INIT(64'h4fb793ce4fb793ce)  
) LUT6_inst9302 (
   .O(to_level1[14]),
   .I0(level2_in[84]),
   .I1(level2_in[85]),
   .I2(level2_in[86]),
   .I3(level2_in[87]),
   .I4(level2_in[88]),
   .I5(level2_in[89])
);

LUT6 #(
   .INIT(64'ha5681747a5681747)  
) LUT6_inst9303 (
   .O(to_level1[15]),
   .I0(level2_in[90]),
   .I1(level2_in[91]),
   .I2(level2_in[92]),
   .I3(level2_in[93]),
   .I4(level2_in[94]),
   .I5(level2_in[95])
);

LUT6 #(
   .INIT(64'he575d0f7e575d0f7)  
) LUT6_inst9304 (
   .O(to_level1[16]),
   .I0(level2_in[96]),
   .I1(level2_in[97]),
   .I2(level2_in[98]),
   .I3(level2_in[99]),
   .I4(level2_in[100]),
   .I5(level2_in[101])
);

LUT6 #(
   .INIT(64'h916b2bea916b2bea)  
) LUT6_inst9305 (
   .O(to_level1[17]),
   .I0(level2_in[102]),
   .I1(level2_in[103]),
   .I2(level2_in[104]),
   .I3(level2_in[105]),
   .I4(level2_in[106]),
   .I5(level2_in[107])
);

LUT6 #(
   .INIT(64'h30507fae30507fae)  
) LUT6_inst9306 (
   .O(to_level1[18]),
   .I0(level2_in[108]),
   .I1(level2_in[109]),
   .I2(level2_in[110]),
   .I3(level2_in[111]),
   .I4(level2_in[112]),
   .I5(level2_in[113])
);

LUT6 #(
   .INIT(64'hd5ef85a6d5ef85a6)  
) LUT6_inst9307 (
   .O(to_level1[19]),
   .I0(level2_in[114]),
   .I1(level2_in[115]),
   .I2(level2_in[116]),
   .I3(level2_in[117]),
   .I4(level2_in[118]),
   .I5(level2_in[119])
);

LUT6 #(
   .INIT(64'hde65a460de65a460)  
) LUT6_inst9308 (
   .O(to_level1[20]),
   .I0(level2_in[120]),
   .I1(level2_in[121]),
   .I2(level2_in[122]),
   .I3(level2_in[123]),
   .I4(level2_in[124]),
   .I5(level2_in[125])
);

LUT6 #(
   .INIT(64'h2913b0642913b064)  
) LUT6_inst9309 (
   .O(to_level1[21]),
   .I0(level2_in[126]),
   .I1(level2_in[127]),
   .I2(level2_in[128]),
   .I3(level2_in[129]),
   .I4(level2_in[130]),
   .I5(level2_in[131])
);

LUT6 #(
   .INIT(64'hef9feb75ef9feb75)  
) LUT6_inst9310 (
   .O(to_level1[22]),
   .I0(level2_in[132]),
   .I1(level2_in[133]),
   .I2(level2_in[134]),
   .I3(level2_in[135]),
   .I4(level2_in[136]),
   .I5(level2_in[137])
);

LUT6 #(
   .INIT(64'h4b46d7d84b46d7d8)  
) LUT6_inst9311 (
   .O(to_level1[23]),
   .I0(level2_in[138]),
   .I1(level2_in[139]),
   .I2(level2_in[140]),
   .I3(level2_in[141]),
   .I4(level2_in[142]),
   .I5(level2_in[143])
);

LUT6 #(
   .INIT(64'h3505b8083505b808)  
) LUT6_inst9312 (
   .O(to_level1[24]),
   .I0(level2_in[144]),
   .I1(level2_in[145]),
   .I2(level2_in[146]),
   .I3(level2_in[147]),
   .I4(level2_in[148]),
   .I5(level2_in[149])
);

LUT6 #(
   .INIT(64'h51fdb0b351fdb0b3)  
) LUT6_inst9313 (
   .O(to_level1[25]),
   .I0(level2_in[150]),
   .I1(level2_in[151]),
   .I2(level2_in[152]),
   .I3(level2_in[153]),
   .I4(level2_in[154]),
   .I5(level2_in[155])
);

LUT6 #(
   .INIT(64'h6c3f20416c3f2041)  
) LUT6_inst9314 (
   .O(to_level1[26]),
   .I0(level2_in[156]),
   .I1(level2_in[157]),
   .I2(level2_in[158]),
   .I3(level2_in[159]),
   .I4(level2_in[160]),
   .I5(level2_in[161])
);

LUT6 #(
   .INIT(64'hdf0a38c3df0a38c3)  
) LUT6_inst9315 (
   .O(to_level1[27]),
   .I0(level2_in[162]),
   .I1(level2_in[163]),
   .I2(level2_in[164]),
   .I3(level2_in[165]),
   .I4(level2_in[166]),
   .I5(level2_in[167])
);

LUT6 #(
   .INIT(64'hf1d58fb2f1d58fb2)  
) LUT6_inst9316 (
   .O(to_level1[28]),
   .I0(level2_in[168]),
   .I1(level2_in[169]),
   .I2(level2_in[170]),
   .I3(level2_in[171]),
   .I4(level2_in[172]),
   .I5(level2_in[173])
);

LUT6 #(
   .INIT(64'hafaf072cafaf072c)  
) LUT6_inst9317 (
   .O(to_level1[29]),
   .I0(level2_in[174]),
   .I1(level2_in[175]),
   .I2(level2_in[176]),
   .I3(level2_in[177]),
   .I4(level2_in[178]),
   .I5(level2_in[179])
);

LUT6 #(
   .INIT(64'h9f44d7fe9f44d7fe)  
) LUT6_inst9318 (
   .O(to_level1[30]),
   .I0(level2_in[180]),
   .I1(level2_in[181]),
   .I2(level2_in[182]),
   .I3(level2_in[183]),
   .I4(level2_in[184]),
   .I5(level2_in[185])
);

LUT6 #(
   .INIT(64'h6ece31206ece3120)  
) LUT6_inst9319 (
   .O(to_level1[31]),
   .I0(level2_in[186]),
   .I1(level2_in[187]),
   .I2(level2_in[188]),
   .I3(level2_in[189]),
   .I4(level2_in[190]),
   .I5(level2_in[191])
);

LUT6 #(
   .INIT(64'h096cc623096cc623)  
) LUT6_inst9320 (
   .O(to_level1[32]),
   .I0(level2_in[192]),
   .I1(level2_in[193]),
   .I2(level2_in[194]),
   .I3(level2_in[195]),
   .I4(level2_in[196]),
   .I5(level2_in[197])
);

LUT6 #(
   .INIT(64'h48faeba948faeba9)  
) LUT6_inst9321 (
   .O(to_level1[33]),
   .I0(level2_in[198]),
   .I1(level2_in[199]),
   .I2(level2_in[200]),
   .I3(level2_in[201]),
   .I4(level2_in[202]),
   .I5(level2_in[203])
);

LUT6 #(
   .INIT(64'h53f9d3f953f9d3f9)  
) LUT6_inst9322 (
   .O(to_level1[34]),
   .I0(level2_in[204]),
   .I1(level2_in[205]),
   .I2(level2_in[206]),
   .I3(level2_in[207]),
   .I4(level2_in[208]),
   .I5(level2_in[209])
);

LUT6 #(
   .INIT(64'h8c7dc8158c7dc815)  
) LUT6_inst9323 (
   .O(to_level1[35]),
   .I0(level2_in[210]),
   .I1(level2_in[211]),
   .I2(level2_in[212]),
   .I3(level2_in[213]),
   .I4(level2_in[214]),
   .I5(level2_in[215])
);
////////////// level 1 starts below:/n
LUT6 #(
   .INIT(64'h2b7ba7a32b7ba7a3)  
) LUT6_inst9324 (
   .O(to_level0[0]),
   .I0(level1_in[0]),
   .I1(level1_in[1]),
   .I2(level1_in[2]),
   .I3(level1_in[3]),
   .I4(level1_in[4]),
   .I5(level1_in[5])
);

LUT6 #(
   .INIT(64'h5bb6f0cf5bb6f0cf)  
) LUT6_inst9325 (
   .O(to_level0[1]),
   .I0(level1_in[6]),
   .I1(level1_in[7]),
   .I2(level1_in[8]),
   .I3(level1_in[9]),
   .I4(level1_in[10]),
   .I5(level1_in[11])
);

LUT6 #(
   .INIT(64'h7683b6517683b651)  
) LUT6_inst9326 (
   .O(to_level0[2]),
   .I0(level1_in[12]),
   .I1(level1_in[13]),
   .I2(level1_in[14]),
   .I3(level1_in[15]),
   .I4(level1_in[16]),
   .I5(level1_in[17])
);

LUT6 #(
   .INIT(64'hff0d4eabff0d4eab)  
) LUT6_inst9327 (
   .O(to_level0[3]),
   .I0(level1_in[18]),
   .I1(level1_in[19]),
   .I2(level1_in[20]),
   .I3(level1_in[21]),
   .I4(level1_in[22]),
   .I5(level1_in[23])
);

LUT6 #(
   .INIT(64'h09eada2609eada26)  
) LUT6_inst9328 (
   .O(to_level0[4]),
   .I0(level1_in[24]),
   .I1(level1_in[25]),
   .I2(level1_in[26]),
   .I3(level1_in[27]),
   .I4(level1_in[28]),
   .I5(level1_in[29])
);

LUT6 #(
   .INIT(64'hf70457b9f70457b9)  
) LUT6_inst9329 (
   .O(to_level0[5]),
   .I0(level1_in[30]),
   .I1(level1_in[31]),
   .I2(level1_in[32]),
   .I3(level1_in[33]),
   .I4(level1_in[34]),
   .I5(level1_in[35])
);
////////////// level 0 starts below:/n
LUT6 #(
   .INIT(64'h8e9f3c048e9f3c04)  
) LUT6_inst9330 (
   .O(data_out_temp),
   .I0(level0_in[0]),
   .I1(level0_in[1]),
   .I2(level0_in[2]),
   .I3(level0_in[3]),
   .I4(level0_in[4]),
   .I5(level0_in[5])
);

endmodule