
module lut_4level_tree4(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [7775:0] data_in,
                       input       data_valid,
                       output  reg data_out     
                       );

wire    [7775:0] to_level4;
(*S="TRUE"*)reg     [7775:0] level4_in;
wire    [1295:0] to_level3;
(*S="TRUE"*)reg     [1295:0] level3_in;
wire    [215:0] to_level2;
(*S="TRUE"*)reg     [215:0] level2_in;
wire    [35:0] to_level1;
(*S="TRUE"*)reg     [35:0] level1_in;
wire    [5:0] to_level0;
(*S="TRUE"*)reg     [5:0] level0_in;
wire          data_out_temp;


assign  to_level4 = data_in;

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level4_in <= 7776'b0;
  else
    level4_in <= to_level4;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level3_in <= 1296'b0;
  else
    level3_in <= to_level3;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level2_in <= 216'b0;
  else
    level2_in <= to_level2;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level1_in <= 36'b0;
  else
    level1_in <= to_level1;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level0_in <= 6'b0;
  else
    level0_in <= to_level0;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    data_out <= 1'b0;
  else
    if(data_valid == 1'b1)
      data_out <= data_out_temp;
    else;
end
////////////// level 4 starts below:/n
LUT6 #(
   .INIT(64'h4e5c4a734e5c4a73)  
) LUT6_inst7776 (
   .O(to_level3[0]),
   .I0(level4_in[0]),
   .I1(level4_in[1]),
   .I2(level4_in[2]),
   .I3(level4_in[3]),
   .I4(level4_in[4]),
   .I5(level4_in[5])
);

LUT6 #(
   .INIT(64'h3615d5a93615d5a9)  
) LUT6_inst7777 (
   .O(to_level3[1]),
   .I0(level4_in[6]),
   .I1(level4_in[7]),
   .I2(level4_in[8]),
   .I3(level4_in[9]),
   .I4(level4_in[10]),
   .I5(level4_in[11])
);

LUT6 #(
   .INIT(64'h2a051f4c2a051f4c)  
) LUT6_inst7778 (
   .O(to_level3[2]),
   .I0(level4_in[12]),
   .I1(level4_in[13]),
   .I2(level4_in[14]),
   .I3(level4_in[15]),
   .I4(level4_in[16]),
   .I5(level4_in[17])
);

LUT6 #(
   .INIT(64'h9c36c5f69c36c5f6)  
) LUT6_inst7779 (
   .O(to_level3[3]),
   .I0(level4_in[18]),
   .I1(level4_in[19]),
   .I2(level4_in[20]),
   .I3(level4_in[21]),
   .I4(level4_in[22]),
   .I5(level4_in[23])
);

LUT6 #(
   .INIT(64'hb338ba39b338ba39)  
) LUT6_inst7780 (
   .O(to_level3[4]),
   .I0(level4_in[24]),
   .I1(level4_in[25]),
   .I2(level4_in[26]),
   .I3(level4_in[27]),
   .I4(level4_in[28]),
   .I5(level4_in[29])
);

LUT6 #(
   .INIT(64'hd57bf3d7d57bf3d7)  
) LUT6_inst7781 (
   .O(to_level3[5]),
   .I0(level4_in[30]),
   .I1(level4_in[31]),
   .I2(level4_in[32]),
   .I3(level4_in[33]),
   .I4(level4_in[34]),
   .I5(level4_in[35])
);

LUT6 #(
   .INIT(64'he9ea4191e9ea4191)  
) LUT6_inst7782 (
   .O(to_level3[6]),
   .I0(level4_in[36]),
   .I1(level4_in[37]),
   .I2(level4_in[38]),
   .I3(level4_in[39]),
   .I4(level4_in[40]),
   .I5(level4_in[41])
);

LUT6 #(
   .INIT(64'h4fecea484fecea48)  
) LUT6_inst7783 (
   .O(to_level3[7]),
   .I0(level4_in[42]),
   .I1(level4_in[43]),
   .I2(level4_in[44]),
   .I3(level4_in[45]),
   .I4(level4_in[46]),
   .I5(level4_in[47])
);

LUT6 #(
   .INIT(64'hed30d429ed30d429)  
) LUT6_inst7784 (
   .O(to_level3[8]),
   .I0(level4_in[48]),
   .I1(level4_in[49]),
   .I2(level4_in[50]),
   .I3(level4_in[51]),
   .I4(level4_in[52]),
   .I5(level4_in[53])
);

LUT6 #(
   .INIT(64'ha7c51126a7c51126)  
) LUT6_inst7785 (
   .O(to_level3[9]),
   .I0(level4_in[54]),
   .I1(level4_in[55]),
   .I2(level4_in[56]),
   .I3(level4_in[57]),
   .I4(level4_in[58]),
   .I5(level4_in[59])
);

LUT6 #(
   .INIT(64'h4ff87e4b4ff87e4b)  
) LUT6_inst7786 (
   .O(to_level3[10]),
   .I0(level4_in[60]),
   .I1(level4_in[61]),
   .I2(level4_in[62]),
   .I3(level4_in[63]),
   .I4(level4_in[64]),
   .I5(level4_in[65])
);

LUT6 #(
   .INIT(64'hf5118450f5118450)  
) LUT6_inst7787 (
   .O(to_level3[11]),
   .I0(level4_in[66]),
   .I1(level4_in[67]),
   .I2(level4_in[68]),
   .I3(level4_in[69]),
   .I4(level4_in[70]),
   .I5(level4_in[71])
);

LUT6 #(
   .INIT(64'h3764cbb73764cbb7)  
) LUT6_inst7788 (
   .O(to_level3[12]),
   .I0(level4_in[72]),
   .I1(level4_in[73]),
   .I2(level4_in[74]),
   .I3(level4_in[75]),
   .I4(level4_in[76]),
   .I5(level4_in[77])
);

LUT6 #(
   .INIT(64'hf6135ff7f6135ff7)  
) LUT6_inst7789 (
   .O(to_level3[13]),
   .I0(level4_in[78]),
   .I1(level4_in[79]),
   .I2(level4_in[80]),
   .I3(level4_in[81]),
   .I4(level4_in[82]),
   .I5(level4_in[83])
);

LUT6 #(
   .INIT(64'h7d94b4187d94b418)  
) LUT6_inst7790 (
   .O(to_level3[14]),
   .I0(level4_in[84]),
   .I1(level4_in[85]),
   .I2(level4_in[86]),
   .I3(level4_in[87]),
   .I4(level4_in[88]),
   .I5(level4_in[89])
);

LUT6 #(
   .INIT(64'he5632472e5632472)  
) LUT6_inst7791 (
   .O(to_level3[15]),
   .I0(level4_in[90]),
   .I1(level4_in[91]),
   .I2(level4_in[92]),
   .I3(level4_in[93]),
   .I4(level4_in[94]),
   .I5(level4_in[95])
);

LUT6 #(
   .INIT(64'h654fb6ff654fb6ff)  
) LUT6_inst7792 (
   .O(to_level3[16]),
   .I0(level4_in[96]),
   .I1(level4_in[97]),
   .I2(level4_in[98]),
   .I3(level4_in[99]),
   .I4(level4_in[100]),
   .I5(level4_in[101])
);

LUT6 #(
   .INIT(64'hf7f35c90f7f35c90)  
) LUT6_inst7793 (
   .O(to_level3[17]),
   .I0(level4_in[102]),
   .I1(level4_in[103]),
   .I2(level4_in[104]),
   .I3(level4_in[105]),
   .I4(level4_in[106]),
   .I5(level4_in[107])
);

LUT6 #(
   .INIT(64'h9a60d0ce9a60d0ce)  
) LUT6_inst7794 (
   .O(to_level3[18]),
   .I0(level4_in[108]),
   .I1(level4_in[109]),
   .I2(level4_in[110]),
   .I3(level4_in[111]),
   .I4(level4_in[112]),
   .I5(level4_in[113])
);

LUT6 #(
   .INIT(64'h612edad6612edad6)  
) LUT6_inst7795 (
   .O(to_level3[19]),
   .I0(level4_in[114]),
   .I1(level4_in[115]),
   .I2(level4_in[116]),
   .I3(level4_in[117]),
   .I4(level4_in[118]),
   .I5(level4_in[119])
);

LUT6 #(
   .INIT(64'h54cc1b1f54cc1b1f)  
) LUT6_inst7796 (
   .O(to_level3[20]),
   .I0(level4_in[120]),
   .I1(level4_in[121]),
   .I2(level4_in[122]),
   .I3(level4_in[123]),
   .I4(level4_in[124]),
   .I5(level4_in[125])
);

LUT6 #(
   .INIT(64'h462f9949462f9949)  
) LUT6_inst7797 (
   .O(to_level3[21]),
   .I0(level4_in[126]),
   .I1(level4_in[127]),
   .I2(level4_in[128]),
   .I3(level4_in[129]),
   .I4(level4_in[130]),
   .I5(level4_in[131])
);

LUT6 #(
   .INIT(64'h278d42c4278d42c4)  
) LUT6_inst7798 (
   .O(to_level3[22]),
   .I0(level4_in[132]),
   .I1(level4_in[133]),
   .I2(level4_in[134]),
   .I3(level4_in[135]),
   .I4(level4_in[136]),
   .I5(level4_in[137])
);

LUT6 #(
   .INIT(64'h10db65b710db65b7)  
) LUT6_inst7799 (
   .O(to_level3[23]),
   .I0(level4_in[138]),
   .I1(level4_in[139]),
   .I2(level4_in[140]),
   .I3(level4_in[141]),
   .I4(level4_in[142]),
   .I5(level4_in[143])
);

LUT6 #(
   .INIT(64'hd91e4f0bd91e4f0b)  
) LUT6_inst7800 (
   .O(to_level3[24]),
   .I0(level4_in[144]),
   .I1(level4_in[145]),
   .I2(level4_in[146]),
   .I3(level4_in[147]),
   .I4(level4_in[148]),
   .I5(level4_in[149])
);

LUT6 #(
   .INIT(64'h780d2602780d2602)  
) LUT6_inst7801 (
   .O(to_level3[25]),
   .I0(level4_in[150]),
   .I1(level4_in[151]),
   .I2(level4_in[152]),
   .I3(level4_in[153]),
   .I4(level4_in[154]),
   .I5(level4_in[155])
);

LUT6 #(
   .INIT(64'hae7416aaae7416aa)  
) LUT6_inst7802 (
   .O(to_level3[26]),
   .I0(level4_in[156]),
   .I1(level4_in[157]),
   .I2(level4_in[158]),
   .I3(level4_in[159]),
   .I4(level4_in[160]),
   .I5(level4_in[161])
);

LUT6 #(
   .INIT(64'ha47e1727a47e1727)  
) LUT6_inst7803 (
   .O(to_level3[27]),
   .I0(level4_in[162]),
   .I1(level4_in[163]),
   .I2(level4_in[164]),
   .I3(level4_in[165]),
   .I4(level4_in[166]),
   .I5(level4_in[167])
);

LUT6 #(
   .INIT(64'h21182bda21182bda)  
) LUT6_inst7804 (
   .O(to_level3[28]),
   .I0(level4_in[168]),
   .I1(level4_in[169]),
   .I2(level4_in[170]),
   .I3(level4_in[171]),
   .I4(level4_in[172]),
   .I5(level4_in[173])
);

LUT6 #(
   .INIT(64'h5c30b50d5c30b50d)  
) LUT6_inst7805 (
   .O(to_level3[29]),
   .I0(level4_in[174]),
   .I1(level4_in[175]),
   .I2(level4_in[176]),
   .I3(level4_in[177]),
   .I4(level4_in[178]),
   .I5(level4_in[179])
);

LUT6 #(
   .INIT(64'hc02f2eb0c02f2eb0)  
) LUT6_inst7806 (
   .O(to_level3[30]),
   .I0(level4_in[180]),
   .I1(level4_in[181]),
   .I2(level4_in[182]),
   .I3(level4_in[183]),
   .I4(level4_in[184]),
   .I5(level4_in[185])
);

LUT6 #(
   .INIT(64'h0778120a0778120a)  
) LUT6_inst7807 (
   .O(to_level3[31]),
   .I0(level4_in[186]),
   .I1(level4_in[187]),
   .I2(level4_in[188]),
   .I3(level4_in[189]),
   .I4(level4_in[190]),
   .I5(level4_in[191])
);

LUT6 #(
   .INIT(64'h93c7563893c75638)  
) LUT6_inst7808 (
   .O(to_level3[32]),
   .I0(level4_in[192]),
   .I1(level4_in[193]),
   .I2(level4_in[194]),
   .I3(level4_in[195]),
   .I4(level4_in[196]),
   .I5(level4_in[197])
);

LUT6 #(
   .INIT(64'he6e7b711e6e7b711)  
) LUT6_inst7809 (
   .O(to_level3[33]),
   .I0(level4_in[198]),
   .I1(level4_in[199]),
   .I2(level4_in[200]),
   .I3(level4_in[201]),
   .I4(level4_in[202]),
   .I5(level4_in[203])
);

LUT6 #(
   .INIT(64'h88e1c94d88e1c94d)  
) LUT6_inst7810 (
   .O(to_level3[34]),
   .I0(level4_in[204]),
   .I1(level4_in[205]),
   .I2(level4_in[206]),
   .I3(level4_in[207]),
   .I4(level4_in[208]),
   .I5(level4_in[209])
);

LUT6 #(
   .INIT(64'h3ca6076a3ca6076a)  
) LUT6_inst7811 (
   .O(to_level3[35]),
   .I0(level4_in[210]),
   .I1(level4_in[211]),
   .I2(level4_in[212]),
   .I3(level4_in[213]),
   .I4(level4_in[214]),
   .I5(level4_in[215])
);

LUT6 #(
   .INIT(64'h8cb727f68cb727f6)  
) LUT6_inst7812 (
   .O(to_level3[36]),
   .I0(level4_in[216]),
   .I1(level4_in[217]),
   .I2(level4_in[218]),
   .I3(level4_in[219]),
   .I4(level4_in[220]),
   .I5(level4_in[221])
);

LUT6 #(
   .INIT(64'h378e2e0b378e2e0b)  
) LUT6_inst7813 (
   .O(to_level3[37]),
   .I0(level4_in[222]),
   .I1(level4_in[223]),
   .I2(level4_in[224]),
   .I3(level4_in[225]),
   .I4(level4_in[226]),
   .I5(level4_in[227])
);

LUT6 #(
   .INIT(64'hc87b169dc87b169d)  
) LUT6_inst7814 (
   .O(to_level3[38]),
   .I0(level4_in[228]),
   .I1(level4_in[229]),
   .I2(level4_in[230]),
   .I3(level4_in[231]),
   .I4(level4_in[232]),
   .I5(level4_in[233])
);

LUT6 #(
   .INIT(64'h6d2359e56d2359e5)  
) LUT6_inst7815 (
   .O(to_level3[39]),
   .I0(level4_in[234]),
   .I1(level4_in[235]),
   .I2(level4_in[236]),
   .I3(level4_in[237]),
   .I4(level4_in[238]),
   .I5(level4_in[239])
);

LUT6 #(
   .INIT(64'ha5de68baa5de68ba)  
) LUT6_inst7816 (
   .O(to_level3[40]),
   .I0(level4_in[240]),
   .I1(level4_in[241]),
   .I2(level4_in[242]),
   .I3(level4_in[243]),
   .I4(level4_in[244]),
   .I5(level4_in[245])
);

LUT6 #(
   .INIT(64'h840ecebb840ecebb)  
) LUT6_inst7817 (
   .O(to_level3[41]),
   .I0(level4_in[246]),
   .I1(level4_in[247]),
   .I2(level4_in[248]),
   .I3(level4_in[249]),
   .I4(level4_in[250]),
   .I5(level4_in[251])
);

LUT6 #(
   .INIT(64'hdbebd89edbebd89e)  
) LUT6_inst7818 (
   .O(to_level3[42]),
   .I0(level4_in[252]),
   .I1(level4_in[253]),
   .I2(level4_in[254]),
   .I3(level4_in[255]),
   .I4(level4_in[256]),
   .I5(level4_in[257])
);

LUT6 #(
   .INIT(64'hee95fa4eee95fa4e)  
) LUT6_inst7819 (
   .O(to_level3[43]),
   .I0(level4_in[258]),
   .I1(level4_in[259]),
   .I2(level4_in[260]),
   .I3(level4_in[261]),
   .I4(level4_in[262]),
   .I5(level4_in[263])
);

LUT6 #(
   .INIT(64'h9b70a10c9b70a10c)  
) LUT6_inst7820 (
   .O(to_level3[44]),
   .I0(level4_in[264]),
   .I1(level4_in[265]),
   .I2(level4_in[266]),
   .I3(level4_in[267]),
   .I4(level4_in[268]),
   .I5(level4_in[269])
);

LUT6 #(
   .INIT(64'h5faad9a65faad9a6)  
) LUT6_inst7821 (
   .O(to_level3[45]),
   .I0(level4_in[270]),
   .I1(level4_in[271]),
   .I2(level4_in[272]),
   .I3(level4_in[273]),
   .I4(level4_in[274]),
   .I5(level4_in[275])
);

LUT6 #(
   .INIT(64'he6eb6e75e6eb6e75)  
) LUT6_inst7822 (
   .O(to_level3[46]),
   .I0(level4_in[276]),
   .I1(level4_in[277]),
   .I2(level4_in[278]),
   .I3(level4_in[279]),
   .I4(level4_in[280]),
   .I5(level4_in[281])
);

LUT6 #(
   .INIT(64'h4a1fae2c4a1fae2c)  
) LUT6_inst7823 (
   .O(to_level3[47]),
   .I0(level4_in[282]),
   .I1(level4_in[283]),
   .I2(level4_in[284]),
   .I3(level4_in[285]),
   .I4(level4_in[286]),
   .I5(level4_in[287])
);

LUT6 #(
   .INIT(64'h696e2d4c696e2d4c)  
) LUT6_inst7824 (
   .O(to_level3[48]),
   .I0(level4_in[288]),
   .I1(level4_in[289]),
   .I2(level4_in[290]),
   .I3(level4_in[291]),
   .I4(level4_in[292]),
   .I5(level4_in[293])
);

LUT6 #(
   .INIT(64'h2e3563852e356385)  
) LUT6_inst7825 (
   .O(to_level3[49]),
   .I0(level4_in[294]),
   .I1(level4_in[295]),
   .I2(level4_in[296]),
   .I3(level4_in[297]),
   .I4(level4_in[298]),
   .I5(level4_in[299])
);

LUT6 #(
   .INIT(64'h9541ccf99541ccf9)  
) LUT6_inst7826 (
   .O(to_level3[50]),
   .I0(level4_in[300]),
   .I1(level4_in[301]),
   .I2(level4_in[302]),
   .I3(level4_in[303]),
   .I4(level4_in[304]),
   .I5(level4_in[305])
);

LUT6 #(
   .INIT(64'h27f1ba0a27f1ba0a)  
) LUT6_inst7827 (
   .O(to_level3[51]),
   .I0(level4_in[306]),
   .I1(level4_in[307]),
   .I2(level4_in[308]),
   .I3(level4_in[309]),
   .I4(level4_in[310]),
   .I5(level4_in[311])
);

LUT6 #(
   .INIT(64'h1dc4c5fc1dc4c5fc)  
) LUT6_inst7828 (
   .O(to_level3[52]),
   .I0(level4_in[312]),
   .I1(level4_in[313]),
   .I2(level4_in[314]),
   .I3(level4_in[315]),
   .I4(level4_in[316]),
   .I5(level4_in[317])
);

LUT6 #(
   .INIT(64'hb2dc20b6b2dc20b6)  
) LUT6_inst7829 (
   .O(to_level3[53]),
   .I0(level4_in[318]),
   .I1(level4_in[319]),
   .I2(level4_in[320]),
   .I3(level4_in[321]),
   .I4(level4_in[322]),
   .I5(level4_in[323])
);

LUT6 #(
   .INIT(64'h8c70b3f98c70b3f9)  
) LUT6_inst7830 (
   .O(to_level3[54]),
   .I0(level4_in[324]),
   .I1(level4_in[325]),
   .I2(level4_in[326]),
   .I3(level4_in[327]),
   .I4(level4_in[328]),
   .I5(level4_in[329])
);

LUT6 #(
   .INIT(64'h5117215951172159)  
) LUT6_inst7831 (
   .O(to_level3[55]),
   .I0(level4_in[330]),
   .I1(level4_in[331]),
   .I2(level4_in[332]),
   .I3(level4_in[333]),
   .I4(level4_in[334]),
   .I5(level4_in[335])
);

LUT6 #(
   .INIT(64'hd12b1334d12b1334)  
) LUT6_inst7832 (
   .O(to_level3[56]),
   .I0(level4_in[336]),
   .I1(level4_in[337]),
   .I2(level4_in[338]),
   .I3(level4_in[339]),
   .I4(level4_in[340]),
   .I5(level4_in[341])
);

LUT6 #(
   .INIT(64'hf5f9569bf5f9569b)  
) LUT6_inst7833 (
   .O(to_level3[57]),
   .I0(level4_in[342]),
   .I1(level4_in[343]),
   .I2(level4_in[344]),
   .I3(level4_in[345]),
   .I4(level4_in[346]),
   .I5(level4_in[347])
);

LUT6 #(
   .INIT(64'h7927973679279736)  
) LUT6_inst7834 (
   .O(to_level3[58]),
   .I0(level4_in[348]),
   .I1(level4_in[349]),
   .I2(level4_in[350]),
   .I3(level4_in[351]),
   .I4(level4_in[352]),
   .I5(level4_in[353])
);

LUT6 #(
   .INIT(64'hdcb8995ddcb8995d)  
) LUT6_inst7835 (
   .O(to_level3[59]),
   .I0(level4_in[354]),
   .I1(level4_in[355]),
   .I2(level4_in[356]),
   .I3(level4_in[357]),
   .I4(level4_in[358]),
   .I5(level4_in[359])
);

LUT6 #(
   .INIT(64'h2779344e2779344e)  
) LUT6_inst7836 (
   .O(to_level3[60]),
   .I0(level4_in[360]),
   .I1(level4_in[361]),
   .I2(level4_in[362]),
   .I3(level4_in[363]),
   .I4(level4_in[364]),
   .I5(level4_in[365])
);

LUT6 #(
   .INIT(64'he8a3087be8a3087b)  
) LUT6_inst7837 (
   .O(to_level3[61]),
   .I0(level4_in[366]),
   .I1(level4_in[367]),
   .I2(level4_in[368]),
   .I3(level4_in[369]),
   .I4(level4_in[370]),
   .I5(level4_in[371])
);

LUT6 #(
   .INIT(64'h61935a4561935a45)  
) LUT6_inst7838 (
   .O(to_level3[62]),
   .I0(level4_in[372]),
   .I1(level4_in[373]),
   .I2(level4_in[374]),
   .I3(level4_in[375]),
   .I4(level4_in[376]),
   .I5(level4_in[377])
);

LUT6 #(
   .INIT(64'hc87c474fc87c474f)  
) LUT6_inst7839 (
   .O(to_level3[63]),
   .I0(level4_in[378]),
   .I1(level4_in[379]),
   .I2(level4_in[380]),
   .I3(level4_in[381]),
   .I4(level4_in[382]),
   .I5(level4_in[383])
);

LUT6 #(
   .INIT(64'h7810013c7810013c)  
) LUT6_inst7840 (
   .O(to_level3[64]),
   .I0(level4_in[384]),
   .I1(level4_in[385]),
   .I2(level4_in[386]),
   .I3(level4_in[387]),
   .I4(level4_in[388]),
   .I5(level4_in[389])
);

LUT6 #(
   .INIT(64'hc62fbe82c62fbe82)  
) LUT6_inst7841 (
   .O(to_level3[65]),
   .I0(level4_in[390]),
   .I1(level4_in[391]),
   .I2(level4_in[392]),
   .I3(level4_in[393]),
   .I4(level4_in[394]),
   .I5(level4_in[395])
);

LUT6 #(
   .INIT(64'h735cb1c2735cb1c2)  
) LUT6_inst7842 (
   .O(to_level3[66]),
   .I0(level4_in[396]),
   .I1(level4_in[397]),
   .I2(level4_in[398]),
   .I3(level4_in[399]),
   .I4(level4_in[400]),
   .I5(level4_in[401])
);

LUT6 #(
   .INIT(64'h6b62515e6b62515e)  
) LUT6_inst7843 (
   .O(to_level3[67]),
   .I0(level4_in[402]),
   .I1(level4_in[403]),
   .I2(level4_in[404]),
   .I3(level4_in[405]),
   .I4(level4_in[406]),
   .I5(level4_in[407])
);

LUT6 #(
   .INIT(64'h87dff9f287dff9f2)  
) LUT6_inst7844 (
   .O(to_level3[68]),
   .I0(level4_in[408]),
   .I1(level4_in[409]),
   .I2(level4_in[410]),
   .I3(level4_in[411]),
   .I4(level4_in[412]),
   .I5(level4_in[413])
);

LUT6 #(
   .INIT(64'hf04adccff04adccf)  
) LUT6_inst7845 (
   .O(to_level3[69]),
   .I0(level4_in[414]),
   .I1(level4_in[415]),
   .I2(level4_in[416]),
   .I3(level4_in[417]),
   .I4(level4_in[418]),
   .I5(level4_in[419])
);

LUT6 #(
   .INIT(64'he5570f0ae5570f0a)  
) LUT6_inst7846 (
   .O(to_level3[70]),
   .I0(level4_in[420]),
   .I1(level4_in[421]),
   .I2(level4_in[422]),
   .I3(level4_in[423]),
   .I4(level4_in[424]),
   .I5(level4_in[425])
);

LUT6 #(
   .INIT(64'h23f93d8a23f93d8a)  
) LUT6_inst7847 (
   .O(to_level3[71]),
   .I0(level4_in[426]),
   .I1(level4_in[427]),
   .I2(level4_in[428]),
   .I3(level4_in[429]),
   .I4(level4_in[430]),
   .I5(level4_in[431])
);

LUT6 #(
   .INIT(64'h20d1468920d14689)  
) LUT6_inst7848 (
   .O(to_level3[72]),
   .I0(level4_in[432]),
   .I1(level4_in[433]),
   .I2(level4_in[434]),
   .I3(level4_in[435]),
   .I4(level4_in[436]),
   .I5(level4_in[437])
);

LUT6 #(
   .INIT(64'he3324b47e3324b47)  
) LUT6_inst7849 (
   .O(to_level3[73]),
   .I0(level4_in[438]),
   .I1(level4_in[439]),
   .I2(level4_in[440]),
   .I3(level4_in[441]),
   .I4(level4_in[442]),
   .I5(level4_in[443])
);

LUT6 #(
   .INIT(64'h37f43a7237f43a72)  
) LUT6_inst7850 (
   .O(to_level3[74]),
   .I0(level4_in[444]),
   .I1(level4_in[445]),
   .I2(level4_in[446]),
   .I3(level4_in[447]),
   .I4(level4_in[448]),
   .I5(level4_in[449])
);

LUT6 #(
   .INIT(64'ha80b42cba80b42cb)  
) LUT6_inst7851 (
   .O(to_level3[75]),
   .I0(level4_in[450]),
   .I1(level4_in[451]),
   .I2(level4_in[452]),
   .I3(level4_in[453]),
   .I4(level4_in[454]),
   .I5(level4_in[455])
);

LUT6 #(
   .INIT(64'h65cdb79e65cdb79e)  
) LUT6_inst7852 (
   .O(to_level3[76]),
   .I0(level4_in[456]),
   .I1(level4_in[457]),
   .I2(level4_in[458]),
   .I3(level4_in[459]),
   .I4(level4_in[460]),
   .I5(level4_in[461])
);

LUT6 #(
   .INIT(64'h5170a0f25170a0f2)  
) LUT6_inst7853 (
   .O(to_level3[77]),
   .I0(level4_in[462]),
   .I1(level4_in[463]),
   .I2(level4_in[464]),
   .I3(level4_in[465]),
   .I4(level4_in[466]),
   .I5(level4_in[467])
);

LUT6 #(
   .INIT(64'he103f752e103f752)  
) LUT6_inst7854 (
   .O(to_level3[78]),
   .I0(level4_in[468]),
   .I1(level4_in[469]),
   .I2(level4_in[470]),
   .I3(level4_in[471]),
   .I4(level4_in[472]),
   .I5(level4_in[473])
);

LUT6 #(
   .INIT(64'haad069fcaad069fc)  
) LUT6_inst7855 (
   .O(to_level3[79]),
   .I0(level4_in[474]),
   .I1(level4_in[475]),
   .I2(level4_in[476]),
   .I3(level4_in[477]),
   .I4(level4_in[478]),
   .I5(level4_in[479])
);

LUT6 #(
   .INIT(64'h7288c8e67288c8e6)  
) LUT6_inst7856 (
   .O(to_level3[80]),
   .I0(level4_in[480]),
   .I1(level4_in[481]),
   .I2(level4_in[482]),
   .I3(level4_in[483]),
   .I4(level4_in[484]),
   .I5(level4_in[485])
);

LUT6 #(
   .INIT(64'h18f9248f18f9248f)  
) LUT6_inst7857 (
   .O(to_level3[81]),
   .I0(level4_in[486]),
   .I1(level4_in[487]),
   .I2(level4_in[488]),
   .I3(level4_in[489]),
   .I4(level4_in[490]),
   .I5(level4_in[491])
);

LUT6 #(
   .INIT(64'hc3ce8bb5c3ce8bb5)  
) LUT6_inst7858 (
   .O(to_level3[82]),
   .I0(level4_in[492]),
   .I1(level4_in[493]),
   .I2(level4_in[494]),
   .I3(level4_in[495]),
   .I4(level4_in[496]),
   .I5(level4_in[497])
);

LUT6 #(
   .INIT(64'h012c38dc012c38dc)  
) LUT6_inst7859 (
   .O(to_level3[83]),
   .I0(level4_in[498]),
   .I1(level4_in[499]),
   .I2(level4_in[500]),
   .I3(level4_in[501]),
   .I4(level4_in[502]),
   .I5(level4_in[503])
);

LUT6 #(
   .INIT(64'h8d9288158d928815)  
) LUT6_inst7860 (
   .O(to_level3[84]),
   .I0(level4_in[504]),
   .I1(level4_in[505]),
   .I2(level4_in[506]),
   .I3(level4_in[507]),
   .I4(level4_in[508]),
   .I5(level4_in[509])
);

LUT6 #(
   .INIT(64'h1b3eb0cf1b3eb0cf)  
) LUT6_inst7861 (
   .O(to_level3[85]),
   .I0(level4_in[510]),
   .I1(level4_in[511]),
   .I2(level4_in[512]),
   .I3(level4_in[513]),
   .I4(level4_in[514]),
   .I5(level4_in[515])
);

LUT6 #(
   .INIT(64'ha5caeecea5caeece)  
) LUT6_inst7862 (
   .O(to_level3[86]),
   .I0(level4_in[516]),
   .I1(level4_in[517]),
   .I2(level4_in[518]),
   .I3(level4_in[519]),
   .I4(level4_in[520]),
   .I5(level4_in[521])
);

LUT6 #(
   .INIT(64'heffde80feffde80f)  
) LUT6_inst7863 (
   .O(to_level3[87]),
   .I0(level4_in[522]),
   .I1(level4_in[523]),
   .I2(level4_in[524]),
   .I3(level4_in[525]),
   .I4(level4_in[526]),
   .I5(level4_in[527])
);

LUT6 #(
   .INIT(64'h32b9d6a732b9d6a7)  
) LUT6_inst7864 (
   .O(to_level3[88]),
   .I0(level4_in[528]),
   .I1(level4_in[529]),
   .I2(level4_in[530]),
   .I3(level4_in[531]),
   .I4(level4_in[532]),
   .I5(level4_in[533])
);

LUT6 #(
   .INIT(64'h88fdfa4788fdfa47)  
) LUT6_inst7865 (
   .O(to_level3[89]),
   .I0(level4_in[534]),
   .I1(level4_in[535]),
   .I2(level4_in[536]),
   .I3(level4_in[537]),
   .I4(level4_in[538]),
   .I5(level4_in[539])
);

LUT6 #(
   .INIT(64'hb90da561b90da561)  
) LUT6_inst7866 (
   .O(to_level3[90]),
   .I0(level4_in[540]),
   .I1(level4_in[541]),
   .I2(level4_in[542]),
   .I3(level4_in[543]),
   .I4(level4_in[544]),
   .I5(level4_in[545])
);

LUT6 #(
   .INIT(64'h7bd1632f7bd1632f)  
) LUT6_inst7867 (
   .O(to_level3[91]),
   .I0(level4_in[546]),
   .I1(level4_in[547]),
   .I2(level4_in[548]),
   .I3(level4_in[549]),
   .I4(level4_in[550]),
   .I5(level4_in[551])
);

LUT6 #(
   .INIT(64'h1627000d1627000d)  
) LUT6_inst7868 (
   .O(to_level3[92]),
   .I0(level4_in[552]),
   .I1(level4_in[553]),
   .I2(level4_in[554]),
   .I3(level4_in[555]),
   .I4(level4_in[556]),
   .I5(level4_in[557])
);

LUT6 #(
   .INIT(64'hb4531e94b4531e94)  
) LUT6_inst7869 (
   .O(to_level3[93]),
   .I0(level4_in[558]),
   .I1(level4_in[559]),
   .I2(level4_in[560]),
   .I3(level4_in[561]),
   .I4(level4_in[562]),
   .I5(level4_in[563])
);

LUT6 #(
   .INIT(64'h18f6197918f61979)  
) LUT6_inst7870 (
   .O(to_level3[94]),
   .I0(level4_in[564]),
   .I1(level4_in[565]),
   .I2(level4_in[566]),
   .I3(level4_in[567]),
   .I4(level4_in[568]),
   .I5(level4_in[569])
);

LUT6 #(
   .INIT(64'h199141b7199141b7)  
) LUT6_inst7871 (
   .O(to_level3[95]),
   .I0(level4_in[570]),
   .I1(level4_in[571]),
   .I2(level4_in[572]),
   .I3(level4_in[573]),
   .I4(level4_in[574]),
   .I5(level4_in[575])
);

LUT6 #(
   .INIT(64'hf8715789f8715789)  
) LUT6_inst7872 (
   .O(to_level3[96]),
   .I0(level4_in[576]),
   .I1(level4_in[577]),
   .I2(level4_in[578]),
   .I3(level4_in[579]),
   .I4(level4_in[580]),
   .I5(level4_in[581])
);

LUT6 #(
   .INIT(64'h1df6f4141df6f414)  
) LUT6_inst7873 (
   .O(to_level3[97]),
   .I0(level4_in[582]),
   .I1(level4_in[583]),
   .I2(level4_in[584]),
   .I3(level4_in[585]),
   .I4(level4_in[586]),
   .I5(level4_in[587])
);

LUT6 #(
   .INIT(64'h167111d3167111d3)  
) LUT6_inst7874 (
   .O(to_level3[98]),
   .I0(level4_in[588]),
   .I1(level4_in[589]),
   .I2(level4_in[590]),
   .I3(level4_in[591]),
   .I4(level4_in[592]),
   .I5(level4_in[593])
);

LUT6 #(
   .INIT(64'h4382bd0b4382bd0b)  
) LUT6_inst7875 (
   .O(to_level3[99]),
   .I0(level4_in[594]),
   .I1(level4_in[595]),
   .I2(level4_in[596]),
   .I3(level4_in[597]),
   .I4(level4_in[598]),
   .I5(level4_in[599])
);

LUT6 #(
   .INIT(64'hcfca6956cfca6956)  
) LUT6_inst7876 (
   .O(to_level3[100]),
   .I0(level4_in[600]),
   .I1(level4_in[601]),
   .I2(level4_in[602]),
   .I3(level4_in[603]),
   .I4(level4_in[604]),
   .I5(level4_in[605])
);

LUT6 #(
   .INIT(64'h3be9273c3be9273c)  
) LUT6_inst7877 (
   .O(to_level3[101]),
   .I0(level4_in[606]),
   .I1(level4_in[607]),
   .I2(level4_in[608]),
   .I3(level4_in[609]),
   .I4(level4_in[610]),
   .I5(level4_in[611])
);

LUT6 #(
   .INIT(64'h6ca735246ca73524)  
) LUT6_inst7878 (
   .O(to_level3[102]),
   .I0(level4_in[612]),
   .I1(level4_in[613]),
   .I2(level4_in[614]),
   .I3(level4_in[615]),
   .I4(level4_in[616]),
   .I5(level4_in[617])
);

LUT6 #(
   .INIT(64'hcc77a150cc77a150)  
) LUT6_inst7879 (
   .O(to_level3[103]),
   .I0(level4_in[618]),
   .I1(level4_in[619]),
   .I2(level4_in[620]),
   .I3(level4_in[621]),
   .I4(level4_in[622]),
   .I5(level4_in[623])
);

LUT6 #(
   .INIT(64'ha87198bfa87198bf)  
) LUT6_inst7880 (
   .O(to_level3[104]),
   .I0(level4_in[624]),
   .I1(level4_in[625]),
   .I2(level4_in[626]),
   .I3(level4_in[627]),
   .I4(level4_in[628]),
   .I5(level4_in[629])
);

LUT6 #(
   .INIT(64'hfc7dc213fc7dc213)  
) LUT6_inst7881 (
   .O(to_level3[105]),
   .I0(level4_in[630]),
   .I1(level4_in[631]),
   .I2(level4_in[632]),
   .I3(level4_in[633]),
   .I4(level4_in[634]),
   .I5(level4_in[635])
);

LUT6 #(
   .INIT(64'h9e3dcef29e3dcef2)  
) LUT6_inst7882 (
   .O(to_level3[106]),
   .I0(level4_in[636]),
   .I1(level4_in[637]),
   .I2(level4_in[638]),
   .I3(level4_in[639]),
   .I4(level4_in[640]),
   .I5(level4_in[641])
);

LUT6 #(
   .INIT(64'h6e5d78006e5d7800)  
) LUT6_inst7883 (
   .O(to_level3[107]),
   .I0(level4_in[642]),
   .I1(level4_in[643]),
   .I2(level4_in[644]),
   .I3(level4_in[645]),
   .I4(level4_in[646]),
   .I5(level4_in[647])
);

LUT6 #(
   .INIT(64'hcd631598cd631598)  
) LUT6_inst7884 (
   .O(to_level3[108]),
   .I0(level4_in[648]),
   .I1(level4_in[649]),
   .I2(level4_in[650]),
   .I3(level4_in[651]),
   .I4(level4_in[652]),
   .I5(level4_in[653])
);

LUT6 #(
   .INIT(64'h2890cfe72890cfe7)  
) LUT6_inst7885 (
   .O(to_level3[109]),
   .I0(level4_in[654]),
   .I1(level4_in[655]),
   .I2(level4_in[656]),
   .I3(level4_in[657]),
   .I4(level4_in[658]),
   .I5(level4_in[659])
);

LUT6 #(
   .INIT(64'h873697d9873697d9)  
) LUT6_inst7886 (
   .O(to_level3[110]),
   .I0(level4_in[660]),
   .I1(level4_in[661]),
   .I2(level4_in[662]),
   .I3(level4_in[663]),
   .I4(level4_in[664]),
   .I5(level4_in[665])
);

LUT6 #(
   .INIT(64'h2fd16dfb2fd16dfb)  
) LUT6_inst7887 (
   .O(to_level3[111]),
   .I0(level4_in[666]),
   .I1(level4_in[667]),
   .I2(level4_in[668]),
   .I3(level4_in[669]),
   .I4(level4_in[670]),
   .I5(level4_in[671])
);

LUT6 #(
   .INIT(64'hbcb692f6bcb692f6)  
) LUT6_inst7888 (
   .O(to_level3[112]),
   .I0(level4_in[672]),
   .I1(level4_in[673]),
   .I2(level4_in[674]),
   .I3(level4_in[675]),
   .I4(level4_in[676]),
   .I5(level4_in[677])
);

LUT6 #(
   .INIT(64'hff69abc9ff69abc9)  
) LUT6_inst7889 (
   .O(to_level3[113]),
   .I0(level4_in[678]),
   .I1(level4_in[679]),
   .I2(level4_in[680]),
   .I3(level4_in[681]),
   .I4(level4_in[682]),
   .I5(level4_in[683])
);

LUT6 #(
   .INIT(64'h3d01372b3d01372b)  
) LUT6_inst7890 (
   .O(to_level3[114]),
   .I0(level4_in[684]),
   .I1(level4_in[685]),
   .I2(level4_in[686]),
   .I3(level4_in[687]),
   .I4(level4_in[688]),
   .I5(level4_in[689])
);

LUT6 #(
   .INIT(64'h3ad85d543ad85d54)  
) LUT6_inst7891 (
   .O(to_level3[115]),
   .I0(level4_in[690]),
   .I1(level4_in[691]),
   .I2(level4_in[692]),
   .I3(level4_in[693]),
   .I4(level4_in[694]),
   .I5(level4_in[695])
);

LUT6 #(
   .INIT(64'hee3160b3ee3160b3)  
) LUT6_inst7892 (
   .O(to_level3[116]),
   .I0(level4_in[696]),
   .I1(level4_in[697]),
   .I2(level4_in[698]),
   .I3(level4_in[699]),
   .I4(level4_in[700]),
   .I5(level4_in[701])
);

LUT6 #(
   .INIT(64'h8a8f719e8a8f719e)  
) LUT6_inst7893 (
   .O(to_level3[117]),
   .I0(level4_in[702]),
   .I1(level4_in[703]),
   .I2(level4_in[704]),
   .I3(level4_in[705]),
   .I4(level4_in[706]),
   .I5(level4_in[707])
);

LUT6 #(
   .INIT(64'hcca7ea3bcca7ea3b)  
) LUT6_inst7894 (
   .O(to_level3[118]),
   .I0(level4_in[708]),
   .I1(level4_in[709]),
   .I2(level4_in[710]),
   .I3(level4_in[711]),
   .I4(level4_in[712]),
   .I5(level4_in[713])
);

LUT6 #(
   .INIT(64'hd499c403d499c403)  
) LUT6_inst7895 (
   .O(to_level3[119]),
   .I0(level4_in[714]),
   .I1(level4_in[715]),
   .I2(level4_in[716]),
   .I3(level4_in[717]),
   .I4(level4_in[718]),
   .I5(level4_in[719])
);

LUT6 #(
   .INIT(64'h15e3929015e39290)  
) LUT6_inst7896 (
   .O(to_level3[120]),
   .I0(level4_in[720]),
   .I1(level4_in[721]),
   .I2(level4_in[722]),
   .I3(level4_in[723]),
   .I4(level4_in[724]),
   .I5(level4_in[725])
);

LUT6 #(
   .INIT(64'h5a152f325a152f32)  
) LUT6_inst7897 (
   .O(to_level3[121]),
   .I0(level4_in[726]),
   .I1(level4_in[727]),
   .I2(level4_in[728]),
   .I3(level4_in[729]),
   .I4(level4_in[730]),
   .I5(level4_in[731])
);

LUT6 #(
   .INIT(64'h88307b3488307b34)  
) LUT6_inst7898 (
   .O(to_level3[122]),
   .I0(level4_in[732]),
   .I1(level4_in[733]),
   .I2(level4_in[734]),
   .I3(level4_in[735]),
   .I4(level4_in[736]),
   .I5(level4_in[737])
);

LUT6 #(
   .INIT(64'h9bf3cfc69bf3cfc6)  
) LUT6_inst7899 (
   .O(to_level3[123]),
   .I0(level4_in[738]),
   .I1(level4_in[739]),
   .I2(level4_in[740]),
   .I3(level4_in[741]),
   .I4(level4_in[742]),
   .I5(level4_in[743])
);

LUT6 #(
   .INIT(64'h393bcb4f393bcb4f)  
) LUT6_inst7900 (
   .O(to_level3[124]),
   .I0(level4_in[744]),
   .I1(level4_in[745]),
   .I2(level4_in[746]),
   .I3(level4_in[747]),
   .I4(level4_in[748]),
   .I5(level4_in[749])
);

LUT6 #(
   .INIT(64'hd8691172d8691172)  
) LUT6_inst7901 (
   .O(to_level3[125]),
   .I0(level4_in[750]),
   .I1(level4_in[751]),
   .I2(level4_in[752]),
   .I3(level4_in[753]),
   .I4(level4_in[754]),
   .I5(level4_in[755])
);

LUT6 #(
   .INIT(64'he0606564e0606564)  
) LUT6_inst7902 (
   .O(to_level3[126]),
   .I0(level4_in[756]),
   .I1(level4_in[757]),
   .I2(level4_in[758]),
   .I3(level4_in[759]),
   .I4(level4_in[760]),
   .I5(level4_in[761])
);

LUT6 #(
   .INIT(64'h04f22b6c04f22b6c)  
) LUT6_inst7903 (
   .O(to_level3[127]),
   .I0(level4_in[762]),
   .I1(level4_in[763]),
   .I2(level4_in[764]),
   .I3(level4_in[765]),
   .I4(level4_in[766]),
   .I5(level4_in[767])
);

LUT6 #(
   .INIT(64'h4e037f4a4e037f4a)  
) LUT6_inst7904 (
   .O(to_level3[128]),
   .I0(level4_in[768]),
   .I1(level4_in[769]),
   .I2(level4_in[770]),
   .I3(level4_in[771]),
   .I4(level4_in[772]),
   .I5(level4_in[773])
);

LUT6 #(
   .INIT(64'hd7768503d7768503)  
) LUT6_inst7905 (
   .O(to_level3[129]),
   .I0(level4_in[774]),
   .I1(level4_in[775]),
   .I2(level4_in[776]),
   .I3(level4_in[777]),
   .I4(level4_in[778]),
   .I5(level4_in[779])
);

LUT6 #(
   .INIT(64'h9a59e3ac9a59e3ac)  
) LUT6_inst7906 (
   .O(to_level3[130]),
   .I0(level4_in[780]),
   .I1(level4_in[781]),
   .I2(level4_in[782]),
   .I3(level4_in[783]),
   .I4(level4_in[784]),
   .I5(level4_in[785])
);

LUT6 #(
   .INIT(64'hfe42767cfe42767c)  
) LUT6_inst7907 (
   .O(to_level3[131]),
   .I0(level4_in[786]),
   .I1(level4_in[787]),
   .I2(level4_in[788]),
   .I3(level4_in[789]),
   .I4(level4_in[790]),
   .I5(level4_in[791])
);

LUT6 #(
   .INIT(64'h7da2723c7da2723c)  
) LUT6_inst7908 (
   .O(to_level3[132]),
   .I0(level4_in[792]),
   .I1(level4_in[793]),
   .I2(level4_in[794]),
   .I3(level4_in[795]),
   .I4(level4_in[796]),
   .I5(level4_in[797])
);

LUT6 #(
   .INIT(64'h22642a6c22642a6c)  
) LUT6_inst7909 (
   .O(to_level3[133]),
   .I0(level4_in[798]),
   .I1(level4_in[799]),
   .I2(level4_in[800]),
   .I3(level4_in[801]),
   .I4(level4_in[802]),
   .I5(level4_in[803])
);

LUT6 #(
   .INIT(64'h5585c2f45585c2f4)  
) LUT6_inst7910 (
   .O(to_level3[134]),
   .I0(level4_in[804]),
   .I1(level4_in[805]),
   .I2(level4_in[806]),
   .I3(level4_in[807]),
   .I4(level4_in[808]),
   .I5(level4_in[809])
);

LUT6 #(
   .INIT(64'h51c7bf8151c7bf81)  
) LUT6_inst7911 (
   .O(to_level3[135]),
   .I0(level4_in[810]),
   .I1(level4_in[811]),
   .I2(level4_in[812]),
   .I3(level4_in[813]),
   .I4(level4_in[814]),
   .I5(level4_in[815])
);

LUT6 #(
   .INIT(64'h29ca885829ca8858)  
) LUT6_inst7912 (
   .O(to_level3[136]),
   .I0(level4_in[816]),
   .I1(level4_in[817]),
   .I2(level4_in[818]),
   .I3(level4_in[819]),
   .I4(level4_in[820]),
   .I5(level4_in[821])
);

LUT6 #(
   .INIT(64'hcaf86e3acaf86e3a)  
) LUT6_inst7913 (
   .O(to_level3[137]),
   .I0(level4_in[822]),
   .I1(level4_in[823]),
   .I2(level4_in[824]),
   .I3(level4_in[825]),
   .I4(level4_in[826]),
   .I5(level4_in[827])
);

LUT6 #(
   .INIT(64'h18c0903718c09037)  
) LUT6_inst7914 (
   .O(to_level3[138]),
   .I0(level4_in[828]),
   .I1(level4_in[829]),
   .I2(level4_in[830]),
   .I3(level4_in[831]),
   .I4(level4_in[832]),
   .I5(level4_in[833])
);

LUT6 #(
   .INIT(64'h3ad5b4073ad5b407)  
) LUT6_inst7915 (
   .O(to_level3[139]),
   .I0(level4_in[834]),
   .I1(level4_in[835]),
   .I2(level4_in[836]),
   .I3(level4_in[837]),
   .I4(level4_in[838]),
   .I5(level4_in[839])
);

LUT6 #(
   .INIT(64'hee7c0712ee7c0712)  
) LUT6_inst7916 (
   .O(to_level3[140]),
   .I0(level4_in[840]),
   .I1(level4_in[841]),
   .I2(level4_in[842]),
   .I3(level4_in[843]),
   .I4(level4_in[844]),
   .I5(level4_in[845])
);

LUT6 #(
   .INIT(64'hed2270bded2270bd)  
) LUT6_inst7917 (
   .O(to_level3[141]),
   .I0(level4_in[846]),
   .I1(level4_in[847]),
   .I2(level4_in[848]),
   .I3(level4_in[849]),
   .I4(level4_in[850]),
   .I5(level4_in[851])
);

LUT6 #(
   .INIT(64'he37f6826e37f6826)  
) LUT6_inst7918 (
   .O(to_level3[142]),
   .I0(level4_in[852]),
   .I1(level4_in[853]),
   .I2(level4_in[854]),
   .I3(level4_in[855]),
   .I4(level4_in[856]),
   .I5(level4_in[857])
);

LUT6 #(
   .INIT(64'hd23ae653d23ae653)  
) LUT6_inst7919 (
   .O(to_level3[143]),
   .I0(level4_in[858]),
   .I1(level4_in[859]),
   .I2(level4_in[860]),
   .I3(level4_in[861]),
   .I4(level4_in[862]),
   .I5(level4_in[863])
);

LUT6 #(
   .INIT(64'h4033c4864033c486)  
) LUT6_inst7920 (
   .O(to_level3[144]),
   .I0(level4_in[864]),
   .I1(level4_in[865]),
   .I2(level4_in[866]),
   .I3(level4_in[867]),
   .I4(level4_in[868]),
   .I5(level4_in[869])
);

LUT6 #(
   .INIT(64'hee80005bee80005b)  
) LUT6_inst7921 (
   .O(to_level3[145]),
   .I0(level4_in[870]),
   .I1(level4_in[871]),
   .I2(level4_in[872]),
   .I3(level4_in[873]),
   .I4(level4_in[874]),
   .I5(level4_in[875])
);

LUT6 #(
   .INIT(64'h0e24fa550e24fa55)  
) LUT6_inst7922 (
   .O(to_level3[146]),
   .I0(level4_in[876]),
   .I1(level4_in[877]),
   .I2(level4_in[878]),
   .I3(level4_in[879]),
   .I4(level4_in[880]),
   .I5(level4_in[881])
);

LUT6 #(
   .INIT(64'hba2164cdba2164cd)  
) LUT6_inst7923 (
   .O(to_level3[147]),
   .I0(level4_in[882]),
   .I1(level4_in[883]),
   .I2(level4_in[884]),
   .I3(level4_in[885]),
   .I4(level4_in[886]),
   .I5(level4_in[887])
);

LUT6 #(
   .INIT(64'h2be985d12be985d1)  
) LUT6_inst7924 (
   .O(to_level3[148]),
   .I0(level4_in[888]),
   .I1(level4_in[889]),
   .I2(level4_in[890]),
   .I3(level4_in[891]),
   .I4(level4_in[892]),
   .I5(level4_in[893])
);

LUT6 #(
   .INIT(64'h2bdb8f4e2bdb8f4e)  
) LUT6_inst7925 (
   .O(to_level3[149]),
   .I0(level4_in[894]),
   .I1(level4_in[895]),
   .I2(level4_in[896]),
   .I3(level4_in[897]),
   .I4(level4_in[898]),
   .I5(level4_in[899])
);

LUT6 #(
   .INIT(64'hea1ed37cea1ed37c)  
) LUT6_inst7926 (
   .O(to_level3[150]),
   .I0(level4_in[900]),
   .I1(level4_in[901]),
   .I2(level4_in[902]),
   .I3(level4_in[903]),
   .I4(level4_in[904]),
   .I5(level4_in[905])
);

LUT6 #(
   .INIT(64'h4b24de5f4b24de5f)  
) LUT6_inst7927 (
   .O(to_level3[151]),
   .I0(level4_in[906]),
   .I1(level4_in[907]),
   .I2(level4_in[908]),
   .I3(level4_in[909]),
   .I4(level4_in[910]),
   .I5(level4_in[911])
);

LUT6 #(
   .INIT(64'h85e2710785e27107)  
) LUT6_inst7928 (
   .O(to_level3[152]),
   .I0(level4_in[912]),
   .I1(level4_in[913]),
   .I2(level4_in[914]),
   .I3(level4_in[915]),
   .I4(level4_in[916]),
   .I5(level4_in[917])
);

LUT6 #(
   .INIT(64'h777a0c84777a0c84)  
) LUT6_inst7929 (
   .O(to_level3[153]),
   .I0(level4_in[918]),
   .I1(level4_in[919]),
   .I2(level4_in[920]),
   .I3(level4_in[921]),
   .I4(level4_in[922]),
   .I5(level4_in[923])
);

LUT6 #(
   .INIT(64'hf0b912eaf0b912ea)  
) LUT6_inst7930 (
   .O(to_level3[154]),
   .I0(level4_in[924]),
   .I1(level4_in[925]),
   .I2(level4_in[926]),
   .I3(level4_in[927]),
   .I4(level4_in[928]),
   .I5(level4_in[929])
);

LUT6 #(
   .INIT(64'h6537b64c6537b64c)  
) LUT6_inst7931 (
   .O(to_level3[155]),
   .I0(level4_in[930]),
   .I1(level4_in[931]),
   .I2(level4_in[932]),
   .I3(level4_in[933]),
   .I4(level4_in[934]),
   .I5(level4_in[935])
);

LUT6 #(
   .INIT(64'h8bd09e008bd09e00)  
) LUT6_inst7932 (
   .O(to_level3[156]),
   .I0(level4_in[936]),
   .I1(level4_in[937]),
   .I2(level4_in[938]),
   .I3(level4_in[939]),
   .I4(level4_in[940]),
   .I5(level4_in[941])
);

LUT6 #(
   .INIT(64'h701f3a4f701f3a4f)  
) LUT6_inst7933 (
   .O(to_level3[157]),
   .I0(level4_in[942]),
   .I1(level4_in[943]),
   .I2(level4_in[944]),
   .I3(level4_in[945]),
   .I4(level4_in[946]),
   .I5(level4_in[947])
);

LUT6 #(
   .INIT(64'h120d6710120d6710)  
) LUT6_inst7934 (
   .O(to_level3[158]),
   .I0(level4_in[948]),
   .I1(level4_in[949]),
   .I2(level4_in[950]),
   .I3(level4_in[951]),
   .I4(level4_in[952]),
   .I5(level4_in[953])
);

LUT6 #(
   .INIT(64'hc3da1d77c3da1d77)  
) LUT6_inst7935 (
   .O(to_level3[159]),
   .I0(level4_in[954]),
   .I1(level4_in[955]),
   .I2(level4_in[956]),
   .I3(level4_in[957]),
   .I4(level4_in[958]),
   .I5(level4_in[959])
);

LUT6 #(
   .INIT(64'h62e175a862e175a8)  
) LUT6_inst7936 (
   .O(to_level3[160]),
   .I0(level4_in[960]),
   .I1(level4_in[961]),
   .I2(level4_in[962]),
   .I3(level4_in[963]),
   .I4(level4_in[964]),
   .I5(level4_in[965])
);

LUT6 #(
   .INIT(64'h3eca89583eca8958)  
) LUT6_inst7937 (
   .O(to_level3[161]),
   .I0(level4_in[966]),
   .I1(level4_in[967]),
   .I2(level4_in[968]),
   .I3(level4_in[969]),
   .I4(level4_in[970]),
   .I5(level4_in[971])
);

LUT6 #(
   .INIT(64'h1b3e51451b3e5145)  
) LUT6_inst7938 (
   .O(to_level3[162]),
   .I0(level4_in[972]),
   .I1(level4_in[973]),
   .I2(level4_in[974]),
   .I3(level4_in[975]),
   .I4(level4_in[976]),
   .I5(level4_in[977])
);

LUT6 #(
   .INIT(64'h97ab95cc97ab95cc)  
) LUT6_inst7939 (
   .O(to_level3[163]),
   .I0(level4_in[978]),
   .I1(level4_in[979]),
   .I2(level4_in[980]),
   .I3(level4_in[981]),
   .I4(level4_in[982]),
   .I5(level4_in[983])
);

LUT6 #(
   .INIT(64'haba16ea0aba16ea0)  
) LUT6_inst7940 (
   .O(to_level3[164]),
   .I0(level4_in[984]),
   .I1(level4_in[985]),
   .I2(level4_in[986]),
   .I3(level4_in[987]),
   .I4(level4_in[988]),
   .I5(level4_in[989])
);

LUT6 #(
   .INIT(64'hce070d9ace070d9a)  
) LUT6_inst7941 (
   .O(to_level3[165]),
   .I0(level4_in[990]),
   .I1(level4_in[991]),
   .I2(level4_in[992]),
   .I3(level4_in[993]),
   .I4(level4_in[994]),
   .I5(level4_in[995])
);

LUT6 #(
   .INIT(64'hec1de1b4ec1de1b4)  
) LUT6_inst7942 (
   .O(to_level3[166]),
   .I0(level4_in[996]),
   .I1(level4_in[997]),
   .I2(level4_in[998]),
   .I3(level4_in[999]),
   .I4(level4_in[1000]),
   .I5(level4_in[1001])
);

LUT6 #(
   .INIT(64'hfc049016fc049016)  
) LUT6_inst7943 (
   .O(to_level3[167]),
   .I0(level4_in[1002]),
   .I1(level4_in[1003]),
   .I2(level4_in[1004]),
   .I3(level4_in[1005]),
   .I4(level4_in[1006]),
   .I5(level4_in[1007])
);

LUT6 #(
   .INIT(64'hdbe530acdbe530ac)  
) LUT6_inst7944 (
   .O(to_level3[168]),
   .I0(level4_in[1008]),
   .I1(level4_in[1009]),
   .I2(level4_in[1010]),
   .I3(level4_in[1011]),
   .I4(level4_in[1012]),
   .I5(level4_in[1013])
);

LUT6 #(
   .INIT(64'h78cd47c678cd47c6)  
) LUT6_inst7945 (
   .O(to_level3[169]),
   .I0(level4_in[1014]),
   .I1(level4_in[1015]),
   .I2(level4_in[1016]),
   .I3(level4_in[1017]),
   .I4(level4_in[1018]),
   .I5(level4_in[1019])
);

LUT6 #(
   .INIT(64'hd1d7c85cd1d7c85c)  
) LUT6_inst7946 (
   .O(to_level3[170]),
   .I0(level4_in[1020]),
   .I1(level4_in[1021]),
   .I2(level4_in[1022]),
   .I3(level4_in[1023]),
   .I4(level4_in[1024]),
   .I5(level4_in[1025])
);

LUT6 #(
   .INIT(64'h357c320b357c320b)  
) LUT6_inst7947 (
   .O(to_level3[171]),
   .I0(level4_in[1026]),
   .I1(level4_in[1027]),
   .I2(level4_in[1028]),
   .I3(level4_in[1029]),
   .I4(level4_in[1030]),
   .I5(level4_in[1031])
);

LUT6 #(
   .INIT(64'hc1237638c1237638)  
) LUT6_inst7948 (
   .O(to_level3[172]),
   .I0(level4_in[1032]),
   .I1(level4_in[1033]),
   .I2(level4_in[1034]),
   .I3(level4_in[1035]),
   .I4(level4_in[1036]),
   .I5(level4_in[1037])
);

LUT6 #(
   .INIT(64'hab62cc80ab62cc80)  
) LUT6_inst7949 (
   .O(to_level3[173]),
   .I0(level4_in[1038]),
   .I1(level4_in[1039]),
   .I2(level4_in[1040]),
   .I3(level4_in[1041]),
   .I4(level4_in[1042]),
   .I5(level4_in[1043])
);

LUT6 #(
   .INIT(64'h2fe676512fe67651)  
) LUT6_inst7950 (
   .O(to_level3[174]),
   .I0(level4_in[1044]),
   .I1(level4_in[1045]),
   .I2(level4_in[1046]),
   .I3(level4_in[1047]),
   .I4(level4_in[1048]),
   .I5(level4_in[1049])
);

LUT6 #(
   .INIT(64'hfe060d30fe060d30)  
) LUT6_inst7951 (
   .O(to_level3[175]),
   .I0(level4_in[1050]),
   .I1(level4_in[1051]),
   .I2(level4_in[1052]),
   .I3(level4_in[1053]),
   .I4(level4_in[1054]),
   .I5(level4_in[1055])
);

LUT6 #(
   .INIT(64'h570979c0570979c0)  
) LUT6_inst7952 (
   .O(to_level3[176]),
   .I0(level4_in[1056]),
   .I1(level4_in[1057]),
   .I2(level4_in[1058]),
   .I3(level4_in[1059]),
   .I4(level4_in[1060]),
   .I5(level4_in[1061])
);

LUT6 #(
   .INIT(64'hff777e61ff777e61)  
) LUT6_inst7953 (
   .O(to_level3[177]),
   .I0(level4_in[1062]),
   .I1(level4_in[1063]),
   .I2(level4_in[1064]),
   .I3(level4_in[1065]),
   .I4(level4_in[1066]),
   .I5(level4_in[1067])
);

LUT6 #(
   .INIT(64'h6042ee7c6042ee7c)  
) LUT6_inst7954 (
   .O(to_level3[178]),
   .I0(level4_in[1068]),
   .I1(level4_in[1069]),
   .I2(level4_in[1070]),
   .I3(level4_in[1071]),
   .I4(level4_in[1072]),
   .I5(level4_in[1073])
);

LUT6 #(
   .INIT(64'hbd216610bd216610)  
) LUT6_inst7955 (
   .O(to_level3[179]),
   .I0(level4_in[1074]),
   .I1(level4_in[1075]),
   .I2(level4_in[1076]),
   .I3(level4_in[1077]),
   .I4(level4_in[1078]),
   .I5(level4_in[1079])
);

LUT6 #(
   .INIT(64'h9da502a89da502a8)  
) LUT6_inst7956 (
   .O(to_level3[180]),
   .I0(level4_in[1080]),
   .I1(level4_in[1081]),
   .I2(level4_in[1082]),
   .I3(level4_in[1083]),
   .I4(level4_in[1084]),
   .I5(level4_in[1085])
);

LUT6 #(
   .INIT(64'h254af2e8254af2e8)  
) LUT6_inst7957 (
   .O(to_level3[181]),
   .I0(level4_in[1086]),
   .I1(level4_in[1087]),
   .I2(level4_in[1088]),
   .I3(level4_in[1089]),
   .I4(level4_in[1090]),
   .I5(level4_in[1091])
);

LUT6 #(
   .INIT(64'h2b5cd2aa2b5cd2aa)  
) LUT6_inst7958 (
   .O(to_level3[182]),
   .I0(level4_in[1092]),
   .I1(level4_in[1093]),
   .I2(level4_in[1094]),
   .I3(level4_in[1095]),
   .I4(level4_in[1096]),
   .I5(level4_in[1097])
);

LUT6 #(
   .INIT(64'h6db9513d6db9513d)  
) LUT6_inst7959 (
   .O(to_level3[183]),
   .I0(level4_in[1098]),
   .I1(level4_in[1099]),
   .I2(level4_in[1100]),
   .I3(level4_in[1101]),
   .I4(level4_in[1102]),
   .I5(level4_in[1103])
);

LUT6 #(
   .INIT(64'hcbb0ad37cbb0ad37)  
) LUT6_inst7960 (
   .O(to_level3[184]),
   .I0(level4_in[1104]),
   .I1(level4_in[1105]),
   .I2(level4_in[1106]),
   .I3(level4_in[1107]),
   .I4(level4_in[1108]),
   .I5(level4_in[1109])
);

LUT6 #(
   .INIT(64'h0745ad570745ad57)  
) LUT6_inst7961 (
   .O(to_level3[185]),
   .I0(level4_in[1110]),
   .I1(level4_in[1111]),
   .I2(level4_in[1112]),
   .I3(level4_in[1113]),
   .I4(level4_in[1114]),
   .I5(level4_in[1115])
);

LUT6 #(
   .INIT(64'h4cd4a59c4cd4a59c)  
) LUT6_inst7962 (
   .O(to_level3[186]),
   .I0(level4_in[1116]),
   .I1(level4_in[1117]),
   .I2(level4_in[1118]),
   .I3(level4_in[1119]),
   .I4(level4_in[1120]),
   .I5(level4_in[1121])
);

LUT6 #(
   .INIT(64'hf3d774cbf3d774cb)  
) LUT6_inst7963 (
   .O(to_level3[187]),
   .I0(level4_in[1122]),
   .I1(level4_in[1123]),
   .I2(level4_in[1124]),
   .I3(level4_in[1125]),
   .I4(level4_in[1126]),
   .I5(level4_in[1127])
);

LUT6 #(
   .INIT(64'h441f8499441f8499)  
) LUT6_inst7964 (
   .O(to_level3[188]),
   .I0(level4_in[1128]),
   .I1(level4_in[1129]),
   .I2(level4_in[1130]),
   .I3(level4_in[1131]),
   .I4(level4_in[1132]),
   .I5(level4_in[1133])
);

LUT6 #(
   .INIT(64'hb55f8305b55f8305)  
) LUT6_inst7965 (
   .O(to_level3[189]),
   .I0(level4_in[1134]),
   .I1(level4_in[1135]),
   .I2(level4_in[1136]),
   .I3(level4_in[1137]),
   .I4(level4_in[1138]),
   .I5(level4_in[1139])
);

LUT6 #(
   .INIT(64'hb9e65bd9b9e65bd9)  
) LUT6_inst7966 (
   .O(to_level3[190]),
   .I0(level4_in[1140]),
   .I1(level4_in[1141]),
   .I2(level4_in[1142]),
   .I3(level4_in[1143]),
   .I4(level4_in[1144]),
   .I5(level4_in[1145])
);

LUT6 #(
   .INIT(64'h7f3113137f311313)  
) LUT6_inst7967 (
   .O(to_level3[191]),
   .I0(level4_in[1146]),
   .I1(level4_in[1147]),
   .I2(level4_in[1148]),
   .I3(level4_in[1149]),
   .I4(level4_in[1150]),
   .I5(level4_in[1151])
);

LUT6 #(
   .INIT(64'h903593ce903593ce)  
) LUT6_inst7968 (
   .O(to_level3[192]),
   .I0(level4_in[1152]),
   .I1(level4_in[1153]),
   .I2(level4_in[1154]),
   .I3(level4_in[1155]),
   .I4(level4_in[1156]),
   .I5(level4_in[1157])
);

LUT6 #(
   .INIT(64'h5bfb2c2d5bfb2c2d)  
) LUT6_inst7969 (
   .O(to_level3[193]),
   .I0(level4_in[1158]),
   .I1(level4_in[1159]),
   .I2(level4_in[1160]),
   .I3(level4_in[1161]),
   .I4(level4_in[1162]),
   .I5(level4_in[1163])
);

LUT6 #(
   .INIT(64'ha12b86faa12b86fa)  
) LUT6_inst7970 (
   .O(to_level3[194]),
   .I0(level4_in[1164]),
   .I1(level4_in[1165]),
   .I2(level4_in[1166]),
   .I3(level4_in[1167]),
   .I4(level4_in[1168]),
   .I5(level4_in[1169])
);

LUT6 #(
   .INIT(64'h46e7343246e73432)  
) LUT6_inst7971 (
   .O(to_level3[195]),
   .I0(level4_in[1170]),
   .I1(level4_in[1171]),
   .I2(level4_in[1172]),
   .I3(level4_in[1173]),
   .I4(level4_in[1174]),
   .I5(level4_in[1175])
);

LUT6 #(
   .INIT(64'h83c146ea83c146ea)  
) LUT6_inst7972 (
   .O(to_level3[196]),
   .I0(level4_in[1176]),
   .I1(level4_in[1177]),
   .I2(level4_in[1178]),
   .I3(level4_in[1179]),
   .I4(level4_in[1180]),
   .I5(level4_in[1181])
);

LUT6 #(
   .INIT(64'h5adadbc05adadbc0)  
) LUT6_inst7973 (
   .O(to_level3[197]),
   .I0(level4_in[1182]),
   .I1(level4_in[1183]),
   .I2(level4_in[1184]),
   .I3(level4_in[1185]),
   .I4(level4_in[1186]),
   .I5(level4_in[1187])
);

LUT6 #(
   .INIT(64'h3987ab6e3987ab6e)  
) LUT6_inst7974 (
   .O(to_level3[198]),
   .I0(level4_in[1188]),
   .I1(level4_in[1189]),
   .I2(level4_in[1190]),
   .I3(level4_in[1191]),
   .I4(level4_in[1192]),
   .I5(level4_in[1193])
);

LUT6 #(
   .INIT(64'hc7676f3bc7676f3b)  
) LUT6_inst7975 (
   .O(to_level3[199]),
   .I0(level4_in[1194]),
   .I1(level4_in[1195]),
   .I2(level4_in[1196]),
   .I3(level4_in[1197]),
   .I4(level4_in[1198]),
   .I5(level4_in[1199])
);

LUT6 #(
   .INIT(64'hd80daab7d80daab7)  
) LUT6_inst7976 (
   .O(to_level3[200]),
   .I0(level4_in[1200]),
   .I1(level4_in[1201]),
   .I2(level4_in[1202]),
   .I3(level4_in[1203]),
   .I4(level4_in[1204]),
   .I5(level4_in[1205])
);

LUT6 #(
   .INIT(64'h3e168ae03e168ae0)  
) LUT6_inst7977 (
   .O(to_level3[201]),
   .I0(level4_in[1206]),
   .I1(level4_in[1207]),
   .I2(level4_in[1208]),
   .I3(level4_in[1209]),
   .I4(level4_in[1210]),
   .I5(level4_in[1211])
);

LUT6 #(
   .INIT(64'hf27c808af27c808a)  
) LUT6_inst7978 (
   .O(to_level3[202]),
   .I0(level4_in[1212]),
   .I1(level4_in[1213]),
   .I2(level4_in[1214]),
   .I3(level4_in[1215]),
   .I4(level4_in[1216]),
   .I5(level4_in[1217])
);

LUT6 #(
   .INIT(64'h997dfa15997dfa15)  
) LUT6_inst7979 (
   .O(to_level3[203]),
   .I0(level4_in[1218]),
   .I1(level4_in[1219]),
   .I2(level4_in[1220]),
   .I3(level4_in[1221]),
   .I4(level4_in[1222]),
   .I5(level4_in[1223])
);

LUT6 #(
   .INIT(64'h9281bc139281bc13)  
) LUT6_inst7980 (
   .O(to_level3[204]),
   .I0(level4_in[1224]),
   .I1(level4_in[1225]),
   .I2(level4_in[1226]),
   .I3(level4_in[1227]),
   .I4(level4_in[1228]),
   .I5(level4_in[1229])
);

LUT6 #(
   .INIT(64'haa4ade68aa4ade68)  
) LUT6_inst7981 (
   .O(to_level3[205]),
   .I0(level4_in[1230]),
   .I1(level4_in[1231]),
   .I2(level4_in[1232]),
   .I3(level4_in[1233]),
   .I4(level4_in[1234]),
   .I5(level4_in[1235])
);

LUT6 #(
   .INIT(64'h73b7fa9573b7fa95)  
) LUT6_inst7982 (
   .O(to_level3[206]),
   .I0(level4_in[1236]),
   .I1(level4_in[1237]),
   .I2(level4_in[1238]),
   .I3(level4_in[1239]),
   .I4(level4_in[1240]),
   .I5(level4_in[1241])
);

LUT6 #(
   .INIT(64'h8d8ecc998d8ecc99)  
) LUT6_inst7983 (
   .O(to_level3[207]),
   .I0(level4_in[1242]),
   .I1(level4_in[1243]),
   .I2(level4_in[1244]),
   .I3(level4_in[1245]),
   .I4(level4_in[1246]),
   .I5(level4_in[1247])
);

LUT6 #(
   .INIT(64'hfd41cacffd41cacf)  
) LUT6_inst7984 (
   .O(to_level3[208]),
   .I0(level4_in[1248]),
   .I1(level4_in[1249]),
   .I2(level4_in[1250]),
   .I3(level4_in[1251]),
   .I4(level4_in[1252]),
   .I5(level4_in[1253])
);

LUT6 #(
   .INIT(64'h6b790f146b790f14)  
) LUT6_inst7985 (
   .O(to_level3[209]),
   .I0(level4_in[1254]),
   .I1(level4_in[1255]),
   .I2(level4_in[1256]),
   .I3(level4_in[1257]),
   .I4(level4_in[1258]),
   .I5(level4_in[1259])
);

LUT6 #(
   .INIT(64'h6d842dac6d842dac)  
) LUT6_inst7986 (
   .O(to_level3[210]),
   .I0(level4_in[1260]),
   .I1(level4_in[1261]),
   .I2(level4_in[1262]),
   .I3(level4_in[1263]),
   .I4(level4_in[1264]),
   .I5(level4_in[1265])
);

LUT6 #(
   .INIT(64'h5b107e995b107e99)  
) LUT6_inst7987 (
   .O(to_level3[211]),
   .I0(level4_in[1266]),
   .I1(level4_in[1267]),
   .I2(level4_in[1268]),
   .I3(level4_in[1269]),
   .I4(level4_in[1270]),
   .I5(level4_in[1271])
);

LUT6 #(
   .INIT(64'h3ebf00433ebf0043)  
) LUT6_inst7988 (
   .O(to_level3[212]),
   .I0(level4_in[1272]),
   .I1(level4_in[1273]),
   .I2(level4_in[1274]),
   .I3(level4_in[1275]),
   .I4(level4_in[1276]),
   .I5(level4_in[1277])
);

LUT6 #(
   .INIT(64'h85f8f6b785f8f6b7)  
) LUT6_inst7989 (
   .O(to_level3[213]),
   .I0(level4_in[1278]),
   .I1(level4_in[1279]),
   .I2(level4_in[1280]),
   .I3(level4_in[1281]),
   .I4(level4_in[1282]),
   .I5(level4_in[1283])
);

LUT6 #(
   .INIT(64'hc87912e0c87912e0)  
) LUT6_inst7990 (
   .O(to_level3[214]),
   .I0(level4_in[1284]),
   .I1(level4_in[1285]),
   .I2(level4_in[1286]),
   .I3(level4_in[1287]),
   .I4(level4_in[1288]),
   .I5(level4_in[1289])
);

LUT6 #(
   .INIT(64'h445147a8445147a8)  
) LUT6_inst7991 (
   .O(to_level3[215]),
   .I0(level4_in[1290]),
   .I1(level4_in[1291]),
   .I2(level4_in[1292]),
   .I3(level4_in[1293]),
   .I4(level4_in[1294]),
   .I5(level4_in[1295])
);

LUT6 #(
   .INIT(64'hd2973f3ad2973f3a)  
) LUT6_inst7992 (
   .O(to_level3[216]),
   .I0(level4_in[1296]),
   .I1(level4_in[1297]),
   .I2(level4_in[1298]),
   .I3(level4_in[1299]),
   .I4(level4_in[1300]),
   .I5(level4_in[1301])
);

LUT6 #(
   .INIT(64'h35824bd735824bd7)  
) LUT6_inst7993 (
   .O(to_level3[217]),
   .I0(level4_in[1302]),
   .I1(level4_in[1303]),
   .I2(level4_in[1304]),
   .I3(level4_in[1305]),
   .I4(level4_in[1306]),
   .I5(level4_in[1307])
);

LUT6 #(
   .INIT(64'h85895e4585895e45)  
) LUT6_inst7994 (
   .O(to_level3[218]),
   .I0(level4_in[1308]),
   .I1(level4_in[1309]),
   .I2(level4_in[1310]),
   .I3(level4_in[1311]),
   .I4(level4_in[1312]),
   .I5(level4_in[1313])
);

LUT6 #(
   .INIT(64'h60cf116e60cf116e)  
) LUT6_inst7995 (
   .O(to_level3[219]),
   .I0(level4_in[1314]),
   .I1(level4_in[1315]),
   .I2(level4_in[1316]),
   .I3(level4_in[1317]),
   .I4(level4_in[1318]),
   .I5(level4_in[1319])
);

LUT6 #(
   .INIT(64'h7e23c5e47e23c5e4)  
) LUT6_inst7996 (
   .O(to_level3[220]),
   .I0(level4_in[1320]),
   .I1(level4_in[1321]),
   .I2(level4_in[1322]),
   .I3(level4_in[1323]),
   .I4(level4_in[1324]),
   .I5(level4_in[1325])
);

LUT6 #(
   .INIT(64'ha174280ea174280e)  
) LUT6_inst7997 (
   .O(to_level3[221]),
   .I0(level4_in[1326]),
   .I1(level4_in[1327]),
   .I2(level4_in[1328]),
   .I3(level4_in[1329]),
   .I4(level4_in[1330]),
   .I5(level4_in[1331])
);

LUT6 #(
   .INIT(64'hfe253997fe253997)  
) LUT6_inst7998 (
   .O(to_level3[222]),
   .I0(level4_in[1332]),
   .I1(level4_in[1333]),
   .I2(level4_in[1334]),
   .I3(level4_in[1335]),
   .I4(level4_in[1336]),
   .I5(level4_in[1337])
);

LUT6 #(
   .INIT(64'h3332665933326659)  
) LUT6_inst7999 (
   .O(to_level3[223]),
   .I0(level4_in[1338]),
   .I1(level4_in[1339]),
   .I2(level4_in[1340]),
   .I3(level4_in[1341]),
   .I4(level4_in[1342]),
   .I5(level4_in[1343])
);

LUT6 #(
   .INIT(64'hf109d2b4f109d2b4)  
) LUT6_inst8000 (
   .O(to_level3[224]),
   .I0(level4_in[1344]),
   .I1(level4_in[1345]),
   .I2(level4_in[1346]),
   .I3(level4_in[1347]),
   .I4(level4_in[1348]),
   .I5(level4_in[1349])
);

LUT6 #(
   .INIT(64'h583575ad583575ad)  
) LUT6_inst8001 (
   .O(to_level3[225]),
   .I0(level4_in[1350]),
   .I1(level4_in[1351]),
   .I2(level4_in[1352]),
   .I3(level4_in[1353]),
   .I4(level4_in[1354]),
   .I5(level4_in[1355])
);

LUT6 #(
   .INIT(64'h6639aab36639aab3)  
) LUT6_inst8002 (
   .O(to_level3[226]),
   .I0(level4_in[1356]),
   .I1(level4_in[1357]),
   .I2(level4_in[1358]),
   .I3(level4_in[1359]),
   .I4(level4_in[1360]),
   .I5(level4_in[1361])
);

LUT6 #(
   .INIT(64'h26008ecb26008ecb)  
) LUT6_inst8003 (
   .O(to_level3[227]),
   .I0(level4_in[1362]),
   .I1(level4_in[1363]),
   .I2(level4_in[1364]),
   .I3(level4_in[1365]),
   .I4(level4_in[1366]),
   .I5(level4_in[1367])
);

LUT6 #(
   .INIT(64'h303b26f4303b26f4)  
) LUT6_inst8004 (
   .O(to_level3[228]),
   .I0(level4_in[1368]),
   .I1(level4_in[1369]),
   .I2(level4_in[1370]),
   .I3(level4_in[1371]),
   .I4(level4_in[1372]),
   .I5(level4_in[1373])
);

LUT6 #(
   .INIT(64'heff7cf26eff7cf26)  
) LUT6_inst8005 (
   .O(to_level3[229]),
   .I0(level4_in[1374]),
   .I1(level4_in[1375]),
   .I2(level4_in[1376]),
   .I3(level4_in[1377]),
   .I4(level4_in[1378]),
   .I5(level4_in[1379])
);

LUT6 #(
   .INIT(64'h68ed2b3d68ed2b3d)  
) LUT6_inst8006 (
   .O(to_level3[230]),
   .I0(level4_in[1380]),
   .I1(level4_in[1381]),
   .I2(level4_in[1382]),
   .I3(level4_in[1383]),
   .I4(level4_in[1384]),
   .I5(level4_in[1385])
);

LUT6 #(
   .INIT(64'hfceb4609fceb4609)  
) LUT6_inst8007 (
   .O(to_level3[231]),
   .I0(level4_in[1386]),
   .I1(level4_in[1387]),
   .I2(level4_in[1388]),
   .I3(level4_in[1389]),
   .I4(level4_in[1390]),
   .I5(level4_in[1391])
);

LUT6 #(
   .INIT(64'h4b3a10a14b3a10a1)  
) LUT6_inst8008 (
   .O(to_level3[232]),
   .I0(level4_in[1392]),
   .I1(level4_in[1393]),
   .I2(level4_in[1394]),
   .I3(level4_in[1395]),
   .I4(level4_in[1396]),
   .I5(level4_in[1397])
);

LUT6 #(
   .INIT(64'h17fd4eb317fd4eb3)  
) LUT6_inst8009 (
   .O(to_level3[233]),
   .I0(level4_in[1398]),
   .I1(level4_in[1399]),
   .I2(level4_in[1400]),
   .I3(level4_in[1401]),
   .I4(level4_in[1402]),
   .I5(level4_in[1403])
);

LUT6 #(
   .INIT(64'h95c8f3dc95c8f3dc)  
) LUT6_inst8010 (
   .O(to_level3[234]),
   .I0(level4_in[1404]),
   .I1(level4_in[1405]),
   .I2(level4_in[1406]),
   .I3(level4_in[1407]),
   .I4(level4_in[1408]),
   .I5(level4_in[1409])
);

LUT6 #(
   .INIT(64'h71f1375f71f1375f)  
) LUT6_inst8011 (
   .O(to_level3[235]),
   .I0(level4_in[1410]),
   .I1(level4_in[1411]),
   .I2(level4_in[1412]),
   .I3(level4_in[1413]),
   .I4(level4_in[1414]),
   .I5(level4_in[1415])
);

LUT6 #(
   .INIT(64'h89c0c4ec89c0c4ec)  
) LUT6_inst8012 (
   .O(to_level3[236]),
   .I0(level4_in[1416]),
   .I1(level4_in[1417]),
   .I2(level4_in[1418]),
   .I3(level4_in[1419]),
   .I4(level4_in[1420]),
   .I5(level4_in[1421])
);

LUT6 #(
   .INIT(64'hd512cf70d512cf70)  
) LUT6_inst8013 (
   .O(to_level3[237]),
   .I0(level4_in[1422]),
   .I1(level4_in[1423]),
   .I2(level4_in[1424]),
   .I3(level4_in[1425]),
   .I4(level4_in[1426]),
   .I5(level4_in[1427])
);

LUT6 #(
   .INIT(64'hdc0b0dfcdc0b0dfc)  
) LUT6_inst8014 (
   .O(to_level3[238]),
   .I0(level4_in[1428]),
   .I1(level4_in[1429]),
   .I2(level4_in[1430]),
   .I3(level4_in[1431]),
   .I4(level4_in[1432]),
   .I5(level4_in[1433])
);

LUT6 #(
   .INIT(64'hb9ae6dcbb9ae6dcb)  
) LUT6_inst8015 (
   .O(to_level3[239]),
   .I0(level4_in[1434]),
   .I1(level4_in[1435]),
   .I2(level4_in[1436]),
   .I3(level4_in[1437]),
   .I4(level4_in[1438]),
   .I5(level4_in[1439])
);

LUT6 #(
   .INIT(64'h4b37c1bd4b37c1bd)  
) LUT6_inst8016 (
   .O(to_level3[240]),
   .I0(level4_in[1440]),
   .I1(level4_in[1441]),
   .I2(level4_in[1442]),
   .I3(level4_in[1443]),
   .I4(level4_in[1444]),
   .I5(level4_in[1445])
);

LUT6 #(
   .INIT(64'h4c90ed7f4c90ed7f)  
) LUT6_inst8017 (
   .O(to_level3[241]),
   .I0(level4_in[1446]),
   .I1(level4_in[1447]),
   .I2(level4_in[1448]),
   .I3(level4_in[1449]),
   .I4(level4_in[1450]),
   .I5(level4_in[1451])
);

LUT6 #(
   .INIT(64'h3ef4d20e3ef4d20e)  
) LUT6_inst8018 (
   .O(to_level3[242]),
   .I0(level4_in[1452]),
   .I1(level4_in[1453]),
   .I2(level4_in[1454]),
   .I3(level4_in[1455]),
   .I4(level4_in[1456]),
   .I5(level4_in[1457])
);

LUT6 #(
   .INIT(64'hc009c440c009c440)  
) LUT6_inst8019 (
   .O(to_level3[243]),
   .I0(level4_in[1458]),
   .I1(level4_in[1459]),
   .I2(level4_in[1460]),
   .I3(level4_in[1461]),
   .I4(level4_in[1462]),
   .I5(level4_in[1463])
);

LUT6 #(
   .INIT(64'h2921abdc2921abdc)  
) LUT6_inst8020 (
   .O(to_level3[244]),
   .I0(level4_in[1464]),
   .I1(level4_in[1465]),
   .I2(level4_in[1466]),
   .I3(level4_in[1467]),
   .I4(level4_in[1468]),
   .I5(level4_in[1469])
);

LUT6 #(
   .INIT(64'h830ca3b4830ca3b4)  
) LUT6_inst8021 (
   .O(to_level3[245]),
   .I0(level4_in[1470]),
   .I1(level4_in[1471]),
   .I2(level4_in[1472]),
   .I3(level4_in[1473]),
   .I4(level4_in[1474]),
   .I5(level4_in[1475])
);

LUT6 #(
   .INIT(64'hca9fac56ca9fac56)  
) LUT6_inst8022 (
   .O(to_level3[246]),
   .I0(level4_in[1476]),
   .I1(level4_in[1477]),
   .I2(level4_in[1478]),
   .I3(level4_in[1479]),
   .I4(level4_in[1480]),
   .I5(level4_in[1481])
);

LUT6 #(
   .INIT(64'h0a57d9e80a57d9e8)  
) LUT6_inst8023 (
   .O(to_level3[247]),
   .I0(level4_in[1482]),
   .I1(level4_in[1483]),
   .I2(level4_in[1484]),
   .I3(level4_in[1485]),
   .I4(level4_in[1486]),
   .I5(level4_in[1487])
);

LUT6 #(
   .INIT(64'he491431ae491431a)  
) LUT6_inst8024 (
   .O(to_level3[248]),
   .I0(level4_in[1488]),
   .I1(level4_in[1489]),
   .I2(level4_in[1490]),
   .I3(level4_in[1491]),
   .I4(level4_in[1492]),
   .I5(level4_in[1493])
);

LUT6 #(
   .INIT(64'h1b8ae00c1b8ae00c)  
) LUT6_inst8025 (
   .O(to_level3[249]),
   .I0(level4_in[1494]),
   .I1(level4_in[1495]),
   .I2(level4_in[1496]),
   .I3(level4_in[1497]),
   .I4(level4_in[1498]),
   .I5(level4_in[1499])
);

LUT6 #(
   .INIT(64'hd503462fd503462f)  
) LUT6_inst8026 (
   .O(to_level3[250]),
   .I0(level4_in[1500]),
   .I1(level4_in[1501]),
   .I2(level4_in[1502]),
   .I3(level4_in[1503]),
   .I4(level4_in[1504]),
   .I5(level4_in[1505])
);

LUT6 #(
   .INIT(64'he647a95ee647a95e)  
) LUT6_inst8027 (
   .O(to_level3[251]),
   .I0(level4_in[1506]),
   .I1(level4_in[1507]),
   .I2(level4_in[1508]),
   .I3(level4_in[1509]),
   .I4(level4_in[1510]),
   .I5(level4_in[1511])
);

LUT6 #(
   .INIT(64'h55257d3b55257d3b)  
) LUT6_inst8028 (
   .O(to_level3[252]),
   .I0(level4_in[1512]),
   .I1(level4_in[1513]),
   .I2(level4_in[1514]),
   .I3(level4_in[1515]),
   .I4(level4_in[1516]),
   .I5(level4_in[1517])
);

LUT6 #(
   .INIT(64'h6f7730346f773034)  
) LUT6_inst8029 (
   .O(to_level3[253]),
   .I0(level4_in[1518]),
   .I1(level4_in[1519]),
   .I2(level4_in[1520]),
   .I3(level4_in[1521]),
   .I4(level4_in[1522]),
   .I5(level4_in[1523])
);

LUT6 #(
   .INIT(64'hdc043c95dc043c95)  
) LUT6_inst8030 (
   .O(to_level3[254]),
   .I0(level4_in[1524]),
   .I1(level4_in[1525]),
   .I2(level4_in[1526]),
   .I3(level4_in[1527]),
   .I4(level4_in[1528]),
   .I5(level4_in[1529])
);

LUT6 #(
   .INIT(64'h1917206419172064)  
) LUT6_inst8031 (
   .O(to_level3[255]),
   .I0(level4_in[1530]),
   .I1(level4_in[1531]),
   .I2(level4_in[1532]),
   .I3(level4_in[1533]),
   .I4(level4_in[1534]),
   .I5(level4_in[1535])
);

LUT6 #(
   .INIT(64'h8e867da78e867da7)  
) LUT6_inst8032 (
   .O(to_level3[256]),
   .I0(level4_in[1536]),
   .I1(level4_in[1537]),
   .I2(level4_in[1538]),
   .I3(level4_in[1539]),
   .I4(level4_in[1540]),
   .I5(level4_in[1541])
);

LUT6 #(
   .INIT(64'h40bfa1f040bfa1f0)  
) LUT6_inst8033 (
   .O(to_level3[257]),
   .I0(level4_in[1542]),
   .I1(level4_in[1543]),
   .I2(level4_in[1544]),
   .I3(level4_in[1545]),
   .I4(level4_in[1546]),
   .I5(level4_in[1547])
);

LUT6 #(
   .INIT(64'h8692b9ac8692b9ac)  
) LUT6_inst8034 (
   .O(to_level3[258]),
   .I0(level4_in[1548]),
   .I1(level4_in[1549]),
   .I2(level4_in[1550]),
   .I3(level4_in[1551]),
   .I4(level4_in[1552]),
   .I5(level4_in[1553])
);

LUT6 #(
   .INIT(64'h5140ada05140ada0)  
) LUT6_inst8035 (
   .O(to_level3[259]),
   .I0(level4_in[1554]),
   .I1(level4_in[1555]),
   .I2(level4_in[1556]),
   .I3(level4_in[1557]),
   .I4(level4_in[1558]),
   .I5(level4_in[1559])
);

LUT6 #(
   .INIT(64'hcb2b46facb2b46fa)  
) LUT6_inst8036 (
   .O(to_level3[260]),
   .I0(level4_in[1560]),
   .I1(level4_in[1561]),
   .I2(level4_in[1562]),
   .I3(level4_in[1563]),
   .I4(level4_in[1564]),
   .I5(level4_in[1565])
);

LUT6 #(
   .INIT(64'h987af1d9987af1d9)  
) LUT6_inst8037 (
   .O(to_level3[261]),
   .I0(level4_in[1566]),
   .I1(level4_in[1567]),
   .I2(level4_in[1568]),
   .I3(level4_in[1569]),
   .I4(level4_in[1570]),
   .I5(level4_in[1571])
);

LUT6 #(
   .INIT(64'h814a8a4a814a8a4a)  
) LUT6_inst8038 (
   .O(to_level3[262]),
   .I0(level4_in[1572]),
   .I1(level4_in[1573]),
   .I2(level4_in[1574]),
   .I3(level4_in[1575]),
   .I4(level4_in[1576]),
   .I5(level4_in[1577])
);

LUT6 #(
   .INIT(64'h96c95ebb96c95ebb)  
) LUT6_inst8039 (
   .O(to_level3[263]),
   .I0(level4_in[1578]),
   .I1(level4_in[1579]),
   .I2(level4_in[1580]),
   .I3(level4_in[1581]),
   .I4(level4_in[1582]),
   .I5(level4_in[1583])
);

LUT6 #(
   .INIT(64'h4e98ac954e98ac95)  
) LUT6_inst8040 (
   .O(to_level3[264]),
   .I0(level4_in[1584]),
   .I1(level4_in[1585]),
   .I2(level4_in[1586]),
   .I3(level4_in[1587]),
   .I4(level4_in[1588]),
   .I5(level4_in[1589])
);

LUT6 #(
   .INIT(64'h3c8caf593c8caf59)  
) LUT6_inst8041 (
   .O(to_level3[265]),
   .I0(level4_in[1590]),
   .I1(level4_in[1591]),
   .I2(level4_in[1592]),
   .I3(level4_in[1593]),
   .I4(level4_in[1594]),
   .I5(level4_in[1595])
);

LUT6 #(
   .INIT(64'hd5f62b5cd5f62b5c)  
) LUT6_inst8042 (
   .O(to_level3[266]),
   .I0(level4_in[1596]),
   .I1(level4_in[1597]),
   .I2(level4_in[1598]),
   .I3(level4_in[1599]),
   .I4(level4_in[1600]),
   .I5(level4_in[1601])
);

LUT6 #(
   .INIT(64'he703f3f4e703f3f4)  
) LUT6_inst8043 (
   .O(to_level3[267]),
   .I0(level4_in[1602]),
   .I1(level4_in[1603]),
   .I2(level4_in[1604]),
   .I3(level4_in[1605]),
   .I4(level4_in[1606]),
   .I5(level4_in[1607])
);

LUT6 #(
   .INIT(64'h92fcc7bf92fcc7bf)  
) LUT6_inst8044 (
   .O(to_level3[268]),
   .I0(level4_in[1608]),
   .I1(level4_in[1609]),
   .I2(level4_in[1610]),
   .I3(level4_in[1611]),
   .I4(level4_in[1612]),
   .I5(level4_in[1613])
);

LUT6 #(
   .INIT(64'h77d6cad277d6cad2)  
) LUT6_inst8045 (
   .O(to_level3[269]),
   .I0(level4_in[1614]),
   .I1(level4_in[1615]),
   .I2(level4_in[1616]),
   .I3(level4_in[1617]),
   .I4(level4_in[1618]),
   .I5(level4_in[1619])
);

LUT6 #(
   .INIT(64'h81ecba9081ecba90)  
) LUT6_inst8046 (
   .O(to_level3[270]),
   .I0(level4_in[1620]),
   .I1(level4_in[1621]),
   .I2(level4_in[1622]),
   .I3(level4_in[1623]),
   .I4(level4_in[1624]),
   .I5(level4_in[1625])
);

LUT6 #(
   .INIT(64'h9cbffbbe9cbffbbe)  
) LUT6_inst8047 (
   .O(to_level3[271]),
   .I0(level4_in[1626]),
   .I1(level4_in[1627]),
   .I2(level4_in[1628]),
   .I3(level4_in[1629]),
   .I4(level4_in[1630]),
   .I5(level4_in[1631])
);

LUT6 #(
   .INIT(64'h7bd2b9a27bd2b9a2)  
) LUT6_inst8048 (
   .O(to_level3[272]),
   .I0(level4_in[1632]),
   .I1(level4_in[1633]),
   .I2(level4_in[1634]),
   .I3(level4_in[1635]),
   .I4(level4_in[1636]),
   .I5(level4_in[1637])
);

LUT6 #(
   .INIT(64'hace511baace511ba)  
) LUT6_inst8049 (
   .O(to_level3[273]),
   .I0(level4_in[1638]),
   .I1(level4_in[1639]),
   .I2(level4_in[1640]),
   .I3(level4_in[1641]),
   .I4(level4_in[1642]),
   .I5(level4_in[1643])
);

LUT6 #(
   .INIT(64'heedd15aceedd15ac)  
) LUT6_inst8050 (
   .O(to_level3[274]),
   .I0(level4_in[1644]),
   .I1(level4_in[1645]),
   .I2(level4_in[1646]),
   .I3(level4_in[1647]),
   .I4(level4_in[1648]),
   .I5(level4_in[1649])
);

LUT6 #(
   .INIT(64'h0417756104177561)  
) LUT6_inst8051 (
   .O(to_level3[275]),
   .I0(level4_in[1650]),
   .I1(level4_in[1651]),
   .I2(level4_in[1652]),
   .I3(level4_in[1653]),
   .I4(level4_in[1654]),
   .I5(level4_in[1655])
);

LUT6 #(
   .INIT(64'h97050b6c97050b6c)  
) LUT6_inst8052 (
   .O(to_level3[276]),
   .I0(level4_in[1656]),
   .I1(level4_in[1657]),
   .I2(level4_in[1658]),
   .I3(level4_in[1659]),
   .I4(level4_in[1660]),
   .I5(level4_in[1661])
);

LUT6 #(
   .INIT(64'h3993151a3993151a)  
) LUT6_inst8053 (
   .O(to_level3[277]),
   .I0(level4_in[1662]),
   .I1(level4_in[1663]),
   .I2(level4_in[1664]),
   .I3(level4_in[1665]),
   .I4(level4_in[1666]),
   .I5(level4_in[1667])
);

LUT6 #(
   .INIT(64'h4ddaaa184ddaaa18)  
) LUT6_inst8054 (
   .O(to_level3[278]),
   .I0(level4_in[1668]),
   .I1(level4_in[1669]),
   .I2(level4_in[1670]),
   .I3(level4_in[1671]),
   .I4(level4_in[1672]),
   .I5(level4_in[1673])
);

LUT6 #(
   .INIT(64'hcaa422f8caa422f8)  
) LUT6_inst8055 (
   .O(to_level3[279]),
   .I0(level4_in[1674]),
   .I1(level4_in[1675]),
   .I2(level4_in[1676]),
   .I3(level4_in[1677]),
   .I4(level4_in[1678]),
   .I5(level4_in[1679])
);

LUT6 #(
   .INIT(64'h0ae902110ae90211)  
) LUT6_inst8056 (
   .O(to_level3[280]),
   .I0(level4_in[1680]),
   .I1(level4_in[1681]),
   .I2(level4_in[1682]),
   .I3(level4_in[1683]),
   .I4(level4_in[1684]),
   .I5(level4_in[1685])
);

LUT6 #(
   .INIT(64'hc337c721c337c721)  
) LUT6_inst8057 (
   .O(to_level3[281]),
   .I0(level4_in[1686]),
   .I1(level4_in[1687]),
   .I2(level4_in[1688]),
   .I3(level4_in[1689]),
   .I4(level4_in[1690]),
   .I5(level4_in[1691])
);

LUT6 #(
   .INIT(64'h466c8862466c8862)  
) LUT6_inst8058 (
   .O(to_level3[282]),
   .I0(level4_in[1692]),
   .I1(level4_in[1693]),
   .I2(level4_in[1694]),
   .I3(level4_in[1695]),
   .I4(level4_in[1696]),
   .I5(level4_in[1697])
);

LUT6 #(
   .INIT(64'h9e7a64a69e7a64a6)  
) LUT6_inst8059 (
   .O(to_level3[283]),
   .I0(level4_in[1698]),
   .I1(level4_in[1699]),
   .I2(level4_in[1700]),
   .I3(level4_in[1701]),
   .I4(level4_in[1702]),
   .I5(level4_in[1703])
);

LUT6 #(
   .INIT(64'hf120a598f120a598)  
) LUT6_inst8060 (
   .O(to_level3[284]),
   .I0(level4_in[1704]),
   .I1(level4_in[1705]),
   .I2(level4_in[1706]),
   .I3(level4_in[1707]),
   .I4(level4_in[1708]),
   .I5(level4_in[1709])
);

LUT6 #(
   .INIT(64'h3772d8d13772d8d1)  
) LUT6_inst8061 (
   .O(to_level3[285]),
   .I0(level4_in[1710]),
   .I1(level4_in[1711]),
   .I2(level4_in[1712]),
   .I3(level4_in[1713]),
   .I4(level4_in[1714]),
   .I5(level4_in[1715])
);

LUT6 #(
   .INIT(64'h9c8d7eed9c8d7eed)  
) LUT6_inst8062 (
   .O(to_level3[286]),
   .I0(level4_in[1716]),
   .I1(level4_in[1717]),
   .I2(level4_in[1718]),
   .I3(level4_in[1719]),
   .I4(level4_in[1720]),
   .I5(level4_in[1721])
);

LUT6 #(
   .INIT(64'h4ada5b5e4ada5b5e)  
) LUT6_inst8063 (
   .O(to_level3[287]),
   .I0(level4_in[1722]),
   .I1(level4_in[1723]),
   .I2(level4_in[1724]),
   .I3(level4_in[1725]),
   .I4(level4_in[1726]),
   .I5(level4_in[1727])
);

LUT6 #(
   .INIT(64'h83d77dae83d77dae)  
) LUT6_inst8064 (
   .O(to_level3[288]),
   .I0(level4_in[1728]),
   .I1(level4_in[1729]),
   .I2(level4_in[1730]),
   .I3(level4_in[1731]),
   .I4(level4_in[1732]),
   .I5(level4_in[1733])
);

LUT6 #(
   .INIT(64'h6c75b9226c75b922)  
) LUT6_inst8065 (
   .O(to_level3[289]),
   .I0(level4_in[1734]),
   .I1(level4_in[1735]),
   .I2(level4_in[1736]),
   .I3(level4_in[1737]),
   .I4(level4_in[1738]),
   .I5(level4_in[1739])
);

LUT6 #(
   .INIT(64'h1961ecfd1961ecfd)  
) LUT6_inst8066 (
   .O(to_level3[290]),
   .I0(level4_in[1740]),
   .I1(level4_in[1741]),
   .I2(level4_in[1742]),
   .I3(level4_in[1743]),
   .I4(level4_in[1744]),
   .I5(level4_in[1745])
);

LUT6 #(
   .INIT(64'hf2a1aafaf2a1aafa)  
) LUT6_inst8067 (
   .O(to_level3[291]),
   .I0(level4_in[1746]),
   .I1(level4_in[1747]),
   .I2(level4_in[1748]),
   .I3(level4_in[1749]),
   .I4(level4_in[1750]),
   .I5(level4_in[1751])
);

LUT6 #(
   .INIT(64'h5f9ab0245f9ab024)  
) LUT6_inst8068 (
   .O(to_level3[292]),
   .I0(level4_in[1752]),
   .I1(level4_in[1753]),
   .I2(level4_in[1754]),
   .I3(level4_in[1755]),
   .I4(level4_in[1756]),
   .I5(level4_in[1757])
);

LUT6 #(
   .INIT(64'h8f9b7df08f9b7df0)  
) LUT6_inst8069 (
   .O(to_level3[293]),
   .I0(level4_in[1758]),
   .I1(level4_in[1759]),
   .I2(level4_in[1760]),
   .I3(level4_in[1761]),
   .I4(level4_in[1762]),
   .I5(level4_in[1763])
);

LUT6 #(
   .INIT(64'hcfe8e2bfcfe8e2bf)  
) LUT6_inst8070 (
   .O(to_level3[294]),
   .I0(level4_in[1764]),
   .I1(level4_in[1765]),
   .I2(level4_in[1766]),
   .I3(level4_in[1767]),
   .I4(level4_in[1768]),
   .I5(level4_in[1769])
);

LUT6 #(
   .INIT(64'hce1ba249ce1ba249)  
) LUT6_inst8071 (
   .O(to_level3[295]),
   .I0(level4_in[1770]),
   .I1(level4_in[1771]),
   .I2(level4_in[1772]),
   .I3(level4_in[1773]),
   .I4(level4_in[1774]),
   .I5(level4_in[1775])
);

LUT6 #(
   .INIT(64'hea4058adea4058ad)  
) LUT6_inst8072 (
   .O(to_level3[296]),
   .I0(level4_in[1776]),
   .I1(level4_in[1777]),
   .I2(level4_in[1778]),
   .I3(level4_in[1779]),
   .I4(level4_in[1780]),
   .I5(level4_in[1781])
);

LUT6 #(
   .INIT(64'hc9edb6ebc9edb6eb)  
) LUT6_inst8073 (
   .O(to_level3[297]),
   .I0(level4_in[1782]),
   .I1(level4_in[1783]),
   .I2(level4_in[1784]),
   .I3(level4_in[1785]),
   .I4(level4_in[1786]),
   .I5(level4_in[1787])
);

LUT6 #(
   .INIT(64'hda103242da103242)  
) LUT6_inst8074 (
   .O(to_level3[298]),
   .I0(level4_in[1788]),
   .I1(level4_in[1789]),
   .I2(level4_in[1790]),
   .I3(level4_in[1791]),
   .I4(level4_in[1792]),
   .I5(level4_in[1793])
);

LUT6 #(
   .INIT(64'h14cd68fc14cd68fc)  
) LUT6_inst8075 (
   .O(to_level3[299]),
   .I0(level4_in[1794]),
   .I1(level4_in[1795]),
   .I2(level4_in[1796]),
   .I3(level4_in[1797]),
   .I4(level4_in[1798]),
   .I5(level4_in[1799])
);

LUT6 #(
   .INIT(64'h054ceeb6054ceeb6)  
) LUT6_inst8076 (
   .O(to_level3[300]),
   .I0(level4_in[1800]),
   .I1(level4_in[1801]),
   .I2(level4_in[1802]),
   .I3(level4_in[1803]),
   .I4(level4_in[1804]),
   .I5(level4_in[1805])
);

LUT6 #(
   .INIT(64'ha9afd8b8a9afd8b8)  
) LUT6_inst8077 (
   .O(to_level3[301]),
   .I0(level4_in[1806]),
   .I1(level4_in[1807]),
   .I2(level4_in[1808]),
   .I3(level4_in[1809]),
   .I4(level4_in[1810]),
   .I5(level4_in[1811])
);

LUT6 #(
   .INIT(64'h9e844caa9e844caa)  
) LUT6_inst8078 (
   .O(to_level3[302]),
   .I0(level4_in[1812]),
   .I1(level4_in[1813]),
   .I2(level4_in[1814]),
   .I3(level4_in[1815]),
   .I4(level4_in[1816]),
   .I5(level4_in[1817])
);

LUT6 #(
   .INIT(64'h5fbaaebc5fbaaebc)  
) LUT6_inst8079 (
   .O(to_level3[303]),
   .I0(level4_in[1818]),
   .I1(level4_in[1819]),
   .I2(level4_in[1820]),
   .I3(level4_in[1821]),
   .I4(level4_in[1822]),
   .I5(level4_in[1823])
);

LUT6 #(
   .INIT(64'h885f9cca885f9cca)  
) LUT6_inst8080 (
   .O(to_level3[304]),
   .I0(level4_in[1824]),
   .I1(level4_in[1825]),
   .I2(level4_in[1826]),
   .I3(level4_in[1827]),
   .I4(level4_in[1828]),
   .I5(level4_in[1829])
);

LUT6 #(
   .INIT(64'hb693e6e1b693e6e1)  
) LUT6_inst8081 (
   .O(to_level3[305]),
   .I0(level4_in[1830]),
   .I1(level4_in[1831]),
   .I2(level4_in[1832]),
   .I3(level4_in[1833]),
   .I4(level4_in[1834]),
   .I5(level4_in[1835])
);

LUT6 #(
   .INIT(64'ha72802b0a72802b0)  
) LUT6_inst8082 (
   .O(to_level3[306]),
   .I0(level4_in[1836]),
   .I1(level4_in[1837]),
   .I2(level4_in[1838]),
   .I3(level4_in[1839]),
   .I4(level4_in[1840]),
   .I5(level4_in[1841])
);

LUT6 #(
   .INIT(64'h435399e4435399e4)  
) LUT6_inst8083 (
   .O(to_level3[307]),
   .I0(level4_in[1842]),
   .I1(level4_in[1843]),
   .I2(level4_in[1844]),
   .I3(level4_in[1845]),
   .I4(level4_in[1846]),
   .I5(level4_in[1847])
);

LUT6 #(
   .INIT(64'ha2954b3ea2954b3e)  
) LUT6_inst8084 (
   .O(to_level3[308]),
   .I0(level4_in[1848]),
   .I1(level4_in[1849]),
   .I2(level4_in[1850]),
   .I3(level4_in[1851]),
   .I4(level4_in[1852]),
   .I5(level4_in[1853])
);

LUT6 #(
   .INIT(64'ha3c675f2a3c675f2)  
) LUT6_inst8085 (
   .O(to_level3[309]),
   .I0(level4_in[1854]),
   .I1(level4_in[1855]),
   .I2(level4_in[1856]),
   .I3(level4_in[1857]),
   .I4(level4_in[1858]),
   .I5(level4_in[1859])
);

LUT6 #(
   .INIT(64'h8951374f8951374f)  
) LUT6_inst8086 (
   .O(to_level3[310]),
   .I0(level4_in[1860]),
   .I1(level4_in[1861]),
   .I2(level4_in[1862]),
   .I3(level4_in[1863]),
   .I4(level4_in[1864]),
   .I5(level4_in[1865])
);

LUT6 #(
   .INIT(64'hbd724c13bd724c13)  
) LUT6_inst8087 (
   .O(to_level3[311]),
   .I0(level4_in[1866]),
   .I1(level4_in[1867]),
   .I2(level4_in[1868]),
   .I3(level4_in[1869]),
   .I4(level4_in[1870]),
   .I5(level4_in[1871])
);

LUT6 #(
   .INIT(64'h7f9886497f988649)  
) LUT6_inst8088 (
   .O(to_level3[312]),
   .I0(level4_in[1872]),
   .I1(level4_in[1873]),
   .I2(level4_in[1874]),
   .I3(level4_in[1875]),
   .I4(level4_in[1876]),
   .I5(level4_in[1877])
);

LUT6 #(
   .INIT(64'h77d2e93f77d2e93f)  
) LUT6_inst8089 (
   .O(to_level3[313]),
   .I0(level4_in[1878]),
   .I1(level4_in[1879]),
   .I2(level4_in[1880]),
   .I3(level4_in[1881]),
   .I4(level4_in[1882]),
   .I5(level4_in[1883])
);

LUT6 #(
   .INIT(64'h13de3d1b13de3d1b)  
) LUT6_inst8090 (
   .O(to_level3[314]),
   .I0(level4_in[1884]),
   .I1(level4_in[1885]),
   .I2(level4_in[1886]),
   .I3(level4_in[1887]),
   .I4(level4_in[1888]),
   .I5(level4_in[1889])
);

LUT6 #(
   .INIT(64'h83516d7f83516d7f)  
) LUT6_inst8091 (
   .O(to_level3[315]),
   .I0(level4_in[1890]),
   .I1(level4_in[1891]),
   .I2(level4_in[1892]),
   .I3(level4_in[1893]),
   .I4(level4_in[1894]),
   .I5(level4_in[1895])
);

LUT6 #(
   .INIT(64'h6e4d78266e4d7826)  
) LUT6_inst8092 (
   .O(to_level3[316]),
   .I0(level4_in[1896]),
   .I1(level4_in[1897]),
   .I2(level4_in[1898]),
   .I3(level4_in[1899]),
   .I4(level4_in[1900]),
   .I5(level4_in[1901])
);

LUT6 #(
   .INIT(64'h15a038ff15a038ff)  
) LUT6_inst8093 (
   .O(to_level3[317]),
   .I0(level4_in[1902]),
   .I1(level4_in[1903]),
   .I2(level4_in[1904]),
   .I3(level4_in[1905]),
   .I4(level4_in[1906]),
   .I5(level4_in[1907])
);

LUT6 #(
   .INIT(64'h49ca09b849ca09b8)  
) LUT6_inst8094 (
   .O(to_level3[318]),
   .I0(level4_in[1908]),
   .I1(level4_in[1909]),
   .I2(level4_in[1910]),
   .I3(level4_in[1911]),
   .I4(level4_in[1912]),
   .I5(level4_in[1913])
);

LUT6 #(
   .INIT(64'he2a43150e2a43150)  
) LUT6_inst8095 (
   .O(to_level3[319]),
   .I0(level4_in[1914]),
   .I1(level4_in[1915]),
   .I2(level4_in[1916]),
   .I3(level4_in[1917]),
   .I4(level4_in[1918]),
   .I5(level4_in[1919])
);

LUT6 #(
   .INIT(64'h19160ce519160ce5)  
) LUT6_inst8096 (
   .O(to_level3[320]),
   .I0(level4_in[1920]),
   .I1(level4_in[1921]),
   .I2(level4_in[1922]),
   .I3(level4_in[1923]),
   .I4(level4_in[1924]),
   .I5(level4_in[1925])
);

LUT6 #(
   .INIT(64'hb691f66cb691f66c)  
) LUT6_inst8097 (
   .O(to_level3[321]),
   .I0(level4_in[1926]),
   .I1(level4_in[1927]),
   .I2(level4_in[1928]),
   .I3(level4_in[1929]),
   .I4(level4_in[1930]),
   .I5(level4_in[1931])
);

LUT6 #(
   .INIT(64'h3adf5dc23adf5dc2)  
) LUT6_inst8098 (
   .O(to_level3[322]),
   .I0(level4_in[1932]),
   .I1(level4_in[1933]),
   .I2(level4_in[1934]),
   .I3(level4_in[1935]),
   .I4(level4_in[1936]),
   .I5(level4_in[1937])
);

LUT6 #(
   .INIT(64'h216eafc4216eafc4)  
) LUT6_inst8099 (
   .O(to_level3[323]),
   .I0(level4_in[1938]),
   .I1(level4_in[1939]),
   .I2(level4_in[1940]),
   .I3(level4_in[1941]),
   .I4(level4_in[1942]),
   .I5(level4_in[1943])
);

LUT6 #(
   .INIT(64'h14c2908c14c2908c)  
) LUT6_inst8100 (
   .O(to_level3[324]),
   .I0(level4_in[1944]),
   .I1(level4_in[1945]),
   .I2(level4_in[1946]),
   .I3(level4_in[1947]),
   .I4(level4_in[1948]),
   .I5(level4_in[1949])
);

LUT6 #(
   .INIT(64'hde667b97de667b97)  
) LUT6_inst8101 (
   .O(to_level3[325]),
   .I0(level4_in[1950]),
   .I1(level4_in[1951]),
   .I2(level4_in[1952]),
   .I3(level4_in[1953]),
   .I4(level4_in[1954]),
   .I5(level4_in[1955])
);

LUT6 #(
   .INIT(64'h3dd07ea73dd07ea7)  
) LUT6_inst8102 (
   .O(to_level3[326]),
   .I0(level4_in[1956]),
   .I1(level4_in[1957]),
   .I2(level4_in[1958]),
   .I3(level4_in[1959]),
   .I4(level4_in[1960]),
   .I5(level4_in[1961])
);

LUT6 #(
   .INIT(64'haf0c6ceeaf0c6cee)  
) LUT6_inst8103 (
   .O(to_level3[327]),
   .I0(level4_in[1962]),
   .I1(level4_in[1963]),
   .I2(level4_in[1964]),
   .I3(level4_in[1965]),
   .I4(level4_in[1966]),
   .I5(level4_in[1967])
);

LUT6 #(
   .INIT(64'h5a7c6ef35a7c6ef3)  
) LUT6_inst8104 (
   .O(to_level3[328]),
   .I0(level4_in[1968]),
   .I1(level4_in[1969]),
   .I2(level4_in[1970]),
   .I3(level4_in[1971]),
   .I4(level4_in[1972]),
   .I5(level4_in[1973])
);

LUT6 #(
   .INIT(64'hd74abd94d74abd94)  
) LUT6_inst8105 (
   .O(to_level3[329]),
   .I0(level4_in[1974]),
   .I1(level4_in[1975]),
   .I2(level4_in[1976]),
   .I3(level4_in[1977]),
   .I4(level4_in[1978]),
   .I5(level4_in[1979])
);

LUT6 #(
   .INIT(64'ha05051bba05051bb)  
) LUT6_inst8106 (
   .O(to_level3[330]),
   .I0(level4_in[1980]),
   .I1(level4_in[1981]),
   .I2(level4_in[1982]),
   .I3(level4_in[1983]),
   .I4(level4_in[1984]),
   .I5(level4_in[1985])
);

LUT6 #(
   .INIT(64'h1368b0941368b094)  
) LUT6_inst8107 (
   .O(to_level3[331]),
   .I0(level4_in[1986]),
   .I1(level4_in[1987]),
   .I2(level4_in[1988]),
   .I3(level4_in[1989]),
   .I4(level4_in[1990]),
   .I5(level4_in[1991])
);

LUT6 #(
   .INIT(64'hdddc46e9dddc46e9)  
) LUT6_inst8108 (
   .O(to_level3[332]),
   .I0(level4_in[1992]),
   .I1(level4_in[1993]),
   .I2(level4_in[1994]),
   .I3(level4_in[1995]),
   .I4(level4_in[1996]),
   .I5(level4_in[1997])
);

LUT6 #(
   .INIT(64'h85b8342c85b8342c)  
) LUT6_inst8109 (
   .O(to_level3[333]),
   .I0(level4_in[1998]),
   .I1(level4_in[1999]),
   .I2(level4_in[2000]),
   .I3(level4_in[2001]),
   .I4(level4_in[2002]),
   .I5(level4_in[2003])
);

LUT6 #(
   .INIT(64'h3d0dbb353d0dbb35)  
) LUT6_inst8110 (
   .O(to_level3[334]),
   .I0(level4_in[2004]),
   .I1(level4_in[2005]),
   .I2(level4_in[2006]),
   .I3(level4_in[2007]),
   .I4(level4_in[2008]),
   .I5(level4_in[2009])
);

LUT6 #(
   .INIT(64'h1ddb72b01ddb72b0)  
) LUT6_inst8111 (
   .O(to_level3[335]),
   .I0(level4_in[2010]),
   .I1(level4_in[2011]),
   .I2(level4_in[2012]),
   .I3(level4_in[2013]),
   .I4(level4_in[2014]),
   .I5(level4_in[2015])
);

LUT6 #(
   .INIT(64'hcad6932fcad6932f)  
) LUT6_inst8112 (
   .O(to_level3[336]),
   .I0(level4_in[2016]),
   .I1(level4_in[2017]),
   .I2(level4_in[2018]),
   .I3(level4_in[2019]),
   .I4(level4_in[2020]),
   .I5(level4_in[2021])
);

LUT6 #(
   .INIT(64'h94c3563c94c3563c)  
) LUT6_inst8113 (
   .O(to_level3[337]),
   .I0(level4_in[2022]),
   .I1(level4_in[2023]),
   .I2(level4_in[2024]),
   .I3(level4_in[2025]),
   .I4(level4_in[2026]),
   .I5(level4_in[2027])
);

LUT6 #(
   .INIT(64'h8220c2438220c243)  
) LUT6_inst8114 (
   .O(to_level3[338]),
   .I0(level4_in[2028]),
   .I1(level4_in[2029]),
   .I2(level4_in[2030]),
   .I3(level4_in[2031]),
   .I4(level4_in[2032]),
   .I5(level4_in[2033])
);

LUT6 #(
   .INIT(64'hb5074a13b5074a13)  
) LUT6_inst8115 (
   .O(to_level3[339]),
   .I0(level4_in[2034]),
   .I1(level4_in[2035]),
   .I2(level4_in[2036]),
   .I3(level4_in[2037]),
   .I4(level4_in[2038]),
   .I5(level4_in[2039])
);

LUT6 #(
   .INIT(64'h65db944c65db944c)  
) LUT6_inst8116 (
   .O(to_level3[340]),
   .I0(level4_in[2040]),
   .I1(level4_in[2041]),
   .I2(level4_in[2042]),
   .I3(level4_in[2043]),
   .I4(level4_in[2044]),
   .I5(level4_in[2045])
);

LUT6 #(
   .INIT(64'h19ceed7719ceed77)  
) LUT6_inst8117 (
   .O(to_level3[341]),
   .I0(level4_in[2046]),
   .I1(level4_in[2047]),
   .I2(level4_in[2048]),
   .I3(level4_in[2049]),
   .I4(level4_in[2050]),
   .I5(level4_in[2051])
);

LUT6 #(
   .INIT(64'h8a317cf68a317cf6)  
) LUT6_inst8118 (
   .O(to_level3[342]),
   .I0(level4_in[2052]),
   .I1(level4_in[2053]),
   .I2(level4_in[2054]),
   .I3(level4_in[2055]),
   .I4(level4_in[2056]),
   .I5(level4_in[2057])
);

LUT6 #(
   .INIT(64'hddfc7041ddfc7041)  
) LUT6_inst8119 (
   .O(to_level3[343]),
   .I0(level4_in[2058]),
   .I1(level4_in[2059]),
   .I2(level4_in[2060]),
   .I3(level4_in[2061]),
   .I4(level4_in[2062]),
   .I5(level4_in[2063])
);

LUT6 #(
   .INIT(64'h3cc8f8cc3cc8f8cc)  
) LUT6_inst8120 (
   .O(to_level3[344]),
   .I0(level4_in[2064]),
   .I1(level4_in[2065]),
   .I2(level4_in[2066]),
   .I3(level4_in[2067]),
   .I4(level4_in[2068]),
   .I5(level4_in[2069])
);

LUT6 #(
   .INIT(64'h3177707231777072)  
) LUT6_inst8121 (
   .O(to_level3[345]),
   .I0(level4_in[2070]),
   .I1(level4_in[2071]),
   .I2(level4_in[2072]),
   .I3(level4_in[2073]),
   .I4(level4_in[2074]),
   .I5(level4_in[2075])
);

LUT6 #(
   .INIT(64'h4463815244638152)  
) LUT6_inst8122 (
   .O(to_level3[346]),
   .I0(level4_in[2076]),
   .I1(level4_in[2077]),
   .I2(level4_in[2078]),
   .I3(level4_in[2079]),
   .I4(level4_in[2080]),
   .I5(level4_in[2081])
);

LUT6 #(
   .INIT(64'hee37cee3ee37cee3)  
) LUT6_inst8123 (
   .O(to_level3[347]),
   .I0(level4_in[2082]),
   .I1(level4_in[2083]),
   .I2(level4_in[2084]),
   .I3(level4_in[2085]),
   .I4(level4_in[2086]),
   .I5(level4_in[2087])
);

LUT6 #(
   .INIT(64'he4b62e0de4b62e0d)  
) LUT6_inst8124 (
   .O(to_level3[348]),
   .I0(level4_in[2088]),
   .I1(level4_in[2089]),
   .I2(level4_in[2090]),
   .I3(level4_in[2091]),
   .I4(level4_in[2092]),
   .I5(level4_in[2093])
);

LUT6 #(
   .INIT(64'h212a5ac8212a5ac8)  
) LUT6_inst8125 (
   .O(to_level3[349]),
   .I0(level4_in[2094]),
   .I1(level4_in[2095]),
   .I2(level4_in[2096]),
   .I3(level4_in[2097]),
   .I4(level4_in[2098]),
   .I5(level4_in[2099])
);

LUT6 #(
   .INIT(64'h0cf617110cf61711)  
) LUT6_inst8126 (
   .O(to_level3[350]),
   .I0(level4_in[2100]),
   .I1(level4_in[2101]),
   .I2(level4_in[2102]),
   .I3(level4_in[2103]),
   .I4(level4_in[2104]),
   .I5(level4_in[2105])
);

LUT6 #(
   .INIT(64'h1991dd741991dd74)  
) LUT6_inst8127 (
   .O(to_level3[351]),
   .I0(level4_in[2106]),
   .I1(level4_in[2107]),
   .I2(level4_in[2108]),
   .I3(level4_in[2109]),
   .I4(level4_in[2110]),
   .I5(level4_in[2111])
);

LUT6 #(
   .INIT(64'h3a5c45863a5c4586)  
) LUT6_inst8128 (
   .O(to_level3[352]),
   .I0(level4_in[2112]),
   .I1(level4_in[2113]),
   .I2(level4_in[2114]),
   .I3(level4_in[2115]),
   .I4(level4_in[2116]),
   .I5(level4_in[2117])
);

LUT6 #(
   .INIT(64'h795c63d8795c63d8)  
) LUT6_inst8129 (
   .O(to_level3[353]),
   .I0(level4_in[2118]),
   .I1(level4_in[2119]),
   .I2(level4_in[2120]),
   .I3(level4_in[2121]),
   .I4(level4_in[2122]),
   .I5(level4_in[2123])
);

LUT6 #(
   .INIT(64'h12d6263312d62633)  
) LUT6_inst8130 (
   .O(to_level3[354]),
   .I0(level4_in[2124]),
   .I1(level4_in[2125]),
   .I2(level4_in[2126]),
   .I3(level4_in[2127]),
   .I4(level4_in[2128]),
   .I5(level4_in[2129])
);

LUT6 #(
   .INIT(64'h0980d7480980d748)  
) LUT6_inst8131 (
   .O(to_level3[355]),
   .I0(level4_in[2130]),
   .I1(level4_in[2131]),
   .I2(level4_in[2132]),
   .I3(level4_in[2133]),
   .I4(level4_in[2134]),
   .I5(level4_in[2135])
);

LUT6 #(
   .INIT(64'h26bd1e5d26bd1e5d)  
) LUT6_inst8132 (
   .O(to_level3[356]),
   .I0(level4_in[2136]),
   .I1(level4_in[2137]),
   .I2(level4_in[2138]),
   .I3(level4_in[2139]),
   .I4(level4_in[2140]),
   .I5(level4_in[2141])
);

LUT6 #(
   .INIT(64'hae0217f8ae0217f8)  
) LUT6_inst8133 (
   .O(to_level3[357]),
   .I0(level4_in[2142]),
   .I1(level4_in[2143]),
   .I2(level4_in[2144]),
   .I3(level4_in[2145]),
   .I4(level4_in[2146]),
   .I5(level4_in[2147])
);

LUT6 #(
   .INIT(64'h034d373b034d373b)  
) LUT6_inst8134 (
   .O(to_level3[358]),
   .I0(level4_in[2148]),
   .I1(level4_in[2149]),
   .I2(level4_in[2150]),
   .I3(level4_in[2151]),
   .I4(level4_in[2152]),
   .I5(level4_in[2153])
);

LUT6 #(
   .INIT(64'h6195b6b46195b6b4)  
) LUT6_inst8135 (
   .O(to_level3[359]),
   .I0(level4_in[2154]),
   .I1(level4_in[2155]),
   .I2(level4_in[2156]),
   .I3(level4_in[2157]),
   .I4(level4_in[2158]),
   .I5(level4_in[2159])
);

LUT6 #(
   .INIT(64'hb737f8a1b737f8a1)  
) LUT6_inst8136 (
   .O(to_level3[360]),
   .I0(level4_in[2160]),
   .I1(level4_in[2161]),
   .I2(level4_in[2162]),
   .I3(level4_in[2163]),
   .I4(level4_in[2164]),
   .I5(level4_in[2165])
);

LUT6 #(
   .INIT(64'h9fbdaf6e9fbdaf6e)  
) LUT6_inst8137 (
   .O(to_level3[361]),
   .I0(level4_in[2166]),
   .I1(level4_in[2167]),
   .I2(level4_in[2168]),
   .I3(level4_in[2169]),
   .I4(level4_in[2170]),
   .I5(level4_in[2171])
);

LUT6 #(
   .INIT(64'h80c092df80c092df)  
) LUT6_inst8138 (
   .O(to_level3[362]),
   .I0(level4_in[2172]),
   .I1(level4_in[2173]),
   .I2(level4_in[2174]),
   .I3(level4_in[2175]),
   .I4(level4_in[2176]),
   .I5(level4_in[2177])
);

LUT6 #(
   .INIT(64'h0df0e5e30df0e5e3)  
) LUT6_inst8139 (
   .O(to_level3[363]),
   .I0(level4_in[2178]),
   .I1(level4_in[2179]),
   .I2(level4_in[2180]),
   .I3(level4_in[2181]),
   .I4(level4_in[2182]),
   .I5(level4_in[2183])
);

LUT6 #(
   .INIT(64'h44b6f68344b6f683)  
) LUT6_inst8140 (
   .O(to_level3[364]),
   .I0(level4_in[2184]),
   .I1(level4_in[2185]),
   .I2(level4_in[2186]),
   .I3(level4_in[2187]),
   .I4(level4_in[2188]),
   .I5(level4_in[2189])
);

LUT6 #(
   .INIT(64'h2529f7582529f758)  
) LUT6_inst8141 (
   .O(to_level3[365]),
   .I0(level4_in[2190]),
   .I1(level4_in[2191]),
   .I2(level4_in[2192]),
   .I3(level4_in[2193]),
   .I4(level4_in[2194]),
   .I5(level4_in[2195])
);

LUT6 #(
   .INIT(64'h6771227b6771227b)  
) LUT6_inst8142 (
   .O(to_level3[366]),
   .I0(level4_in[2196]),
   .I1(level4_in[2197]),
   .I2(level4_in[2198]),
   .I3(level4_in[2199]),
   .I4(level4_in[2200]),
   .I5(level4_in[2201])
);

LUT6 #(
   .INIT(64'hff3aa004ff3aa004)  
) LUT6_inst8143 (
   .O(to_level3[367]),
   .I0(level4_in[2202]),
   .I1(level4_in[2203]),
   .I2(level4_in[2204]),
   .I3(level4_in[2205]),
   .I4(level4_in[2206]),
   .I5(level4_in[2207])
);

LUT6 #(
   .INIT(64'h2c62d8fa2c62d8fa)  
) LUT6_inst8144 (
   .O(to_level3[368]),
   .I0(level4_in[2208]),
   .I1(level4_in[2209]),
   .I2(level4_in[2210]),
   .I3(level4_in[2211]),
   .I4(level4_in[2212]),
   .I5(level4_in[2213])
);

LUT6 #(
   .INIT(64'h6f908bc76f908bc7)  
) LUT6_inst8145 (
   .O(to_level3[369]),
   .I0(level4_in[2214]),
   .I1(level4_in[2215]),
   .I2(level4_in[2216]),
   .I3(level4_in[2217]),
   .I4(level4_in[2218]),
   .I5(level4_in[2219])
);

LUT6 #(
   .INIT(64'habde6f81abde6f81)  
) LUT6_inst8146 (
   .O(to_level3[370]),
   .I0(level4_in[2220]),
   .I1(level4_in[2221]),
   .I2(level4_in[2222]),
   .I3(level4_in[2223]),
   .I4(level4_in[2224]),
   .I5(level4_in[2225])
);

LUT6 #(
   .INIT(64'h562dc2fa562dc2fa)  
) LUT6_inst8147 (
   .O(to_level3[371]),
   .I0(level4_in[2226]),
   .I1(level4_in[2227]),
   .I2(level4_in[2228]),
   .I3(level4_in[2229]),
   .I4(level4_in[2230]),
   .I5(level4_in[2231])
);

LUT6 #(
   .INIT(64'hf901f2cff901f2cf)  
) LUT6_inst8148 (
   .O(to_level3[372]),
   .I0(level4_in[2232]),
   .I1(level4_in[2233]),
   .I2(level4_in[2234]),
   .I3(level4_in[2235]),
   .I4(level4_in[2236]),
   .I5(level4_in[2237])
);

LUT6 #(
   .INIT(64'ha59677a2a59677a2)  
) LUT6_inst8149 (
   .O(to_level3[373]),
   .I0(level4_in[2238]),
   .I1(level4_in[2239]),
   .I2(level4_in[2240]),
   .I3(level4_in[2241]),
   .I4(level4_in[2242]),
   .I5(level4_in[2243])
);

LUT6 #(
   .INIT(64'h78a2936578a29365)  
) LUT6_inst8150 (
   .O(to_level3[374]),
   .I0(level4_in[2244]),
   .I1(level4_in[2245]),
   .I2(level4_in[2246]),
   .I3(level4_in[2247]),
   .I4(level4_in[2248]),
   .I5(level4_in[2249])
);

LUT6 #(
   .INIT(64'h653bb9be653bb9be)  
) LUT6_inst8151 (
   .O(to_level3[375]),
   .I0(level4_in[2250]),
   .I1(level4_in[2251]),
   .I2(level4_in[2252]),
   .I3(level4_in[2253]),
   .I4(level4_in[2254]),
   .I5(level4_in[2255])
);

LUT6 #(
   .INIT(64'h7c9354a37c9354a3)  
) LUT6_inst8152 (
   .O(to_level3[376]),
   .I0(level4_in[2256]),
   .I1(level4_in[2257]),
   .I2(level4_in[2258]),
   .I3(level4_in[2259]),
   .I4(level4_in[2260]),
   .I5(level4_in[2261])
);

LUT6 #(
   .INIT(64'h2b4f97f12b4f97f1)  
) LUT6_inst8153 (
   .O(to_level3[377]),
   .I0(level4_in[2262]),
   .I1(level4_in[2263]),
   .I2(level4_in[2264]),
   .I3(level4_in[2265]),
   .I4(level4_in[2266]),
   .I5(level4_in[2267])
);

LUT6 #(
   .INIT(64'h05348b4105348b41)  
) LUT6_inst8154 (
   .O(to_level3[378]),
   .I0(level4_in[2268]),
   .I1(level4_in[2269]),
   .I2(level4_in[2270]),
   .I3(level4_in[2271]),
   .I4(level4_in[2272]),
   .I5(level4_in[2273])
);

LUT6 #(
   .INIT(64'hc916a12cc916a12c)  
) LUT6_inst8155 (
   .O(to_level3[379]),
   .I0(level4_in[2274]),
   .I1(level4_in[2275]),
   .I2(level4_in[2276]),
   .I3(level4_in[2277]),
   .I4(level4_in[2278]),
   .I5(level4_in[2279])
);

LUT6 #(
   .INIT(64'h8e86b3698e86b369)  
) LUT6_inst8156 (
   .O(to_level3[380]),
   .I0(level4_in[2280]),
   .I1(level4_in[2281]),
   .I2(level4_in[2282]),
   .I3(level4_in[2283]),
   .I4(level4_in[2284]),
   .I5(level4_in[2285])
);

LUT6 #(
   .INIT(64'h970a7955970a7955)  
) LUT6_inst8157 (
   .O(to_level3[381]),
   .I0(level4_in[2286]),
   .I1(level4_in[2287]),
   .I2(level4_in[2288]),
   .I3(level4_in[2289]),
   .I4(level4_in[2290]),
   .I5(level4_in[2291])
);

LUT6 #(
   .INIT(64'hff39c132ff39c132)  
) LUT6_inst8158 (
   .O(to_level3[382]),
   .I0(level4_in[2292]),
   .I1(level4_in[2293]),
   .I2(level4_in[2294]),
   .I3(level4_in[2295]),
   .I4(level4_in[2296]),
   .I5(level4_in[2297])
);

LUT6 #(
   .INIT(64'heaea58e6eaea58e6)  
) LUT6_inst8159 (
   .O(to_level3[383]),
   .I0(level4_in[2298]),
   .I1(level4_in[2299]),
   .I2(level4_in[2300]),
   .I3(level4_in[2301]),
   .I4(level4_in[2302]),
   .I5(level4_in[2303])
);

LUT6 #(
   .INIT(64'h20c4428920c44289)  
) LUT6_inst8160 (
   .O(to_level3[384]),
   .I0(level4_in[2304]),
   .I1(level4_in[2305]),
   .I2(level4_in[2306]),
   .I3(level4_in[2307]),
   .I4(level4_in[2308]),
   .I5(level4_in[2309])
);

LUT6 #(
   .INIT(64'haeb12a81aeb12a81)  
) LUT6_inst8161 (
   .O(to_level3[385]),
   .I0(level4_in[2310]),
   .I1(level4_in[2311]),
   .I2(level4_in[2312]),
   .I3(level4_in[2313]),
   .I4(level4_in[2314]),
   .I5(level4_in[2315])
);

LUT6 #(
   .INIT(64'hddb1715cddb1715c)  
) LUT6_inst8162 (
   .O(to_level3[386]),
   .I0(level4_in[2316]),
   .I1(level4_in[2317]),
   .I2(level4_in[2318]),
   .I3(level4_in[2319]),
   .I4(level4_in[2320]),
   .I5(level4_in[2321])
);

LUT6 #(
   .INIT(64'hb4315b90b4315b90)  
) LUT6_inst8163 (
   .O(to_level3[387]),
   .I0(level4_in[2322]),
   .I1(level4_in[2323]),
   .I2(level4_in[2324]),
   .I3(level4_in[2325]),
   .I4(level4_in[2326]),
   .I5(level4_in[2327])
);

LUT6 #(
   .INIT(64'h9f9435919f943591)  
) LUT6_inst8164 (
   .O(to_level3[388]),
   .I0(level4_in[2328]),
   .I1(level4_in[2329]),
   .I2(level4_in[2330]),
   .I3(level4_in[2331]),
   .I4(level4_in[2332]),
   .I5(level4_in[2333])
);

LUT6 #(
   .INIT(64'h29ac691c29ac691c)  
) LUT6_inst8165 (
   .O(to_level3[389]),
   .I0(level4_in[2334]),
   .I1(level4_in[2335]),
   .I2(level4_in[2336]),
   .I3(level4_in[2337]),
   .I4(level4_in[2338]),
   .I5(level4_in[2339])
);

LUT6 #(
   .INIT(64'h5c3967855c396785)  
) LUT6_inst8166 (
   .O(to_level3[390]),
   .I0(level4_in[2340]),
   .I1(level4_in[2341]),
   .I2(level4_in[2342]),
   .I3(level4_in[2343]),
   .I4(level4_in[2344]),
   .I5(level4_in[2345])
);

LUT6 #(
   .INIT(64'h1001b9d61001b9d6)  
) LUT6_inst8167 (
   .O(to_level3[391]),
   .I0(level4_in[2346]),
   .I1(level4_in[2347]),
   .I2(level4_in[2348]),
   .I3(level4_in[2349]),
   .I4(level4_in[2350]),
   .I5(level4_in[2351])
);

LUT6 #(
   .INIT(64'h2ca900d12ca900d1)  
) LUT6_inst8168 (
   .O(to_level3[392]),
   .I0(level4_in[2352]),
   .I1(level4_in[2353]),
   .I2(level4_in[2354]),
   .I3(level4_in[2355]),
   .I4(level4_in[2356]),
   .I5(level4_in[2357])
);

LUT6 #(
   .INIT(64'h1c60b5931c60b593)  
) LUT6_inst8169 (
   .O(to_level3[393]),
   .I0(level4_in[2358]),
   .I1(level4_in[2359]),
   .I2(level4_in[2360]),
   .I3(level4_in[2361]),
   .I4(level4_in[2362]),
   .I5(level4_in[2363])
);

LUT6 #(
   .INIT(64'h858a21a8858a21a8)  
) LUT6_inst8170 (
   .O(to_level3[394]),
   .I0(level4_in[2364]),
   .I1(level4_in[2365]),
   .I2(level4_in[2366]),
   .I3(level4_in[2367]),
   .I4(level4_in[2368]),
   .I5(level4_in[2369])
);

LUT6 #(
   .INIT(64'h1cac31151cac3115)  
) LUT6_inst8171 (
   .O(to_level3[395]),
   .I0(level4_in[2370]),
   .I1(level4_in[2371]),
   .I2(level4_in[2372]),
   .I3(level4_in[2373]),
   .I4(level4_in[2374]),
   .I5(level4_in[2375])
);

LUT6 #(
   .INIT(64'h53032abf53032abf)  
) LUT6_inst8172 (
   .O(to_level3[396]),
   .I0(level4_in[2376]),
   .I1(level4_in[2377]),
   .I2(level4_in[2378]),
   .I3(level4_in[2379]),
   .I4(level4_in[2380]),
   .I5(level4_in[2381])
);

LUT6 #(
   .INIT(64'hb30e3c56b30e3c56)  
) LUT6_inst8173 (
   .O(to_level3[397]),
   .I0(level4_in[2382]),
   .I1(level4_in[2383]),
   .I2(level4_in[2384]),
   .I3(level4_in[2385]),
   .I4(level4_in[2386]),
   .I5(level4_in[2387])
);

LUT6 #(
   .INIT(64'h660ada76660ada76)  
) LUT6_inst8174 (
   .O(to_level3[398]),
   .I0(level4_in[2388]),
   .I1(level4_in[2389]),
   .I2(level4_in[2390]),
   .I3(level4_in[2391]),
   .I4(level4_in[2392]),
   .I5(level4_in[2393])
);

LUT6 #(
   .INIT(64'h11e3429111e34291)  
) LUT6_inst8175 (
   .O(to_level3[399]),
   .I0(level4_in[2394]),
   .I1(level4_in[2395]),
   .I2(level4_in[2396]),
   .I3(level4_in[2397]),
   .I4(level4_in[2398]),
   .I5(level4_in[2399])
);

LUT6 #(
   .INIT(64'he94d7645e94d7645)  
) LUT6_inst8176 (
   .O(to_level3[400]),
   .I0(level4_in[2400]),
   .I1(level4_in[2401]),
   .I2(level4_in[2402]),
   .I3(level4_in[2403]),
   .I4(level4_in[2404]),
   .I5(level4_in[2405])
);

LUT6 #(
   .INIT(64'h41139fac41139fac)  
) LUT6_inst8177 (
   .O(to_level3[401]),
   .I0(level4_in[2406]),
   .I1(level4_in[2407]),
   .I2(level4_in[2408]),
   .I3(level4_in[2409]),
   .I4(level4_in[2410]),
   .I5(level4_in[2411])
);

LUT6 #(
   .INIT(64'h396c2293396c2293)  
) LUT6_inst8178 (
   .O(to_level3[402]),
   .I0(level4_in[2412]),
   .I1(level4_in[2413]),
   .I2(level4_in[2414]),
   .I3(level4_in[2415]),
   .I4(level4_in[2416]),
   .I5(level4_in[2417])
);

LUT6 #(
   .INIT(64'h5eff0db25eff0db2)  
) LUT6_inst8179 (
   .O(to_level3[403]),
   .I0(level4_in[2418]),
   .I1(level4_in[2419]),
   .I2(level4_in[2420]),
   .I3(level4_in[2421]),
   .I4(level4_in[2422]),
   .I5(level4_in[2423])
);

LUT6 #(
   .INIT(64'h9931adc29931adc2)  
) LUT6_inst8180 (
   .O(to_level3[404]),
   .I0(level4_in[2424]),
   .I1(level4_in[2425]),
   .I2(level4_in[2426]),
   .I3(level4_in[2427]),
   .I4(level4_in[2428]),
   .I5(level4_in[2429])
);

LUT6 #(
   .INIT(64'h53685dcd53685dcd)  
) LUT6_inst8181 (
   .O(to_level3[405]),
   .I0(level4_in[2430]),
   .I1(level4_in[2431]),
   .I2(level4_in[2432]),
   .I3(level4_in[2433]),
   .I4(level4_in[2434]),
   .I5(level4_in[2435])
);

LUT6 #(
   .INIT(64'h6fbea7a86fbea7a8)  
) LUT6_inst8182 (
   .O(to_level3[406]),
   .I0(level4_in[2436]),
   .I1(level4_in[2437]),
   .I2(level4_in[2438]),
   .I3(level4_in[2439]),
   .I4(level4_in[2440]),
   .I5(level4_in[2441])
);

LUT6 #(
   .INIT(64'h8d5a21938d5a2193)  
) LUT6_inst8183 (
   .O(to_level3[407]),
   .I0(level4_in[2442]),
   .I1(level4_in[2443]),
   .I2(level4_in[2444]),
   .I3(level4_in[2445]),
   .I4(level4_in[2446]),
   .I5(level4_in[2447])
);

LUT6 #(
   .INIT(64'h5824e3295824e329)  
) LUT6_inst8184 (
   .O(to_level3[408]),
   .I0(level4_in[2448]),
   .I1(level4_in[2449]),
   .I2(level4_in[2450]),
   .I3(level4_in[2451]),
   .I4(level4_in[2452]),
   .I5(level4_in[2453])
);

LUT6 #(
   .INIT(64'h7e5467d97e5467d9)  
) LUT6_inst8185 (
   .O(to_level3[409]),
   .I0(level4_in[2454]),
   .I1(level4_in[2455]),
   .I2(level4_in[2456]),
   .I3(level4_in[2457]),
   .I4(level4_in[2458]),
   .I5(level4_in[2459])
);

LUT6 #(
   .INIT(64'h8f7c67038f7c6703)  
) LUT6_inst8186 (
   .O(to_level3[410]),
   .I0(level4_in[2460]),
   .I1(level4_in[2461]),
   .I2(level4_in[2462]),
   .I3(level4_in[2463]),
   .I4(level4_in[2464]),
   .I5(level4_in[2465])
);

LUT6 #(
   .INIT(64'h4f1710454f171045)  
) LUT6_inst8187 (
   .O(to_level3[411]),
   .I0(level4_in[2466]),
   .I1(level4_in[2467]),
   .I2(level4_in[2468]),
   .I3(level4_in[2469]),
   .I4(level4_in[2470]),
   .I5(level4_in[2471])
);

LUT6 #(
   .INIT(64'h65e7405365e74053)  
) LUT6_inst8188 (
   .O(to_level3[412]),
   .I0(level4_in[2472]),
   .I1(level4_in[2473]),
   .I2(level4_in[2474]),
   .I3(level4_in[2475]),
   .I4(level4_in[2476]),
   .I5(level4_in[2477])
);

LUT6 #(
   .INIT(64'h807aaec2807aaec2)  
) LUT6_inst8189 (
   .O(to_level3[413]),
   .I0(level4_in[2478]),
   .I1(level4_in[2479]),
   .I2(level4_in[2480]),
   .I3(level4_in[2481]),
   .I4(level4_in[2482]),
   .I5(level4_in[2483])
);

LUT6 #(
   .INIT(64'h4daf23254daf2325)  
) LUT6_inst8190 (
   .O(to_level3[414]),
   .I0(level4_in[2484]),
   .I1(level4_in[2485]),
   .I2(level4_in[2486]),
   .I3(level4_in[2487]),
   .I4(level4_in[2488]),
   .I5(level4_in[2489])
);

LUT6 #(
   .INIT(64'h8e98ecbd8e98ecbd)  
) LUT6_inst8191 (
   .O(to_level3[415]),
   .I0(level4_in[2490]),
   .I1(level4_in[2491]),
   .I2(level4_in[2492]),
   .I3(level4_in[2493]),
   .I4(level4_in[2494]),
   .I5(level4_in[2495])
);

LUT6 #(
   .INIT(64'h06884c3b06884c3b)  
) LUT6_inst8192 (
   .O(to_level3[416]),
   .I0(level4_in[2496]),
   .I1(level4_in[2497]),
   .I2(level4_in[2498]),
   .I3(level4_in[2499]),
   .I4(level4_in[2500]),
   .I5(level4_in[2501])
);

LUT6 #(
   .INIT(64'h70e955af70e955af)  
) LUT6_inst8193 (
   .O(to_level3[417]),
   .I0(level4_in[2502]),
   .I1(level4_in[2503]),
   .I2(level4_in[2504]),
   .I3(level4_in[2505]),
   .I4(level4_in[2506]),
   .I5(level4_in[2507])
);

LUT6 #(
   .INIT(64'h7389685573896855)  
) LUT6_inst8194 (
   .O(to_level3[418]),
   .I0(level4_in[2508]),
   .I1(level4_in[2509]),
   .I2(level4_in[2510]),
   .I3(level4_in[2511]),
   .I4(level4_in[2512]),
   .I5(level4_in[2513])
);

LUT6 #(
   .INIT(64'h5d9b35d65d9b35d6)  
) LUT6_inst8195 (
   .O(to_level3[419]),
   .I0(level4_in[2514]),
   .I1(level4_in[2515]),
   .I2(level4_in[2516]),
   .I3(level4_in[2517]),
   .I4(level4_in[2518]),
   .I5(level4_in[2519])
);

LUT6 #(
   .INIT(64'h98932e6198932e61)  
) LUT6_inst8196 (
   .O(to_level3[420]),
   .I0(level4_in[2520]),
   .I1(level4_in[2521]),
   .I2(level4_in[2522]),
   .I3(level4_in[2523]),
   .I4(level4_in[2524]),
   .I5(level4_in[2525])
);

LUT6 #(
   .INIT(64'h5b4d9d3d5b4d9d3d)  
) LUT6_inst8197 (
   .O(to_level3[421]),
   .I0(level4_in[2526]),
   .I1(level4_in[2527]),
   .I2(level4_in[2528]),
   .I3(level4_in[2529]),
   .I4(level4_in[2530]),
   .I5(level4_in[2531])
);

LUT6 #(
   .INIT(64'h42dd29bf42dd29bf)  
) LUT6_inst8198 (
   .O(to_level3[422]),
   .I0(level4_in[2532]),
   .I1(level4_in[2533]),
   .I2(level4_in[2534]),
   .I3(level4_in[2535]),
   .I4(level4_in[2536]),
   .I5(level4_in[2537])
);

LUT6 #(
   .INIT(64'hd5697f6cd5697f6c)  
) LUT6_inst8199 (
   .O(to_level3[423]),
   .I0(level4_in[2538]),
   .I1(level4_in[2539]),
   .I2(level4_in[2540]),
   .I3(level4_in[2541]),
   .I4(level4_in[2542]),
   .I5(level4_in[2543])
);

LUT6 #(
   .INIT(64'hc2eed0acc2eed0ac)  
) LUT6_inst8200 (
   .O(to_level3[424]),
   .I0(level4_in[2544]),
   .I1(level4_in[2545]),
   .I2(level4_in[2546]),
   .I3(level4_in[2547]),
   .I4(level4_in[2548]),
   .I5(level4_in[2549])
);

LUT6 #(
   .INIT(64'h795e193c795e193c)  
) LUT6_inst8201 (
   .O(to_level3[425]),
   .I0(level4_in[2550]),
   .I1(level4_in[2551]),
   .I2(level4_in[2552]),
   .I3(level4_in[2553]),
   .I4(level4_in[2554]),
   .I5(level4_in[2555])
);

LUT6 #(
   .INIT(64'hb7c72561b7c72561)  
) LUT6_inst8202 (
   .O(to_level3[426]),
   .I0(level4_in[2556]),
   .I1(level4_in[2557]),
   .I2(level4_in[2558]),
   .I3(level4_in[2559]),
   .I4(level4_in[2560]),
   .I5(level4_in[2561])
);

LUT6 #(
   .INIT(64'h6c89bd236c89bd23)  
) LUT6_inst8203 (
   .O(to_level3[427]),
   .I0(level4_in[2562]),
   .I1(level4_in[2563]),
   .I2(level4_in[2564]),
   .I3(level4_in[2565]),
   .I4(level4_in[2566]),
   .I5(level4_in[2567])
);

LUT6 #(
   .INIT(64'h46fdeb7546fdeb75)  
) LUT6_inst8204 (
   .O(to_level3[428]),
   .I0(level4_in[2568]),
   .I1(level4_in[2569]),
   .I2(level4_in[2570]),
   .I3(level4_in[2571]),
   .I4(level4_in[2572]),
   .I5(level4_in[2573])
);

LUT6 #(
   .INIT(64'h49801d4049801d40)  
) LUT6_inst8205 (
   .O(to_level3[429]),
   .I0(level4_in[2574]),
   .I1(level4_in[2575]),
   .I2(level4_in[2576]),
   .I3(level4_in[2577]),
   .I4(level4_in[2578]),
   .I5(level4_in[2579])
);

LUT6 #(
   .INIT(64'h35d2cf5f35d2cf5f)  
) LUT6_inst8206 (
   .O(to_level3[430]),
   .I0(level4_in[2580]),
   .I1(level4_in[2581]),
   .I2(level4_in[2582]),
   .I3(level4_in[2583]),
   .I4(level4_in[2584]),
   .I5(level4_in[2585])
);

LUT6 #(
   .INIT(64'h8b1e82a28b1e82a2)  
) LUT6_inst8207 (
   .O(to_level3[431]),
   .I0(level4_in[2586]),
   .I1(level4_in[2587]),
   .I2(level4_in[2588]),
   .I3(level4_in[2589]),
   .I4(level4_in[2590]),
   .I5(level4_in[2591])
);

LUT6 #(
   .INIT(64'h1971974a1971974a)  
) LUT6_inst8208 (
   .O(to_level3[432]),
   .I0(level4_in[2592]),
   .I1(level4_in[2593]),
   .I2(level4_in[2594]),
   .I3(level4_in[2595]),
   .I4(level4_in[2596]),
   .I5(level4_in[2597])
);

LUT6 #(
   .INIT(64'h5487bb035487bb03)  
) LUT6_inst8209 (
   .O(to_level3[433]),
   .I0(level4_in[2598]),
   .I1(level4_in[2599]),
   .I2(level4_in[2600]),
   .I3(level4_in[2601]),
   .I4(level4_in[2602]),
   .I5(level4_in[2603])
);

LUT6 #(
   .INIT(64'h49f4188349f41883)  
) LUT6_inst8210 (
   .O(to_level3[434]),
   .I0(level4_in[2604]),
   .I1(level4_in[2605]),
   .I2(level4_in[2606]),
   .I3(level4_in[2607]),
   .I4(level4_in[2608]),
   .I5(level4_in[2609])
);

LUT6 #(
   .INIT(64'hd9774274d9774274)  
) LUT6_inst8211 (
   .O(to_level3[435]),
   .I0(level4_in[2610]),
   .I1(level4_in[2611]),
   .I2(level4_in[2612]),
   .I3(level4_in[2613]),
   .I4(level4_in[2614]),
   .I5(level4_in[2615])
);

LUT6 #(
   .INIT(64'h4d75af8e4d75af8e)  
) LUT6_inst8212 (
   .O(to_level3[436]),
   .I0(level4_in[2616]),
   .I1(level4_in[2617]),
   .I2(level4_in[2618]),
   .I3(level4_in[2619]),
   .I4(level4_in[2620]),
   .I5(level4_in[2621])
);

LUT6 #(
   .INIT(64'h5b6e99d35b6e99d3)  
) LUT6_inst8213 (
   .O(to_level3[437]),
   .I0(level4_in[2622]),
   .I1(level4_in[2623]),
   .I2(level4_in[2624]),
   .I3(level4_in[2625]),
   .I4(level4_in[2626]),
   .I5(level4_in[2627])
);

LUT6 #(
   .INIT(64'h8770c1c88770c1c8)  
) LUT6_inst8214 (
   .O(to_level3[438]),
   .I0(level4_in[2628]),
   .I1(level4_in[2629]),
   .I2(level4_in[2630]),
   .I3(level4_in[2631]),
   .I4(level4_in[2632]),
   .I5(level4_in[2633])
);

LUT6 #(
   .INIT(64'h317201e9317201e9)  
) LUT6_inst8215 (
   .O(to_level3[439]),
   .I0(level4_in[2634]),
   .I1(level4_in[2635]),
   .I2(level4_in[2636]),
   .I3(level4_in[2637]),
   .I4(level4_in[2638]),
   .I5(level4_in[2639])
);

LUT6 #(
   .INIT(64'hfba3ce59fba3ce59)  
) LUT6_inst8216 (
   .O(to_level3[440]),
   .I0(level4_in[2640]),
   .I1(level4_in[2641]),
   .I2(level4_in[2642]),
   .I3(level4_in[2643]),
   .I4(level4_in[2644]),
   .I5(level4_in[2645])
);

LUT6 #(
   .INIT(64'h36c00a3236c00a32)  
) LUT6_inst8217 (
   .O(to_level3[441]),
   .I0(level4_in[2646]),
   .I1(level4_in[2647]),
   .I2(level4_in[2648]),
   .I3(level4_in[2649]),
   .I4(level4_in[2650]),
   .I5(level4_in[2651])
);

LUT6 #(
   .INIT(64'hcd363fb1cd363fb1)  
) LUT6_inst8218 (
   .O(to_level3[442]),
   .I0(level4_in[2652]),
   .I1(level4_in[2653]),
   .I2(level4_in[2654]),
   .I3(level4_in[2655]),
   .I4(level4_in[2656]),
   .I5(level4_in[2657])
);

LUT6 #(
   .INIT(64'h9a5555579a555557)  
) LUT6_inst8219 (
   .O(to_level3[443]),
   .I0(level4_in[2658]),
   .I1(level4_in[2659]),
   .I2(level4_in[2660]),
   .I3(level4_in[2661]),
   .I4(level4_in[2662]),
   .I5(level4_in[2663])
);

LUT6 #(
   .INIT(64'ha5f20f05a5f20f05)  
) LUT6_inst8220 (
   .O(to_level3[444]),
   .I0(level4_in[2664]),
   .I1(level4_in[2665]),
   .I2(level4_in[2666]),
   .I3(level4_in[2667]),
   .I4(level4_in[2668]),
   .I5(level4_in[2669])
);

LUT6 #(
   .INIT(64'h1685044716850447)  
) LUT6_inst8221 (
   .O(to_level3[445]),
   .I0(level4_in[2670]),
   .I1(level4_in[2671]),
   .I2(level4_in[2672]),
   .I3(level4_in[2673]),
   .I4(level4_in[2674]),
   .I5(level4_in[2675])
);

LUT6 #(
   .INIT(64'hf0507514f0507514)  
) LUT6_inst8222 (
   .O(to_level3[446]),
   .I0(level4_in[2676]),
   .I1(level4_in[2677]),
   .I2(level4_in[2678]),
   .I3(level4_in[2679]),
   .I4(level4_in[2680]),
   .I5(level4_in[2681])
);

LUT6 #(
   .INIT(64'h11c7930611c79306)  
) LUT6_inst8223 (
   .O(to_level3[447]),
   .I0(level4_in[2682]),
   .I1(level4_in[2683]),
   .I2(level4_in[2684]),
   .I3(level4_in[2685]),
   .I4(level4_in[2686]),
   .I5(level4_in[2687])
);

LUT6 #(
   .INIT(64'hd4b24d93d4b24d93)  
) LUT6_inst8224 (
   .O(to_level3[448]),
   .I0(level4_in[2688]),
   .I1(level4_in[2689]),
   .I2(level4_in[2690]),
   .I3(level4_in[2691]),
   .I4(level4_in[2692]),
   .I5(level4_in[2693])
);

LUT6 #(
   .INIT(64'h081f2e4e081f2e4e)  
) LUT6_inst8225 (
   .O(to_level3[449]),
   .I0(level4_in[2694]),
   .I1(level4_in[2695]),
   .I2(level4_in[2696]),
   .I3(level4_in[2697]),
   .I4(level4_in[2698]),
   .I5(level4_in[2699])
);

LUT6 #(
   .INIT(64'h4e69164a4e69164a)  
) LUT6_inst8226 (
   .O(to_level3[450]),
   .I0(level4_in[2700]),
   .I1(level4_in[2701]),
   .I2(level4_in[2702]),
   .I3(level4_in[2703]),
   .I4(level4_in[2704]),
   .I5(level4_in[2705])
);

LUT6 #(
   .INIT(64'h0cc8a0130cc8a013)  
) LUT6_inst8227 (
   .O(to_level3[451]),
   .I0(level4_in[2706]),
   .I1(level4_in[2707]),
   .I2(level4_in[2708]),
   .I3(level4_in[2709]),
   .I4(level4_in[2710]),
   .I5(level4_in[2711])
);

LUT6 #(
   .INIT(64'h3bb315083bb31508)  
) LUT6_inst8228 (
   .O(to_level3[452]),
   .I0(level4_in[2712]),
   .I1(level4_in[2713]),
   .I2(level4_in[2714]),
   .I3(level4_in[2715]),
   .I4(level4_in[2716]),
   .I5(level4_in[2717])
);

LUT6 #(
   .INIT(64'h7c1ecc567c1ecc56)  
) LUT6_inst8229 (
   .O(to_level3[453]),
   .I0(level4_in[2718]),
   .I1(level4_in[2719]),
   .I2(level4_in[2720]),
   .I3(level4_in[2721]),
   .I4(level4_in[2722]),
   .I5(level4_in[2723])
);

LUT6 #(
   .INIT(64'hef5476d3ef5476d3)  
) LUT6_inst8230 (
   .O(to_level3[454]),
   .I0(level4_in[2724]),
   .I1(level4_in[2725]),
   .I2(level4_in[2726]),
   .I3(level4_in[2727]),
   .I4(level4_in[2728]),
   .I5(level4_in[2729])
);

LUT6 #(
   .INIT(64'hcbd73482cbd73482)  
) LUT6_inst8231 (
   .O(to_level3[455]),
   .I0(level4_in[2730]),
   .I1(level4_in[2731]),
   .I2(level4_in[2732]),
   .I3(level4_in[2733]),
   .I4(level4_in[2734]),
   .I5(level4_in[2735])
);

LUT6 #(
   .INIT(64'ha52f823ea52f823e)  
) LUT6_inst8232 (
   .O(to_level3[456]),
   .I0(level4_in[2736]),
   .I1(level4_in[2737]),
   .I2(level4_in[2738]),
   .I3(level4_in[2739]),
   .I4(level4_in[2740]),
   .I5(level4_in[2741])
);

LUT6 #(
   .INIT(64'heecfc654eecfc654)  
) LUT6_inst8233 (
   .O(to_level3[457]),
   .I0(level4_in[2742]),
   .I1(level4_in[2743]),
   .I2(level4_in[2744]),
   .I3(level4_in[2745]),
   .I4(level4_in[2746]),
   .I5(level4_in[2747])
);

LUT6 #(
   .INIT(64'h52939b1352939b13)  
) LUT6_inst8234 (
   .O(to_level3[458]),
   .I0(level4_in[2748]),
   .I1(level4_in[2749]),
   .I2(level4_in[2750]),
   .I3(level4_in[2751]),
   .I4(level4_in[2752]),
   .I5(level4_in[2753])
);

LUT6 #(
   .INIT(64'h04cf755704cf7557)  
) LUT6_inst8235 (
   .O(to_level3[459]),
   .I0(level4_in[2754]),
   .I1(level4_in[2755]),
   .I2(level4_in[2756]),
   .I3(level4_in[2757]),
   .I4(level4_in[2758]),
   .I5(level4_in[2759])
);

LUT6 #(
   .INIT(64'h25af730125af7301)  
) LUT6_inst8236 (
   .O(to_level3[460]),
   .I0(level4_in[2760]),
   .I1(level4_in[2761]),
   .I2(level4_in[2762]),
   .I3(level4_in[2763]),
   .I4(level4_in[2764]),
   .I5(level4_in[2765])
);

LUT6 #(
   .INIT(64'h02bac35002bac350)  
) LUT6_inst8237 (
   .O(to_level3[461]),
   .I0(level4_in[2766]),
   .I1(level4_in[2767]),
   .I2(level4_in[2768]),
   .I3(level4_in[2769]),
   .I4(level4_in[2770]),
   .I5(level4_in[2771])
);

LUT6 #(
   .INIT(64'h1ef419411ef41941)  
) LUT6_inst8238 (
   .O(to_level3[462]),
   .I0(level4_in[2772]),
   .I1(level4_in[2773]),
   .I2(level4_in[2774]),
   .I3(level4_in[2775]),
   .I4(level4_in[2776]),
   .I5(level4_in[2777])
);

LUT6 #(
   .INIT(64'h78e67b5078e67b50)  
) LUT6_inst8239 (
   .O(to_level3[463]),
   .I0(level4_in[2778]),
   .I1(level4_in[2779]),
   .I2(level4_in[2780]),
   .I3(level4_in[2781]),
   .I4(level4_in[2782]),
   .I5(level4_in[2783])
);

LUT6 #(
   .INIT(64'he8174414e8174414)  
) LUT6_inst8240 (
   .O(to_level3[464]),
   .I0(level4_in[2784]),
   .I1(level4_in[2785]),
   .I2(level4_in[2786]),
   .I3(level4_in[2787]),
   .I4(level4_in[2788]),
   .I5(level4_in[2789])
);

LUT6 #(
   .INIT(64'ha3e50af8a3e50af8)  
) LUT6_inst8241 (
   .O(to_level3[465]),
   .I0(level4_in[2790]),
   .I1(level4_in[2791]),
   .I2(level4_in[2792]),
   .I3(level4_in[2793]),
   .I4(level4_in[2794]),
   .I5(level4_in[2795])
);

LUT6 #(
   .INIT(64'h0391489a0391489a)  
) LUT6_inst8242 (
   .O(to_level3[466]),
   .I0(level4_in[2796]),
   .I1(level4_in[2797]),
   .I2(level4_in[2798]),
   .I3(level4_in[2799]),
   .I4(level4_in[2800]),
   .I5(level4_in[2801])
);

LUT6 #(
   .INIT(64'hf0d0ad4bf0d0ad4b)  
) LUT6_inst8243 (
   .O(to_level3[467]),
   .I0(level4_in[2802]),
   .I1(level4_in[2803]),
   .I2(level4_in[2804]),
   .I3(level4_in[2805]),
   .I4(level4_in[2806]),
   .I5(level4_in[2807])
);

LUT6 #(
   .INIT(64'h2107340f2107340f)  
) LUT6_inst8244 (
   .O(to_level3[468]),
   .I0(level4_in[2808]),
   .I1(level4_in[2809]),
   .I2(level4_in[2810]),
   .I3(level4_in[2811]),
   .I4(level4_in[2812]),
   .I5(level4_in[2813])
);

LUT6 #(
   .INIT(64'hd7a1651dd7a1651d)  
) LUT6_inst8245 (
   .O(to_level3[469]),
   .I0(level4_in[2814]),
   .I1(level4_in[2815]),
   .I2(level4_in[2816]),
   .I3(level4_in[2817]),
   .I4(level4_in[2818]),
   .I5(level4_in[2819])
);

LUT6 #(
   .INIT(64'hfb221cf0fb221cf0)  
) LUT6_inst8246 (
   .O(to_level3[470]),
   .I0(level4_in[2820]),
   .I1(level4_in[2821]),
   .I2(level4_in[2822]),
   .I3(level4_in[2823]),
   .I4(level4_in[2824]),
   .I5(level4_in[2825])
);

LUT6 #(
   .INIT(64'hbbcd54dcbbcd54dc)  
) LUT6_inst8247 (
   .O(to_level3[471]),
   .I0(level4_in[2826]),
   .I1(level4_in[2827]),
   .I2(level4_in[2828]),
   .I3(level4_in[2829]),
   .I4(level4_in[2830]),
   .I5(level4_in[2831])
);

LUT6 #(
   .INIT(64'h7f2c015b7f2c015b)  
) LUT6_inst8248 (
   .O(to_level3[472]),
   .I0(level4_in[2832]),
   .I1(level4_in[2833]),
   .I2(level4_in[2834]),
   .I3(level4_in[2835]),
   .I4(level4_in[2836]),
   .I5(level4_in[2837])
);

LUT6 #(
   .INIT(64'h9bbd9a379bbd9a37)  
) LUT6_inst8249 (
   .O(to_level3[473]),
   .I0(level4_in[2838]),
   .I1(level4_in[2839]),
   .I2(level4_in[2840]),
   .I3(level4_in[2841]),
   .I4(level4_in[2842]),
   .I5(level4_in[2843])
);

LUT6 #(
   .INIT(64'hf7aa2d86f7aa2d86)  
) LUT6_inst8250 (
   .O(to_level3[474]),
   .I0(level4_in[2844]),
   .I1(level4_in[2845]),
   .I2(level4_in[2846]),
   .I3(level4_in[2847]),
   .I4(level4_in[2848]),
   .I5(level4_in[2849])
);

LUT6 #(
   .INIT(64'hd31a7aacd31a7aac)  
) LUT6_inst8251 (
   .O(to_level3[475]),
   .I0(level4_in[2850]),
   .I1(level4_in[2851]),
   .I2(level4_in[2852]),
   .I3(level4_in[2853]),
   .I4(level4_in[2854]),
   .I5(level4_in[2855])
);

LUT6 #(
   .INIT(64'h66c11b8966c11b89)  
) LUT6_inst8252 (
   .O(to_level3[476]),
   .I0(level4_in[2856]),
   .I1(level4_in[2857]),
   .I2(level4_in[2858]),
   .I3(level4_in[2859]),
   .I4(level4_in[2860]),
   .I5(level4_in[2861])
);

LUT6 #(
   .INIT(64'h5464b5e05464b5e0)  
) LUT6_inst8253 (
   .O(to_level3[477]),
   .I0(level4_in[2862]),
   .I1(level4_in[2863]),
   .I2(level4_in[2864]),
   .I3(level4_in[2865]),
   .I4(level4_in[2866]),
   .I5(level4_in[2867])
);

LUT6 #(
   .INIT(64'h4178a2184178a218)  
) LUT6_inst8254 (
   .O(to_level3[478]),
   .I0(level4_in[2868]),
   .I1(level4_in[2869]),
   .I2(level4_in[2870]),
   .I3(level4_in[2871]),
   .I4(level4_in[2872]),
   .I5(level4_in[2873])
);

LUT6 #(
   .INIT(64'hbbbf8718bbbf8718)  
) LUT6_inst8255 (
   .O(to_level3[479]),
   .I0(level4_in[2874]),
   .I1(level4_in[2875]),
   .I2(level4_in[2876]),
   .I3(level4_in[2877]),
   .I4(level4_in[2878]),
   .I5(level4_in[2879])
);

LUT6 #(
   .INIT(64'hd56b70cdd56b70cd)  
) LUT6_inst8256 (
   .O(to_level3[480]),
   .I0(level4_in[2880]),
   .I1(level4_in[2881]),
   .I2(level4_in[2882]),
   .I3(level4_in[2883]),
   .I4(level4_in[2884]),
   .I5(level4_in[2885])
);

LUT6 #(
   .INIT(64'h703cae97703cae97)  
) LUT6_inst8257 (
   .O(to_level3[481]),
   .I0(level4_in[2886]),
   .I1(level4_in[2887]),
   .I2(level4_in[2888]),
   .I3(level4_in[2889]),
   .I4(level4_in[2890]),
   .I5(level4_in[2891])
);

LUT6 #(
   .INIT(64'h3a69a3633a69a363)  
) LUT6_inst8258 (
   .O(to_level3[482]),
   .I0(level4_in[2892]),
   .I1(level4_in[2893]),
   .I2(level4_in[2894]),
   .I3(level4_in[2895]),
   .I4(level4_in[2896]),
   .I5(level4_in[2897])
);

LUT6 #(
   .INIT(64'hece2b682ece2b682)  
) LUT6_inst8259 (
   .O(to_level3[483]),
   .I0(level4_in[2898]),
   .I1(level4_in[2899]),
   .I2(level4_in[2900]),
   .I3(level4_in[2901]),
   .I4(level4_in[2902]),
   .I5(level4_in[2903])
);

LUT6 #(
   .INIT(64'ha22d0270a22d0270)  
) LUT6_inst8260 (
   .O(to_level3[484]),
   .I0(level4_in[2904]),
   .I1(level4_in[2905]),
   .I2(level4_in[2906]),
   .I3(level4_in[2907]),
   .I4(level4_in[2908]),
   .I5(level4_in[2909])
);

LUT6 #(
   .INIT(64'h963a00a0963a00a0)  
) LUT6_inst8261 (
   .O(to_level3[485]),
   .I0(level4_in[2910]),
   .I1(level4_in[2911]),
   .I2(level4_in[2912]),
   .I3(level4_in[2913]),
   .I4(level4_in[2914]),
   .I5(level4_in[2915])
);

LUT6 #(
   .INIT(64'h6dc7982c6dc7982c)  
) LUT6_inst8262 (
   .O(to_level3[486]),
   .I0(level4_in[2916]),
   .I1(level4_in[2917]),
   .I2(level4_in[2918]),
   .I3(level4_in[2919]),
   .I4(level4_in[2920]),
   .I5(level4_in[2921])
);

LUT6 #(
   .INIT(64'h1a76f0501a76f050)  
) LUT6_inst8263 (
   .O(to_level3[487]),
   .I0(level4_in[2922]),
   .I1(level4_in[2923]),
   .I2(level4_in[2924]),
   .I3(level4_in[2925]),
   .I4(level4_in[2926]),
   .I5(level4_in[2927])
);

LUT6 #(
   .INIT(64'hfc7720bffc7720bf)  
) LUT6_inst8264 (
   .O(to_level3[488]),
   .I0(level4_in[2928]),
   .I1(level4_in[2929]),
   .I2(level4_in[2930]),
   .I3(level4_in[2931]),
   .I4(level4_in[2932]),
   .I5(level4_in[2933])
);

LUT6 #(
   .INIT(64'h76def53476def534)  
) LUT6_inst8265 (
   .O(to_level3[489]),
   .I0(level4_in[2934]),
   .I1(level4_in[2935]),
   .I2(level4_in[2936]),
   .I3(level4_in[2937]),
   .I4(level4_in[2938]),
   .I5(level4_in[2939])
);

LUT6 #(
   .INIT(64'h6f26bbf96f26bbf9)  
) LUT6_inst8266 (
   .O(to_level3[490]),
   .I0(level4_in[2940]),
   .I1(level4_in[2941]),
   .I2(level4_in[2942]),
   .I3(level4_in[2943]),
   .I4(level4_in[2944]),
   .I5(level4_in[2945])
);

LUT6 #(
   .INIT(64'h2079b1bc2079b1bc)  
) LUT6_inst8267 (
   .O(to_level3[491]),
   .I0(level4_in[2946]),
   .I1(level4_in[2947]),
   .I2(level4_in[2948]),
   .I3(level4_in[2949]),
   .I4(level4_in[2950]),
   .I5(level4_in[2951])
);

LUT6 #(
   .INIT(64'h1b23cc7c1b23cc7c)  
) LUT6_inst8268 (
   .O(to_level3[492]),
   .I0(level4_in[2952]),
   .I1(level4_in[2953]),
   .I2(level4_in[2954]),
   .I3(level4_in[2955]),
   .I4(level4_in[2956]),
   .I5(level4_in[2957])
);

LUT6 #(
   .INIT(64'h16c5489f16c5489f)  
) LUT6_inst8269 (
   .O(to_level3[493]),
   .I0(level4_in[2958]),
   .I1(level4_in[2959]),
   .I2(level4_in[2960]),
   .I3(level4_in[2961]),
   .I4(level4_in[2962]),
   .I5(level4_in[2963])
);

LUT6 #(
   .INIT(64'h1998046619980466)  
) LUT6_inst8270 (
   .O(to_level3[494]),
   .I0(level4_in[2964]),
   .I1(level4_in[2965]),
   .I2(level4_in[2966]),
   .I3(level4_in[2967]),
   .I4(level4_in[2968]),
   .I5(level4_in[2969])
);

LUT6 #(
   .INIT(64'h026535b6026535b6)  
) LUT6_inst8271 (
   .O(to_level3[495]),
   .I0(level4_in[2970]),
   .I1(level4_in[2971]),
   .I2(level4_in[2972]),
   .I3(level4_in[2973]),
   .I4(level4_in[2974]),
   .I5(level4_in[2975])
);

LUT6 #(
   .INIT(64'h5e6ac7cd5e6ac7cd)  
) LUT6_inst8272 (
   .O(to_level3[496]),
   .I0(level4_in[2976]),
   .I1(level4_in[2977]),
   .I2(level4_in[2978]),
   .I3(level4_in[2979]),
   .I4(level4_in[2980]),
   .I5(level4_in[2981])
);

LUT6 #(
   .INIT(64'h786886a3786886a3)  
) LUT6_inst8273 (
   .O(to_level3[497]),
   .I0(level4_in[2982]),
   .I1(level4_in[2983]),
   .I2(level4_in[2984]),
   .I3(level4_in[2985]),
   .I4(level4_in[2986]),
   .I5(level4_in[2987])
);

LUT6 #(
   .INIT(64'h828cfdb4828cfdb4)  
) LUT6_inst8274 (
   .O(to_level3[498]),
   .I0(level4_in[2988]),
   .I1(level4_in[2989]),
   .I2(level4_in[2990]),
   .I3(level4_in[2991]),
   .I4(level4_in[2992]),
   .I5(level4_in[2993])
);

LUT6 #(
   .INIT(64'hec433751ec433751)  
) LUT6_inst8275 (
   .O(to_level3[499]),
   .I0(level4_in[2994]),
   .I1(level4_in[2995]),
   .I2(level4_in[2996]),
   .I3(level4_in[2997]),
   .I4(level4_in[2998]),
   .I5(level4_in[2999])
);

LUT6 #(
   .INIT(64'h6ff1647c6ff1647c)  
) LUT6_inst8276 (
   .O(to_level3[500]),
   .I0(level4_in[3000]),
   .I1(level4_in[3001]),
   .I2(level4_in[3002]),
   .I3(level4_in[3003]),
   .I4(level4_in[3004]),
   .I5(level4_in[3005])
);

LUT6 #(
   .INIT(64'hd23ceb86d23ceb86)  
) LUT6_inst8277 (
   .O(to_level3[501]),
   .I0(level4_in[3006]),
   .I1(level4_in[3007]),
   .I2(level4_in[3008]),
   .I3(level4_in[3009]),
   .I4(level4_in[3010]),
   .I5(level4_in[3011])
);

LUT6 #(
   .INIT(64'hc6ddc168c6ddc168)  
) LUT6_inst8278 (
   .O(to_level3[502]),
   .I0(level4_in[3012]),
   .I1(level4_in[3013]),
   .I2(level4_in[3014]),
   .I3(level4_in[3015]),
   .I4(level4_in[3016]),
   .I5(level4_in[3017])
);

LUT6 #(
   .INIT(64'h1346549513465495)  
) LUT6_inst8279 (
   .O(to_level3[503]),
   .I0(level4_in[3018]),
   .I1(level4_in[3019]),
   .I2(level4_in[3020]),
   .I3(level4_in[3021]),
   .I4(level4_in[3022]),
   .I5(level4_in[3023])
);

LUT6 #(
   .INIT(64'hedd9c54aedd9c54a)  
) LUT6_inst8280 (
   .O(to_level3[504]),
   .I0(level4_in[3024]),
   .I1(level4_in[3025]),
   .I2(level4_in[3026]),
   .I3(level4_in[3027]),
   .I4(level4_in[3028]),
   .I5(level4_in[3029])
);

LUT6 #(
   .INIT(64'ha85532f2a85532f2)  
) LUT6_inst8281 (
   .O(to_level3[505]),
   .I0(level4_in[3030]),
   .I1(level4_in[3031]),
   .I2(level4_in[3032]),
   .I3(level4_in[3033]),
   .I4(level4_in[3034]),
   .I5(level4_in[3035])
);

LUT6 #(
   .INIT(64'h39d34a8b39d34a8b)  
) LUT6_inst8282 (
   .O(to_level3[506]),
   .I0(level4_in[3036]),
   .I1(level4_in[3037]),
   .I2(level4_in[3038]),
   .I3(level4_in[3039]),
   .I4(level4_in[3040]),
   .I5(level4_in[3041])
);

LUT6 #(
   .INIT(64'h154f992f154f992f)  
) LUT6_inst8283 (
   .O(to_level3[507]),
   .I0(level4_in[3042]),
   .I1(level4_in[3043]),
   .I2(level4_in[3044]),
   .I3(level4_in[3045]),
   .I4(level4_in[3046]),
   .I5(level4_in[3047])
);

LUT6 #(
   .INIT(64'hc47f8cf9c47f8cf9)  
) LUT6_inst8284 (
   .O(to_level3[508]),
   .I0(level4_in[3048]),
   .I1(level4_in[3049]),
   .I2(level4_in[3050]),
   .I3(level4_in[3051]),
   .I4(level4_in[3052]),
   .I5(level4_in[3053])
);

LUT6 #(
   .INIT(64'h6231dac56231dac5)  
) LUT6_inst8285 (
   .O(to_level3[509]),
   .I0(level4_in[3054]),
   .I1(level4_in[3055]),
   .I2(level4_in[3056]),
   .I3(level4_in[3057]),
   .I4(level4_in[3058]),
   .I5(level4_in[3059])
);

LUT6 #(
   .INIT(64'h4a10044c4a10044c)  
) LUT6_inst8286 (
   .O(to_level3[510]),
   .I0(level4_in[3060]),
   .I1(level4_in[3061]),
   .I2(level4_in[3062]),
   .I3(level4_in[3063]),
   .I4(level4_in[3064]),
   .I5(level4_in[3065])
);

LUT6 #(
   .INIT(64'h776bd2d0776bd2d0)  
) LUT6_inst8287 (
   .O(to_level3[511]),
   .I0(level4_in[3066]),
   .I1(level4_in[3067]),
   .I2(level4_in[3068]),
   .I3(level4_in[3069]),
   .I4(level4_in[3070]),
   .I5(level4_in[3071])
);

LUT6 #(
   .INIT(64'h14deff0214deff02)  
) LUT6_inst8288 (
   .O(to_level3[512]),
   .I0(level4_in[3072]),
   .I1(level4_in[3073]),
   .I2(level4_in[3074]),
   .I3(level4_in[3075]),
   .I4(level4_in[3076]),
   .I5(level4_in[3077])
);

LUT6 #(
   .INIT(64'hd39b00b4d39b00b4)  
) LUT6_inst8289 (
   .O(to_level3[513]),
   .I0(level4_in[3078]),
   .I1(level4_in[3079]),
   .I2(level4_in[3080]),
   .I3(level4_in[3081]),
   .I4(level4_in[3082]),
   .I5(level4_in[3083])
);

LUT6 #(
   .INIT(64'h8fb63bac8fb63bac)  
) LUT6_inst8290 (
   .O(to_level3[514]),
   .I0(level4_in[3084]),
   .I1(level4_in[3085]),
   .I2(level4_in[3086]),
   .I3(level4_in[3087]),
   .I4(level4_in[3088]),
   .I5(level4_in[3089])
);

LUT6 #(
   .INIT(64'h18149f4d18149f4d)  
) LUT6_inst8291 (
   .O(to_level3[515]),
   .I0(level4_in[3090]),
   .I1(level4_in[3091]),
   .I2(level4_in[3092]),
   .I3(level4_in[3093]),
   .I4(level4_in[3094]),
   .I5(level4_in[3095])
);

LUT6 #(
   .INIT(64'hf81d30f2f81d30f2)  
) LUT6_inst8292 (
   .O(to_level3[516]),
   .I0(level4_in[3096]),
   .I1(level4_in[3097]),
   .I2(level4_in[3098]),
   .I3(level4_in[3099]),
   .I4(level4_in[3100]),
   .I5(level4_in[3101])
);

LUT6 #(
   .INIT(64'hc5db8336c5db8336)  
) LUT6_inst8293 (
   .O(to_level3[517]),
   .I0(level4_in[3102]),
   .I1(level4_in[3103]),
   .I2(level4_in[3104]),
   .I3(level4_in[3105]),
   .I4(level4_in[3106]),
   .I5(level4_in[3107])
);

LUT6 #(
   .INIT(64'hd6419aa3d6419aa3)  
) LUT6_inst8294 (
   .O(to_level3[518]),
   .I0(level4_in[3108]),
   .I1(level4_in[3109]),
   .I2(level4_in[3110]),
   .I3(level4_in[3111]),
   .I4(level4_in[3112]),
   .I5(level4_in[3113])
);

LUT6 #(
   .INIT(64'hde7fde02de7fde02)  
) LUT6_inst8295 (
   .O(to_level3[519]),
   .I0(level4_in[3114]),
   .I1(level4_in[3115]),
   .I2(level4_in[3116]),
   .I3(level4_in[3117]),
   .I4(level4_in[3118]),
   .I5(level4_in[3119])
);

LUT6 #(
   .INIT(64'hd3fed42ad3fed42a)  
) LUT6_inst8296 (
   .O(to_level3[520]),
   .I0(level4_in[3120]),
   .I1(level4_in[3121]),
   .I2(level4_in[3122]),
   .I3(level4_in[3123]),
   .I4(level4_in[3124]),
   .I5(level4_in[3125])
);

LUT6 #(
   .INIT(64'h4b85b0e74b85b0e7)  
) LUT6_inst8297 (
   .O(to_level3[521]),
   .I0(level4_in[3126]),
   .I1(level4_in[3127]),
   .I2(level4_in[3128]),
   .I3(level4_in[3129]),
   .I4(level4_in[3130]),
   .I5(level4_in[3131])
);

LUT6 #(
   .INIT(64'h188ba01c188ba01c)  
) LUT6_inst8298 (
   .O(to_level3[522]),
   .I0(level4_in[3132]),
   .I1(level4_in[3133]),
   .I2(level4_in[3134]),
   .I3(level4_in[3135]),
   .I4(level4_in[3136]),
   .I5(level4_in[3137])
);

LUT6 #(
   .INIT(64'hdac08d7bdac08d7b)  
) LUT6_inst8299 (
   .O(to_level3[523]),
   .I0(level4_in[3138]),
   .I1(level4_in[3139]),
   .I2(level4_in[3140]),
   .I3(level4_in[3141]),
   .I4(level4_in[3142]),
   .I5(level4_in[3143])
);

LUT6 #(
   .INIT(64'h329211f0329211f0)  
) LUT6_inst8300 (
   .O(to_level3[524]),
   .I0(level4_in[3144]),
   .I1(level4_in[3145]),
   .I2(level4_in[3146]),
   .I3(level4_in[3147]),
   .I4(level4_in[3148]),
   .I5(level4_in[3149])
);

LUT6 #(
   .INIT(64'h81dbd82981dbd829)  
) LUT6_inst8301 (
   .O(to_level3[525]),
   .I0(level4_in[3150]),
   .I1(level4_in[3151]),
   .I2(level4_in[3152]),
   .I3(level4_in[3153]),
   .I4(level4_in[3154]),
   .I5(level4_in[3155])
);

LUT6 #(
   .INIT(64'h63ca98b863ca98b8)  
) LUT6_inst8302 (
   .O(to_level3[526]),
   .I0(level4_in[3156]),
   .I1(level4_in[3157]),
   .I2(level4_in[3158]),
   .I3(level4_in[3159]),
   .I4(level4_in[3160]),
   .I5(level4_in[3161])
);

LUT6 #(
   .INIT(64'h43c5ecfd43c5ecfd)  
) LUT6_inst8303 (
   .O(to_level3[527]),
   .I0(level4_in[3162]),
   .I1(level4_in[3163]),
   .I2(level4_in[3164]),
   .I3(level4_in[3165]),
   .I4(level4_in[3166]),
   .I5(level4_in[3167])
);

LUT6 #(
   .INIT(64'ha7641b8da7641b8d)  
) LUT6_inst8304 (
   .O(to_level3[528]),
   .I0(level4_in[3168]),
   .I1(level4_in[3169]),
   .I2(level4_in[3170]),
   .I3(level4_in[3171]),
   .I4(level4_in[3172]),
   .I5(level4_in[3173])
);

LUT6 #(
   .INIT(64'hcb298930cb298930)  
) LUT6_inst8305 (
   .O(to_level3[529]),
   .I0(level4_in[3174]),
   .I1(level4_in[3175]),
   .I2(level4_in[3176]),
   .I3(level4_in[3177]),
   .I4(level4_in[3178]),
   .I5(level4_in[3179])
);

LUT6 #(
   .INIT(64'hf0d0313af0d0313a)  
) LUT6_inst8306 (
   .O(to_level3[530]),
   .I0(level4_in[3180]),
   .I1(level4_in[3181]),
   .I2(level4_in[3182]),
   .I3(level4_in[3183]),
   .I4(level4_in[3184]),
   .I5(level4_in[3185])
);

LUT6 #(
   .INIT(64'ha9ca2bc0a9ca2bc0)  
) LUT6_inst8307 (
   .O(to_level3[531]),
   .I0(level4_in[3186]),
   .I1(level4_in[3187]),
   .I2(level4_in[3188]),
   .I3(level4_in[3189]),
   .I4(level4_in[3190]),
   .I5(level4_in[3191])
);

LUT6 #(
   .INIT(64'h1f5d5af21f5d5af2)  
) LUT6_inst8308 (
   .O(to_level3[532]),
   .I0(level4_in[3192]),
   .I1(level4_in[3193]),
   .I2(level4_in[3194]),
   .I3(level4_in[3195]),
   .I4(level4_in[3196]),
   .I5(level4_in[3197])
);

LUT6 #(
   .INIT(64'h9659355796593557)  
) LUT6_inst8309 (
   .O(to_level3[533]),
   .I0(level4_in[3198]),
   .I1(level4_in[3199]),
   .I2(level4_in[3200]),
   .I3(level4_in[3201]),
   .I4(level4_in[3202]),
   .I5(level4_in[3203])
);

LUT6 #(
   .INIT(64'h30bcda1c30bcda1c)  
) LUT6_inst8310 (
   .O(to_level3[534]),
   .I0(level4_in[3204]),
   .I1(level4_in[3205]),
   .I2(level4_in[3206]),
   .I3(level4_in[3207]),
   .I4(level4_in[3208]),
   .I5(level4_in[3209])
);

LUT6 #(
   .INIT(64'h7536fa2e7536fa2e)  
) LUT6_inst8311 (
   .O(to_level3[535]),
   .I0(level4_in[3210]),
   .I1(level4_in[3211]),
   .I2(level4_in[3212]),
   .I3(level4_in[3213]),
   .I4(level4_in[3214]),
   .I5(level4_in[3215])
);

LUT6 #(
   .INIT(64'h70b2234070b22340)  
) LUT6_inst8312 (
   .O(to_level3[536]),
   .I0(level4_in[3216]),
   .I1(level4_in[3217]),
   .I2(level4_in[3218]),
   .I3(level4_in[3219]),
   .I4(level4_in[3220]),
   .I5(level4_in[3221])
);

LUT6 #(
   .INIT(64'h87b2fb9c87b2fb9c)  
) LUT6_inst8313 (
   .O(to_level3[537]),
   .I0(level4_in[3222]),
   .I1(level4_in[3223]),
   .I2(level4_in[3224]),
   .I3(level4_in[3225]),
   .I4(level4_in[3226]),
   .I5(level4_in[3227])
);

LUT6 #(
   .INIT(64'haceac1dbaceac1db)  
) LUT6_inst8314 (
   .O(to_level3[538]),
   .I0(level4_in[3228]),
   .I1(level4_in[3229]),
   .I2(level4_in[3230]),
   .I3(level4_in[3231]),
   .I4(level4_in[3232]),
   .I5(level4_in[3233])
);

LUT6 #(
   .INIT(64'h792fdb19792fdb19)  
) LUT6_inst8315 (
   .O(to_level3[539]),
   .I0(level4_in[3234]),
   .I1(level4_in[3235]),
   .I2(level4_in[3236]),
   .I3(level4_in[3237]),
   .I4(level4_in[3238]),
   .I5(level4_in[3239])
);

LUT6 #(
   .INIT(64'he7357e7fe7357e7f)  
) LUT6_inst8316 (
   .O(to_level3[540]),
   .I0(level4_in[3240]),
   .I1(level4_in[3241]),
   .I2(level4_in[3242]),
   .I3(level4_in[3243]),
   .I4(level4_in[3244]),
   .I5(level4_in[3245])
);

LUT6 #(
   .INIT(64'h8c069e128c069e12)  
) LUT6_inst8317 (
   .O(to_level3[541]),
   .I0(level4_in[3246]),
   .I1(level4_in[3247]),
   .I2(level4_in[3248]),
   .I3(level4_in[3249]),
   .I4(level4_in[3250]),
   .I5(level4_in[3251])
);

LUT6 #(
   .INIT(64'h166295da166295da)  
) LUT6_inst8318 (
   .O(to_level3[542]),
   .I0(level4_in[3252]),
   .I1(level4_in[3253]),
   .I2(level4_in[3254]),
   .I3(level4_in[3255]),
   .I4(level4_in[3256]),
   .I5(level4_in[3257])
);

LUT6 #(
   .INIT(64'h8ff5bf868ff5bf86)  
) LUT6_inst8319 (
   .O(to_level3[543]),
   .I0(level4_in[3258]),
   .I1(level4_in[3259]),
   .I2(level4_in[3260]),
   .I3(level4_in[3261]),
   .I4(level4_in[3262]),
   .I5(level4_in[3263])
);

LUT6 #(
   .INIT(64'hb905e34db905e34d)  
) LUT6_inst8320 (
   .O(to_level3[544]),
   .I0(level4_in[3264]),
   .I1(level4_in[3265]),
   .I2(level4_in[3266]),
   .I3(level4_in[3267]),
   .I4(level4_in[3268]),
   .I5(level4_in[3269])
);

LUT6 #(
   .INIT(64'h6a455ebf6a455ebf)  
) LUT6_inst8321 (
   .O(to_level3[545]),
   .I0(level4_in[3270]),
   .I1(level4_in[3271]),
   .I2(level4_in[3272]),
   .I3(level4_in[3273]),
   .I4(level4_in[3274]),
   .I5(level4_in[3275])
);

LUT6 #(
   .INIT(64'h5787d65e5787d65e)  
) LUT6_inst8322 (
   .O(to_level3[546]),
   .I0(level4_in[3276]),
   .I1(level4_in[3277]),
   .I2(level4_in[3278]),
   .I3(level4_in[3279]),
   .I4(level4_in[3280]),
   .I5(level4_in[3281])
);

LUT6 #(
   .INIT(64'hb877587eb877587e)  
) LUT6_inst8323 (
   .O(to_level3[547]),
   .I0(level4_in[3282]),
   .I1(level4_in[3283]),
   .I2(level4_in[3284]),
   .I3(level4_in[3285]),
   .I4(level4_in[3286]),
   .I5(level4_in[3287])
);

LUT6 #(
   .INIT(64'h568bb889568bb889)  
) LUT6_inst8324 (
   .O(to_level3[548]),
   .I0(level4_in[3288]),
   .I1(level4_in[3289]),
   .I2(level4_in[3290]),
   .I3(level4_in[3291]),
   .I4(level4_in[3292]),
   .I5(level4_in[3293])
);

LUT6 #(
   .INIT(64'h41fb5e4141fb5e41)  
) LUT6_inst8325 (
   .O(to_level3[549]),
   .I0(level4_in[3294]),
   .I1(level4_in[3295]),
   .I2(level4_in[3296]),
   .I3(level4_in[3297]),
   .I4(level4_in[3298]),
   .I5(level4_in[3299])
);

LUT6 #(
   .INIT(64'h74fb959274fb9592)  
) LUT6_inst8326 (
   .O(to_level3[550]),
   .I0(level4_in[3300]),
   .I1(level4_in[3301]),
   .I2(level4_in[3302]),
   .I3(level4_in[3303]),
   .I4(level4_in[3304]),
   .I5(level4_in[3305])
);

LUT6 #(
   .INIT(64'h21ed179021ed1790)  
) LUT6_inst8327 (
   .O(to_level3[551]),
   .I0(level4_in[3306]),
   .I1(level4_in[3307]),
   .I2(level4_in[3308]),
   .I3(level4_in[3309]),
   .I4(level4_in[3310]),
   .I5(level4_in[3311])
);

LUT6 #(
   .INIT(64'h64d0b8b964d0b8b9)  
) LUT6_inst8328 (
   .O(to_level3[552]),
   .I0(level4_in[3312]),
   .I1(level4_in[3313]),
   .I2(level4_in[3314]),
   .I3(level4_in[3315]),
   .I4(level4_in[3316]),
   .I5(level4_in[3317])
);

LUT6 #(
   .INIT(64'h872f4187872f4187)  
) LUT6_inst8329 (
   .O(to_level3[553]),
   .I0(level4_in[3318]),
   .I1(level4_in[3319]),
   .I2(level4_in[3320]),
   .I3(level4_in[3321]),
   .I4(level4_in[3322]),
   .I5(level4_in[3323])
);

LUT6 #(
   .INIT(64'h87dc73a787dc73a7)  
) LUT6_inst8330 (
   .O(to_level3[554]),
   .I0(level4_in[3324]),
   .I1(level4_in[3325]),
   .I2(level4_in[3326]),
   .I3(level4_in[3327]),
   .I4(level4_in[3328]),
   .I5(level4_in[3329])
);

LUT6 #(
   .INIT(64'h3bcff19f3bcff19f)  
) LUT6_inst8331 (
   .O(to_level3[555]),
   .I0(level4_in[3330]),
   .I1(level4_in[3331]),
   .I2(level4_in[3332]),
   .I3(level4_in[3333]),
   .I4(level4_in[3334]),
   .I5(level4_in[3335])
);

LUT6 #(
   .INIT(64'ha4268b87a4268b87)  
) LUT6_inst8332 (
   .O(to_level3[556]),
   .I0(level4_in[3336]),
   .I1(level4_in[3337]),
   .I2(level4_in[3338]),
   .I3(level4_in[3339]),
   .I4(level4_in[3340]),
   .I5(level4_in[3341])
);

LUT6 #(
   .INIT(64'h8cf67a278cf67a27)  
) LUT6_inst8333 (
   .O(to_level3[557]),
   .I0(level4_in[3342]),
   .I1(level4_in[3343]),
   .I2(level4_in[3344]),
   .I3(level4_in[3345]),
   .I4(level4_in[3346]),
   .I5(level4_in[3347])
);

LUT6 #(
   .INIT(64'h04b3f08004b3f080)  
) LUT6_inst8334 (
   .O(to_level3[558]),
   .I0(level4_in[3348]),
   .I1(level4_in[3349]),
   .I2(level4_in[3350]),
   .I3(level4_in[3351]),
   .I4(level4_in[3352]),
   .I5(level4_in[3353])
);

LUT6 #(
   .INIT(64'h6420a9206420a920)  
) LUT6_inst8335 (
   .O(to_level3[559]),
   .I0(level4_in[3354]),
   .I1(level4_in[3355]),
   .I2(level4_in[3356]),
   .I3(level4_in[3357]),
   .I4(level4_in[3358]),
   .I5(level4_in[3359])
);

LUT6 #(
   .INIT(64'hfc4e6a60fc4e6a60)  
) LUT6_inst8336 (
   .O(to_level3[560]),
   .I0(level4_in[3360]),
   .I1(level4_in[3361]),
   .I2(level4_in[3362]),
   .I3(level4_in[3363]),
   .I4(level4_in[3364]),
   .I5(level4_in[3365])
);

LUT6 #(
   .INIT(64'hc833fdb9c833fdb9)  
) LUT6_inst8337 (
   .O(to_level3[561]),
   .I0(level4_in[3366]),
   .I1(level4_in[3367]),
   .I2(level4_in[3368]),
   .I3(level4_in[3369]),
   .I4(level4_in[3370]),
   .I5(level4_in[3371])
);

LUT6 #(
   .INIT(64'h66961f1666961f16)  
) LUT6_inst8338 (
   .O(to_level3[562]),
   .I0(level4_in[3372]),
   .I1(level4_in[3373]),
   .I2(level4_in[3374]),
   .I3(level4_in[3375]),
   .I4(level4_in[3376]),
   .I5(level4_in[3377])
);

LUT6 #(
   .INIT(64'h6f8f82b16f8f82b1)  
) LUT6_inst8339 (
   .O(to_level3[563]),
   .I0(level4_in[3378]),
   .I1(level4_in[3379]),
   .I2(level4_in[3380]),
   .I3(level4_in[3381]),
   .I4(level4_in[3382]),
   .I5(level4_in[3383])
);

LUT6 #(
   .INIT(64'h6d6420996d642099)  
) LUT6_inst8340 (
   .O(to_level3[564]),
   .I0(level4_in[3384]),
   .I1(level4_in[3385]),
   .I2(level4_in[3386]),
   .I3(level4_in[3387]),
   .I4(level4_in[3388]),
   .I5(level4_in[3389])
);

LUT6 #(
   .INIT(64'h2d126dab2d126dab)  
) LUT6_inst8341 (
   .O(to_level3[565]),
   .I0(level4_in[3390]),
   .I1(level4_in[3391]),
   .I2(level4_in[3392]),
   .I3(level4_in[3393]),
   .I4(level4_in[3394]),
   .I5(level4_in[3395])
);

LUT6 #(
   .INIT(64'h34c9823534c98235)  
) LUT6_inst8342 (
   .O(to_level3[566]),
   .I0(level4_in[3396]),
   .I1(level4_in[3397]),
   .I2(level4_in[3398]),
   .I3(level4_in[3399]),
   .I4(level4_in[3400]),
   .I5(level4_in[3401])
);

LUT6 #(
   .INIT(64'h0aa882b10aa882b1)  
) LUT6_inst8343 (
   .O(to_level3[567]),
   .I0(level4_in[3402]),
   .I1(level4_in[3403]),
   .I2(level4_in[3404]),
   .I3(level4_in[3405]),
   .I4(level4_in[3406]),
   .I5(level4_in[3407])
);

LUT6 #(
   .INIT(64'h4103577641035776)  
) LUT6_inst8344 (
   .O(to_level3[568]),
   .I0(level4_in[3408]),
   .I1(level4_in[3409]),
   .I2(level4_in[3410]),
   .I3(level4_in[3411]),
   .I4(level4_in[3412]),
   .I5(level4_in[3413])
);

LUT6 #(
   .INIT(64'h620e1040620e1040)  
) LUT6_inst8345 (
   .O(to_level3[569]),
   .I0(level4_in[3414]),
   .I1(level4_in[3415]),
   .I2(level4_in[3416]),
   .I3(level4_in[3417]),
   .I4(level4_in[3418]),
   .I5(level4_in[3419])
);

LUT6 #(
   .INIT(64'h6a0bbb9f6a0bbb9f)  
) LUT6_inst8346 (
   .O(to_level3[570]),
   .I0(level4_in[3420]),
   .I1(level4_in[3421]),
   .I2(level4_in[3422]),
   .I3(level4_in[3423]),
   .I4(level4_in[3424]),
   .I5(level4_in[3425])
);

LUT6 #(
   .INIT(64'h2ad45c842ad45c84)  
) LUT6_inst8347 (
   .O(to_level3[571]),
   .I0(level4_in[3426]),
   .I1(level4_in[3427]),
   .I2(level4_in[3428]),
   .I3(level4_in[3429]),
   .I4(level4_in[3430]),
   .I5(level4_in[3431])
);

LUT6 #(
   .INIT(64'hfa2e2b36fa2e2b36)  
) LUT6_inst8348 (
   .O(to_level3[572]),
   .I0(level4_in[3432]),
   .I1(level4_in[3433]),
   .I2(level4_in[3434]),
   .I3(level4_in[3435]),
   .I4(level4_in[3436]),
   .I5(level4_in[3437])
);

LUT6 #(
   .INIT(64'haafefaefaafefaef)  
) LUT6_inst8349 (
   .O(to_level3[573]),
   .I0(level4_in[3438]),
   .I1(level4_in[3439]),
   .I2(level4_in[3440]),
   .I3(level4_in[3441]),
   .I4(level4_in[3442]),
   .I5(level4_in[3443])
);

LUT6 #(
   .INIT(64'hde888fdbde888fdb)  
) LUT6_inst8350 (
   .O(to_level3[574]),
   .I0(level4_in[3444]),
   .I1(level4_in[3445]),
   .I2(level4_in[3446]),
   .I3(level4_in[3447]),
   .I4(level4_in[3448]),
   .I5(level4_in[3449])
);

LUT6 #(
   .INIT(64'h0ca737440ca73744)  
) LUT6_inst8351 (
   .O(to_level3[575]),
   .I0(level4_in[3450]),
   .I1(level4_in[3451]),
   .I2(level4_in[3452]),
   .I3(level4_in[3453]),
   .I4(level4_in[3454]),
   .I5(level4_in[3455])
);

LUT6 #(
   .INIT(64'he01a66c7e01a66c7)  
) LUT6_inst8352 (
   .O(to_level3[576]),
   .I0(level4_in[3456]),
   .I1(level4_in[3457]),
   .I2(level4_in[3458]),
   .I3(level4_in[3459]),
   .I4(level4_in[3460]),
   .I5(level4_in[3461])
);

LUT6 #(
   .INIT(64'h2055c2c32055c2c3)  
) LUT6_inst8353 (
   .O(to_level3[577]),
   .I0(level4_in[3462]),
   .I1(level4_in[3463]),
   .I2(level4_in[3464]),
   .I3(level4_in[3465]),
   .I4(level4_in[3466]),
   .I5(level4_in[3467])
);

LUT6 #(
   .INIT(64'hbed8c072bed8c072)  
) LUT6_inst8354 (
   .O(to_level3[578]),
   .I0(level4_in[3468]),
   .I1(level4_in[3469]),
   .I2(level4_in[3470]),
   .I3(level4_in[3471]),
   .I4(level4_in[3472]),
   .I5(level4_in[3473])
);

LUT6 #(
   .INIT(64'he824282fe824282f)  
) LUT6_inst8355 (
   .O(to_level3[579]),
   .I0(level4_in[3474]),
   .I1(level4_in[3475]),
   .I2(level4_in[3476]),
   .I3(level4_in[3477]),
   .I4(level4_in[3478]),
   .I5(level4_in[3479])
);

LUT6 #(
   .INIT(64'he6b3964fe6b3964f)  
) LUT6_inst8356 (
   .O(to_level3[580]),
   .I0(level4_in[3480]),
   .I1(level4_in[3481]),
   .I2(level4_in[3482]),
   .I3(level4_in[3483]),
   .I4(level4_in[3484]),
   .I5(level4_in[3485])
);

LUT6 #(
   .INIT(64'h34d3bdec34d3bdec)  
) LUT6_inst8357 (
   .O(to_level3[581]),
   .I0(level4_in[3486]),
   .I1(level4_in[3487]),
   .I2(level4_in[3488]),
   .I3(level4_in[3489]),
   .I4(level4_in[3490]),
   .I5(level4_in[3491])
);

LUT6 #(
   .INIT(64'h31f0b4f431f0b4f4)  
) LUT6_inst8358 (
   .O(to_level3[582]),
   .I0(level4_in[3492]),
   .I1(level4_in[3493]),
   .I2(level4_in[3494]),
   .I3(level4_in[3495]),
   .I4(level4_in[3496]),
   .I5(level4_in[3497])
);

LUT6 #(
   .INIT(64'h2bd9b6362bd9b636)  
) LUT6_inst8359 (
   .O(to_level3[583]),
   .I0(level4_in[3498]),
   .I1(level4_in[3499]),
   .I2(level4_in[3500]),
   .I3(level4_in[3501]),
   .I4(level4_in[3502]),
   .I5(level4_in[3503])
);

LUT6 #(
   .INIT(64'hc916f696c916f696)  
) LUT6_inst8360 (
   .O(to_level3[584]),
   .I0(level4_in[3504]),
   .I1(level4_in[3505]),
   .I2(level4_in[3506]),
   .I3(level4_in[3507]),
   .I4(level4_in[3508]),
   .I5(level4_in[3509])
);

LUT6 #(
   .INIT(64'h43a4b34e43a4b34e)  
) LUT6_inst8361 (
   .O(to_level3[585]),
   .I0(level4_in[3510]),
   .I1(level4_in[3511]),
   .I2(level4_in[3512]),
   .I3(level4_in[3513]),
   .I4(level4_in[3514]),
   .I5(level4_in[3515])
);

LUT6 #(
   .INIT(64'he6335fa3e6335fa3)  
) LUT6_inst8362 (
   .O(to_level3[586]),
   .I0(level4_in[3516]),
   .I1(level4_in[3517]),
   .I2(level4_in[3518]),
   .I3(level4_in[3519]),
   .I4(level4_in[3520]),
   .I5(level4_in[3521])
);

LUT6 #(
   .INIT(64'h7e9049507e904950)  
) LUT6_inst8363 (
   .O(to_level3[587]),
   .I0(level4_in[3522]),
   .I1(level4_in[3523]),
   .I2(level4_in[3524]),
   .I3(level4_in[3525]),
   .I4(level4_in[3526]),
   .I5(level4_in[3527])
);

LUT6 #(
   .INIT(64'h8afa346b8afa346b)  
) LUT6_inst8364 (
   .O(to_level3[588]),
   .I0(level4_in[3528]),
   .I1(level4_in[3529]),
   .I2(level4_in[3530]),
   .I3(level4_in[3531]),
   .I4(level4_in[3532]),
   .I5(level4_in[3533])
);

LUT6 #(
   .INIT(64'h21516bd221516bd2)  
) LUT6_inst8365 (
   .O(to_level3[589]),
   .I0(level4_in[3534]),
   .I1(level4_in[3535]),
   .I2(level4_in[3536]),
   .I3(level4_in[3537]),
   .I4(level4_in[3538]),
   .I5(level4_in[3539])
);

LUT6 #(
   .INIT(64'h368c46c9368c46c9)  
) LUT6_inst8366 (
   .O(to_level3[590]),
   .I0(level4_in[3540]),
   .I1(level4_in[3541]),
   .I2(level4_in[3542]),
   .I3(level4_in[3543]),
   .I4(level4_in[3544]),
   .I5(level4_in[3545])
);

LUT6 #(
   .INIT(64'h80afa66980afa669)  
) LUT6_inst8367 (
   .O(to_level3[591]),
   .I0(level4_in[3546]),
   .I1(level4_in[3547]),
   .I2(level4_in[3548]),
   .I3(level4_in[3549]),
   .I4(level4_in[3550]),
   .I5(level4_in[3551])
);

LUT6 #(
   .INIT(64'h4723dd804723dd80)  
) LUT6_inst8368 (
   .O(to_level3[592]),
   .I0(level4_in[3552]),
   .I1(level4_in[3553]),
   .I2(level4_in[3554]),
   .I3(level4_in[3555]),
   .I4(level4_in[3556]),
   .I5(level4_in[3557])
);

LUT6 #(
   .INIT(64'h99df1b5699df1b56)  
) LUT6_inst8369 (
   .O(to_level3[593]),
   .I0(level4_in[3558]),
   .I1(level4_in[3559]),
   .I2(level4_in[3560]),
   .I3(level4_in[3561]),
   .I4(level4_in[3562]),
   .I5(level4_in[3563])
);

LUT6 #(
   .INIT(64'hfff8df82fff8df82)  
) LUT6_inst8370 (
   .O(to_level3[594]),
   .I0(level4_in[3564]),
   .I1(level4_in[3565]),
   .I2(level4_in[3566]),
   .I3(level4_in[3567]),
   .I4(level4_in[3568]),
   .I5(level4_in[3569])
);

LUT6 #(
   .INIT(64'h4aac873f4aac873f)  
) LUT6_inst8371 (
   .O(to_level3[595]),
   .I0(level4_in[3570]),
   .I1(level4_in[3571]),
   .I2(level4_in[3572]),
   .I3(level4_in[3573]),
   .I4(level4_in[3574]),
   .I5(level4_in[3575])
);

LUT6 #(
   .INIT(64'h7332ff9b7332ff9b)  
) LUT6_inst8372 (
   .O(to_level3[596]),
   .I0(level4_in[3576]),
   .I1(level4_in[3577]),
   .I2(level4_in[3578]),
   .I3(level4_in[3579]),
   .I4(level4_in[3580]),
   .I5(level4_in[3581])
);

LUT6 #(
   .INIT(64'ha091ad8ba091ad8b)  
) LUT6_inst8373 (
   .O(to_level3[597]),
   .I0(level4_in[3582]),
   .I1(level4_in[3583]),
   .I2(level4_in[3584]),
   .I3(level4_in[3585]),
   .I4(level4_in[3586]),
   .I5(level4_in[3587])
);

LUT6 #(
   .INIT(64'h1c3df2ed1c3df2ed)  
) LUT6_inst8374 (
   .O(to_level3[598]),
   .I0(level4_in[3588]),
   .I1(level4_in[3589]),
   .I2(level4_in[3590]),
   .I3(level4_in[3591]),
   .I4(level4_in[3592]),
   .I5(level4_in[3593])
);

LUT6 #(
   .INIT(64'hcdb51368cdb51368)  
) LUT6_inst8375 (
   .O(to_level3[599]),
   .I0(level4_in[3594]),
   .I1(level4_in[3595]),
   .I2(level4_in[3596]),
   .I3(level4_in[3597]),
   .I4(level4_in[3598]),
   .I5(level4_in[3599])
);

LUT6 #(
   .INIT(64'h7bd56a087bd56a08)  
) LUT6_inst8376 (
   .O(to_level3[600]),
   .I0(level4_in[3600]),
   .I1(level4_in[3601]),
   .I2(level4_in[3602]),
   .I3(level4_in[3603]),
   .I4(level4_in[3604]),
   .I5(level4_in[3605])
);

LUT6 #(
   .INIT(64'h5343990853439908)  
) LUT6_inst8377 (
   .O(to_level3[601]),
   .I0(level4_in[3606]),
   .I1(level4_in[3607]),
   .I2(level4_in[3608]),
   .I3(level4_in[3609]),
   .I4(level4_in[3610]),
   .I5(level4_in[3611])
);

LUT6 #(
   .INIT(64'h9d4e33e29d4e33e2)  
) LUT6_inst8378 (
   .O(to_level3[602]),
   .I0(level4_in[3612]),
   .I1(level4_in[3613]),
   .I2(level4_in[3614]),
   .I3(level4_in[3615]),
   .I4(level4_in[3616]),
   .I5(level4_in[3617])
);

LUT6 #(
   .INIT(64'h4167349b4167349b)  
) LUT6_inst8379 (
   .O(to_level3[603]),
   .I0(level4_in[3618]),
   .I1(level4_in[3619]),
   .I2(level4_in[3620]),
   .I3(level4_in[3621]),
   .I4(level4_in[3622]),
   .I5(level4_in[3623])
);

LUT6 #(
   .INIT(64'hf6549b46f6549b46)  
) LUT6_inst8380 (
   .O(to_level3[604]),
   .I0(level4_in[3624]),
   .I1(level4_in[3625]),
   .I2(level4_in[3626]),
   .I3(level4_in[3627]),
   .I4(level4_in[3628]),
   .I5(level4_in[3629])
);

LUT6 #(
   .INIT(64'h1832396718323967)  
) LUT6_inst8381 (
   .O(to_level3[605]),
   .I0(level4_in[3630]),
   .I1(level4_in[3631]),
   .I2(level4_in[3632]),
   .I3(level4_in[3633]),
   .I4(level4_in[3634]),
   .I5(level4_in[3635])
);

LUT6 #(
   .INIT(64'hbc8cfb6abc8cfb6a)  
) LUT6_inst8382 (
   .O(to_level3[606]),
   .I0(level4_in[3636]),
   .I1(level4_in[3637]),
   .I2(level4_in[3638]),
   .I3(level4_in[3639]),
   .I4(level4_in[3640]),
   .I5(level4_in[3641])
);

LUT6 #(
   .INIT(64'h197b7425197b7425)  
) LUT6_inst8383 (
   .O(to_level3[607]),
   .I0(level4_in[3642]),
   .I1(level4_in[3643]),
   .I2(level4_in[3644]),
   .I3(level4_in[3645]),
   .I4(level4_in[3646]),
   .I5(level4_in[3647])
);

LUT6 #(
   .INIT(64'hb14683aab14683aa)  
) LUT6_inst8384 (
   .O(to_level3[608]),
   .I0(level4_in[3648]),
   .I1(level4_in[3649]),
   .I2(level4_in[3650]),
   .I3(level4_in[3651]),
   .I4(level4_in[3652]),
   .I5(level4_in[3653])
);

LUT6 #(
   .INIT(64'h4ef565f94ef565f9)  
) LUT6_inst8385 (
   .O(to_level3[609]),
   .I0(level4_in[3654]),
   .I1(level4_in[3655]),
   .I2(level4_in[3656]),
   .I3(level4_in[3657]),
   .I4(level4_in[3658]),
   .I5(level4_in[3659])
);

LUT6 #(
   .INIT(64'hccd21234ccd21234)  
) LUT6_inst8386 (
   .O(to_level3[610]),
   .I0(level4_in[3660]),
   .I1(level4_in[3661]),
   .I2(level4_in[3662]),
   .I3(level4_in[3663]),
   .I4(level4_in[3664]),
   .I5(level4_in[3665])
);

LUT6 #(
   .INIT(64'hc0481b8ac0481b8a)  
) LUT6_inst8387 (
   .O(to_level3[611]),
   .I0(level4_in[3666]),
   .I1(level4_in[3667]),
   .I2(level4_in[3668]),
   .I3(level4_in[3669]),
   .I4(level4_in[3670]),
   .I5(level4_in[3671])
);

LUT6 #(
   .INIT(64'hb3ad127db3ad127d)  
) LUT6_inst8388 (
   .O(to_level3[612]),
   .I0(level4_in[3672]),
   .I1(level4_in[3673]),
   .I2(level4_in[3674]),
   .I3(level4_in[3675]),
   .I4(level4_in[3676]),
   .I5(level4_in[3677])
);

LUT6 #(
   .INIT(64'h998e9920998e9920)  
) LUT6_inst8389 (
   .O(to_level3[613]),
   .I0(level4_in[3678]),
   .I1(level4_in[3679]),
   .I2(level4_in[3680]),
   .I3(level4_in[3681]),
   .I4(level4_in[3682]),
   .I5(level4_in[3683])
);

LUT6 #(
   .INIT(64'h676a10f1676a10f1)  
) LUT6_inst8390 (
   .O(to_level3[614]),
   .I0(level4_in[3684]),
   .I1(level4_in[3685]),
   .I2(level4_in[3686]),
   .I3(level4_in[3687]),
   .I4(level4_in[3688]),
   .I5(level4_in[3689])
);

LUT6 #(
   .INIT(64'h089ee5fd089ee5fd)  
) LUT6_inst8391 (
   .O(to_level3[615]),
   .I0(level4_in[3690]),
   .I1(level4_in[3691]),
   .I2(level4_in[3692]),
   .I3(level4_in[3693]),
   .I4(level4_in[3694]),
   .I5(level4_in[3695])
);

LUT6 #(
   .INIT(64'h0bfaa8cb0bfaa8cb)  
) LUT6_inst8392 (
   .O(to_level3[616]),
   .I0(level4_in[3696]),
   .I1(level4_in[3697]),
   .I2(level4_in[3698]),
   .I3(level4_in[3699]),
   .I4(level4_in[3700]),
   .I5(level4_in[3701])
);

LUT6 #(
   .INIT(64'hbb4f2f25bb4f2f25)  
) LUT6_inst8393 (
   .O(to_level3[617]),
   .I0(level4_in[3702]),
   .I1(level4_in[3703]),
   .I2(level4_in[3704]),
   .I3(level4_in[3705]),
   .I4(level4_in[3706]),
   .I5(level4_in[3707])
);

LUT6 #(
   .INIT(64'h30e95d5b30e95d5b)  
) LUT6_inst8394 (
   .O(to_level3[618]),
   .I0(level4_in[3708]),
   .I1(level4_in[3709]),
   .I2(level4_in[3710]),
   .I3(level4_in[3711]),
   .I4(level4_in[3712]),
   .I5(level4_in[3713])
);

LUT6 #(
   .INIT(64'hbc6c8dcabc6c8dca)  
) LUT6_inst8395 (
   .O(to_level3[619]),
   .I0(level4_in[3714]),
   .I1(level4_in[3715]),
   .I2(level4_in[3716]),
   .I3(level4_in[3717]),
   .I4(level4_in[3718]),
   .I5(level4_in[3719])
);

LUT6 #(
   .INIT(64'hff1736b7ff1736b7)  
) LUT6_inst8396 (
   .O(to_level3[620]),
   .I0(level4_in[3720]),
   .I1(level4_in[3721]),
   .I2(level4_in[3722]),
   .I3(level4_in[3723]),
   .I4(level4_in[3724]),
   .I5(level4_in[3725])
);

LUT6 #(
   .INIT(64'h9a05c2269a05c226)  
) LUT6_inst8397 (
   .O(to_level3[621]),
   .I0(level4_in[3726]),
   .I1(level4_in[3727]),
   .I2(level4_in[3728]),
   .I3(level4_in[3729]),
   .I4(level4_in[3730]),
   .I5(level4_in[3731])
);

LUT6 #(
   .INIT(64'h034194bd034194bd)  
) LUT6_inst8398 (
   .O(to_level3[622]),
   .I0(level4_in[3732]),
   .I1(level4_in[3733]),
   .I2(level4_in[3734]),
   .I3(level4_in[3735]),
   .I4(level4_in[3736]),
   .I5(level4_in[3737])
);

LUT6 #(
   .INIT(64'hc15efde1c15efde1)  
) LUT6_inst8399 (
   .O(to_level3[623]),
   .I0(level4_in[3738]),
   .I1(level4_in[3739]),
   .I2(level4_in[3740]),
   .I3(level4_in[3741]),
   .I4(level4_in[3742]),
   .I5(level4_in[3743])
);

LUT6 #(
   .INIT(64'hd22d7e26d22d7e26)  
) LUT6_inst8400 (
   .O(to_level3[624]),
   .I0(level4_in[3744]),
   .I1(level4_in[3745]),
   .I2(level4_in[3746]),
   .I3(level4_in[3747]),
   .I4(level4_in[3748]),
   .I5(level4_in[3749])
);

LUT6 #(
   .INIT(64'h57080e2257080e22)  
) LUT6_inst8401 (
   .O(to_level3[625]),
   .I0(level4_in[3750]),
   .I1(level4_in[3751]),
   .I2(level4_in[3752]),
   .I3(level4_in[3753]),
   .I4(level4_in[3754]),
   .I5(level4_in[3755])
);

LUT6 #(
   .INIT(64'hd5217d97d5217d97)  
) LUT6_inst8402 (
   .O(to_level3[626]),
   .I0(level4_in[3756]),
   .I1(level4_in[3757]),
   .I2(level4_in[3758]),
   .I3(level4_in[3759]),
   .I4(level4_in[3760]),
   .I5(level4_in[3761])
);

LUT6 #(
   .INIT(64'h634b3385634b3385)  
) LUT6_inst8403 (
   .O(to_level3[627]),
   .I0(level4_in[3762]),
   .I1(level4_in[3763]),
   .I2(level4_in[3764]),
   .I3(level4_in[3765]),
   .I4(level4_in[3766]),
   .I5(level4_in[3767])
);

LUT6 #(
   .INIT(64'h59d0e2f359d0e2f3)  
) LUT6_inst8404 (
   .O(to_level3[628]),
   .I0(level4_in[3768]),
   .I1(level4_in[3769]),
   .I2(level4_in[3770]),
   .I3(level4_in[3771]),
   .I4(level4_in[3772]),
   .I5(level4_in[3773])
);

LUT6 #(
   .INIT(64'h3aff0f323aff0f32)  
) LUT6_inst8405 (
   .O(to_level3[629]),
   .I0(level4_in[3774]),
   .I1(level4_in[3775]),
   .I2(level4_in[3776]),
   .I3(level4_in[3777]),
   .I4(level4_in[3778]),
   .I5(level4_in[3779])
);

LUT6 #(
   .INIT(64'hd233244fd233244f)  
) LUT6_inst8406 (
   .O(to_level3[630]),
   .I0(level4_in[3780]),
   .I1(level4_in[3781]),
   .I2(level4_in[3782]),
   .I3(level4_in[3783]),
   .I4(level4_in[3784]),
   .I5(level4_in[3785])
);

LUT6 #(
   .INIT(64'hf697ba6df697ba6d)  
) LUT6_inst8407 (
   .O(to_level3[631]),
   .I0(level4_in[3786]),
   .I1(level4_in[3787]),
   .I2(level4_in[3788]),
   .I3(level4_in[3789]),
   .I4(level4_in[3790]),
   .I5(level4_in[3791])
);

LUT6 #(
   .INIT(64'h284285ff284285ff)  
) LUT6_inst8408 (
   .O(to_level3[632]),
   .I0(level4_in[3792]),
   .I1(level4_in[3793]),
   .I2(level4_in[3794]),
   .I3(level4_in[3795]),
   .I4(level4_in[3796]),
   .I5(level4_in[3797])
);

LUT6 #(
   .INIT(64'h84cba21d84cba21d)  
) LUT6_inst8409 (
   .O(to_level3[633]),
   .I0(level4_in[3798]),
   .I1(level4_in[3799]),
   .I2(level4_in[3800]),
   .I3(level4_in[3801]),
   .I4(level4_in[3802]),
   .I5(level4_in[3803])
);

LUT6 #(
   .INIT(64'h50cf73ee50cf73ee)  
) LUT6_inst8410 (
   .O(to_level3[634]),
   .I0(level4_in[3804]),
   .I1(level4_in[3805]),
   .I2(level4_in[3806]),
   .I3(level4_in[3807]),
   .I4(level4_in[3808]),
   .I5(level4_in[3809])
);

LUT6 #(
   .INIT(64'he9f39f67e9f39f67)  
) LUT6_inst8411 (
   .O(to_level3[635]),
   .I0(level4_in[3810]),
   .I1(level4_in[3811]),
   .I2(level4_in[3812]),
   .I3(level4_in[3813]),
   .I4(level4_in[3814]),
   .I5(level4_in[3815])
);

LUT6 #(
   .INIT(64'h17efeacb17efeacb)  
) LUT6_inst8412 (
   .O(to_level3[636]),
   .I0(level4_in[3816]),
   .I1(level4_in[3817]),
   .I2(level4_in[3818]),
   .I3(level4_in[3819]),
   .I4(level4_in[3820]),
   .I5(level4_in[3821])
);

LUT6 #(
   .INIT(64'hdfed6494dfed6494)  
) LUT6_inst8413 (
   .O(to_level3[637]),
   .I0(level4_in[3822]),
   .I1(level4_in[3823]),
   .I2(level4_in[3824]),
   .I3(level4_in[3825]),
   .I4(level4_in[3826]),
   .I5(level4_in[3827])
);

LUT6 #(
   .INIT(64'hcc9805b1cc9805b1)  
) LUT6_inst8414 (
   .O(to_level3[638]),
   .I0(level4_in[3828]),
   .I1(level4_in[3829]),
   .I2(level4_in[3830]),
   .I3(level4_in[3831]),
   .I4(level4_in[3832]),
   .I5(level4_in[3833])
);

LUT6 #(
   .INIT(64'hc19ba043c19ba043)  
) LUT6_inst8415 (
   .O(to_level3[639]),
   .I0(level4_in[3834]),
   .I1(level4_in[3835]),
   .I2(level4_in[3836]),
   .I3(level4_in[3837]),
   .I4(level4_in[3838]),
   .I5(level4_in[3839])
);

LUT6 #(
   .INIT(64'h589483f1589483f1)  
) LUT6_inst8416 (
   .O(to_level3[640]),
   .I0(level4_in[3840]),
   .I1(level4_in[3841]),
   .I2(level4_in[3842]),
   .I3(level4_in[3843]),
   .I4(level4_in[3844]),
   .I5(level4_in[3845])
);

LUT6 #(
   .INIT(64'hee4e537bee4e537b)  
) LUT6_inst8417 (
   .O(to_level3[641]),
   .I0(level4_in[3846]),
   .I1(level4_in[3847]),
   .I2(level4_in[3848]),
   .I3(level4_in[3849]),
   .I4(level4_in[3850]),
   .I5(level4_in[3851])
);

LUT6 #(
   .INIT(64'hbca0e6bcbca0e6bc)  
) LUT6_inst8418 (
   .O(to_level3[642]),
   .I0(level4_in[3852]),
   .I1(level4_in[3853]),
   .I2(level4_in[3854]),
   .I3(level4_in[3855]),
   .I4(level4_in[3856]),
   .I5(level4_in[3857])
);

LUT6 #(
   .INIT(64'h7cfa5bb87cfa5bb8)  
) LUT6_inst8419 (
   .O(to_level3[643]),
   .I0(level4_in[3858]),
   .I1(level4_in[3859]),
   .I2(level4_in[3860]),
   .I3(level4_in[3861]),
   .I4(level4_in[3862]),
   .I5(level4_in[3863])
);

LUT6 #(
   .INIT(64'hf695471ef695471e)  
) LUT6_inst8420 (
   .O(to_level3[644]),
   .I0(level4_in[3864]),
   .I1(level4_in[3865]),
   .I2(level4_in[3866]),
   .I3(level4_in[3867]),
   .I4(level4_in[3868]),
   .I5(level4_in[3869])
);

LUT6 #(
   .INIT(64'h9a164c379a164c37)  
) LUT6_inst8421 (
   .O(to_level3[645]),
   .I0(level4_in[3870]),
   .I1(level4_in[3871]),
   .I2(level4_in[3872]),
   .I3(level4_in[3873]),
   .I4(level4_in[3874]),
   .I5(level4_in[3875])
);

LUT6 #(
   .INIT(64'h0062e3b50062e3b5)  
) LUT6_inst8422 (
   .O(to_level3[646]),
   .I0(level4_in[3876]),
   .I1(level4_in[3877]),
   .I2(level4_in[3878]),
   .I3(level4_in[3879]),
   .I4(level4_in[3880]),
   .I5(level4_in[3881])
);

LUT6 #(
   .INIT(64'hd115ce1fd115ce1f)  
) LUT6_inst8423 (
   .O(to_level3[647]),
   .I0(level4_in[3882]),
   .I1(level4_in[3883]),
   .I2(level4_in[3884]),
   .I3(level4_in[3885]),
   .I4(level4_in[3886]),
   .I5(level4_in[3887])
);

LUT6 #(
   .INIT(64'h6496e8826496e882)  
) LUT6_inst8424 (
   .O(to_level3[648]),
   .I0(level4_in[3888]),
   .I1(level4_in[3889]),
   .I2(level4_in[3890]),
   .I3(level4_in[3891]),
   .I4(level4_in[3892]),
   .I5(level4_in[3893])
);

LUT6 #(
   .INIT(64'he81ba057e81ba057)  
) LUT6_inst8425 (
   .O(to_level3[649]),
   .I0(level4_in[3894]),
   .I1(level4_in[3895]),
   .I2(level4_in[3896]),
   .I3(level4_in[3897]),
   .I4(level4_in[3898]),
   .I5(level4_in[3899])
);

LUT6 #(
   .INIT(64'haeda98b9aeda98b9)  
) LUT6_inst8426 (
   .O(to_level3[650]),
   .I0(level4_in[3900]),
   .I1(level4_in[3901]),
   .I2(level4_in[3902]),
   .I3(level4_in[3903]),
   .I4(level4_in[3904]),
   .I5(level4_in[3905])
);

LUT6 #(
   .INIT(64'h004ec807004ec807)  
) LUT6_inst8427 (
   .O(to_level3[651]),
   .I0(level4_in[3906]),
   .I1(level4_in[3907]),
   .I2(level4_in[3908]),
   .I3(level4_in[3909]),
   .I4(level4_in[3910]),
   .I5(level4_in[3911])
);

LUT6 #(
   .INIT(64'h1ea8ac731ea8ac73)  
) LUT6_inst8428 (
   .O(to_level3[652]),
   .I0(level4_in[3912]),
   .I1(level4_in[3913]),
   .I2(level4_in[3914]),
   .I3(level4_in[3915]),
   .I4(level4_in[3916]),
   .I5(level4_in[3917])
);

LUT6 #(
   .INIT(64'hf13c9c5bf13c9c5b)  
) LUT6_inst8429 (
   .O(to_level3[653]),
   .I0(level4_in[3918]),
   .I1(level4_in[3919]),
   .I2(level4_in[3920]),
   .I3(level4_in[3921]),
   .I4(level4_in[3922]),
   .I5(level4_in[3923])
);

LUT6 #(
   .INIT(64'h962b1376962b1376)  
) LUT6_inst8430 (
   .O(to_level3[654]),
   .I0(level4_in[3924]),
   .I1(level4_in[3925]),
   .I2(level4_in[3926]),
   .I3(level4_in[3927]),
   .I4(level4_in[3928]),
   .I5(level4_in[3929])
);

LUT6 #(
   .INIT(64'h3166c9c33166c9c3)  
) LUT6_inst8431 (
   .O(to_level3[655]),
   .I0(level4_in[3930]),
   .I1(level4_in[3931]),
   .I2(level4_in[3932]),
   .I3(level4_in[3933]),
   .I4(level4_in[3934]),
   .I5(level4_in[3935])
);

LUT6 #(
   .INIT(64'hc755883cc755883c)  
) LUT6_inst8432 (
   .O(to_level3[656]),
   .I0(level4_in[3936]),
   .I1(level4_in[3937]),
   .I2(level4_in[3938]),
   .I3(level4_in[3939]),
   .I4(level4_in[3940]),
   .I5(level4_in[3941])
);

LUT6 #(
   .INIT(64'h2cf8c0582cf8c058)  
) LUT6_inst8433 (
   .O(to_level3[657]),
   .I0(level4_in[3942]),
   .I1(level4_in[3943]),
   .I2(level4_in[3944]),
   .I3(level4_in[3945]),
   .I4(level4_in[3946]),
   .I5(level4_in[3947])
);

LUT6 #(
   .INIT(64'h122a3271122a3271)  
) LUT6_inst8434 (
   .O(to_level3[658]),
   .I0(level4_in[3948]),
   .I1(level4_in[3949]),
   .I2(level4_in[3950]),
   .I3(level4_in[3951]),
   .I4(level4_in[3952]),
   .I5(level4_in[3953])
);

LUT6 #(
   .INIT(64'hf487c09bf487c09b)  
) LUT6_inst8435 (
   .O(to_level3[659]),
   .I0(level4_in[3954]),
   .I1(level4_in[3955]),
   .I2(level4_in[3956]),
   .I3(level4_in[3957]),
   .I4(level4_in[3958]),
   .I5(level4_in[3959])
);

LUT6 #(
   .INIT(64'h3b8823eb3b8823eb)  
) LUT6_inst8436 (
   .O(to_level3[660]),
   .I0(level4_in[3960]),
   .I1(level4_in[3961]),
   .I2(level4_in[3962]),
   .I3(level4_in[3963]),
   .I4(level4_in[3964]),
   .I5(level4_in[3965])
);

LUT6 #(
   .INIT(64'hf457beb9f457beb9)  
) LUT6_inst8437 (
   .O(to_level3[661]),
   .I0(level4_in[3966]),
   .I1(level4_in[3967]),
   .I2(level4_in[3968]),
   .I3(level4_in[3969]),
   .I4(level4_in[3970]),
   .I5(level4_in[3971])
);

LUT6 #(
   .INIT(64'ha0d44374a0d44374)  
) LUT6_inst8438 (
   .O(to_level3[662]),
   .I0(level4_in[3972]),
   .I1(level4_in[3973]),
   .I2(level4_in[3974]),
   .I3(level4_in[3975]),
   .I4(level4_in[3976]),
   .I5(level4_in[3977])
);

LUT6 #(
   .INIT(64'ha1599fbaa1599fba)  
) LUT6_inst8439 (
   .O(to_level3[663]),
   .I0(level4_in[3978]),
   .I1(level4_in[3979]),
   .I2(level4_in[3980]),
   .I3(level4_in[3981]),
   .I4(level4_in[3982]),
   .I5(level4_in[3983])
);

LUT6 #(
   .INIT(64'h6184b4746184b474)  
) LUT6_inst8440 (
   .O(to_level3[664]),
   .I0(level4_in[3984]),
   .I1(level4_in[3985]),
   .I2(level4_in[3986]),
   .I3(level4_in[3987]),
   .I4(level4_in[3988]),
   .I5(level4_in[3989])
);

LUT6 #(
   .INIT(64'hff71758aff71758a)  
) LUT6_inst8441 (
   .O(to_level3[665]),
   .I0(level4_in[3990]),
   .I1(level4_in[3991]),
   .I2(level4_in[3992]),
   .I3(level4_in[3993]),
   .I4(level4_in[3994]),
   .I5(level4_in[3995])
);

LUT6 #(
   .INIT(64'hccb694ccccb694cc)  
) LUT6_inst8442 (
   .O(to_level3[666]),
   .I0(level4_in[3996]),
   .I1(level4_in[3997]),
   .I2(level4_in[3998]),
   .I3(level4_in[3999]),
   .I4(level4_in[4000]),
   .I5(level4_in[4001])
);

LUT6 #(
   .INIT(64'h2bb195222bb19522)  
) LUT6_inst8443 (
   .O(to_level3[667]),
   .I0(level4_in[4002]),
   .I1(level4_in[4003]),
   .I2(level4_in[4004]),
   .I3(level4_in[4005]),
   .I4(level4_in[4006]),
   .I5(level4_in[4007])
);

LUT6 #(
   .INIT(64'h850c41de850c41de)  
) LUT6_inst8444 (
   .O(to_level3[668]),
   .I0(level4_in[4008]),
   .I1(level4_in[4009]),
   .I2(level4_in[4010]),
   .I3(level4_in[4011]),
   .I4(level4_in[4012]),
   .I5(level4_in[4013])
);

LUT6 #(
   .INIT(64'h1a27a6c11a27a6c1)  
) LUT6_inst8445 (
   .O(to_level3[669]),
   .I0(level4_in[4014]),
   .I1(level4_in[4015]),
   .I2(level4_in[4016]),
   .I3(level4_in[4017]),
   .I4(level4_in[4018]),
   .I5(level4_in[4019])
);

LUT6 #(
   .INIT(64'h15d6c5ea15d6c5ea)  
) LUT6_inst8446 (
   .O(to_level3[670]),
   .I0(level4_in[4020]),
   .I1(level4_in[4021]),
   .I2(level4_in[4022]),
   .I3(level4_in[4023]),
   .I4(level4_in[4024]),
   .I5(level4_in[4025])
);

LUT6 #(
   .INIT(64'h4b11c5d74b11c5d7)  
) LUT6_inst8447 (
   .O(to_level3[671]),
   .I0(level4_in[4026]),
   .I1(level4_in[4027]),
   .I2(level4_in[4028]),
   .I3(level4_in[4029]),
   .I4(level4_in[4030]),
   .I5(level4_in[4031])
);

LUT6 #(
   .INIT(64'hce3d61e5ce3d61e5)  
) LUT6_inst8448 (
   .O(to_level3[672]),
   .I0(level4_in[4032]),
   .I1(level4_in[4033]),
   .I2(level4_in[4034]),
   .I3(level4_in[4035]),
   .I4(level4_in[4036]),
   .I5(level4_in[4037])
);

LUT6 #(
   .INIT(64'h2b6ac4632b6ac463)  
) LUT6_inst8449 (
   .O(to_level3[673]),
   .I0(level4_in[4038]),
   .I1(level4_in[4039]),
   .I2(level4_in[4040]),
   .I3(level4_in[4041]),
   .I4(level4_in[4042]),
   .I5(level4_in[4043])
);

LUT6 #(
   .INIT(64'ha86b4606a86b4606)  
) LUT6_inst8450 (
   .O(to_level3[674]),
   .I0(level4_in[4044]),
   .I1(level4_in[4045]),
   .I2(level4_in[4046]),
   .I3(level4_in[4047]),
   .I4(level4_in[4048]),
   .I5(level4_in[4049])
);

LUT6 #(
   .INIT(64'h1455f1c41455f1c4)  
) LUT6_inst8451 (
   .O(to_level3[675]),
   .I0(level4_in[4050]),
   .I1(level4_in[4051]),
   .I2(level4_in[4052]),
   .I3(level4_in[4053]),
   .I4(level4_in[4054]),
   .I5(level4_in[4055])
);

LUT6 #(
   .INIT(64'hba834e5bba834e5b)  
) LUT6_inst8452 (
   .O(to_level3[676]),
   .I0(level4_in[4056]),
   .I1(level4_in[4057]),
   .I2(level4_in[4058]),
   .I3(level4_in[4059]),
   .I4(level4_in[4060]),
   .I5(level4_in[4061])
);

LUT6 #(
   .INIT(64'h61c5c13c61c5c13c)  
) LUT6_inst8453 (
   .O(to_level3[677]),
   .I0(level4_in[4062]),
   .I1(level4_in[4063]),
   .I2(level4_in[4064]),
   .I3(level4_in[4065]),
   .I4(level4_in[4066]),
   .I5(level4_in[4067])
);

LUT6 #(
   .INIT(64'h4523386a4523386a)  
) LUT6_inst8454 (
   .O(to_level3[678]),
   .I0(level4_in[4068]),
   .I1(level4_in[4069]),
   .I2(level4_in[4070]),
   .I3(level4_in[4071]),
   .I4(level4_in[4072]),
   .I5(level4_in[4073])
);

LUT6 #(
   .INIT(64'hb0887aa6b0887aa6)  
) LUT6_inst8455 (
   .O(to_level3[679]),
   .I0(level4_in[4074]),
   .I1(level4_in[4075]),
   .I2(level4_in[4076]),
   .I3(level4_in[4077]),
   .I4(level4_in[4078]),
   .I5(level4_in[4079])
);

LUT6 #(
   .INIT(64'heff5efd4eff5efd4)  
) LUT6_inst8456 (
   .O(to_level3[680]),
   .I0(level4_in[4080]),
   .I1(level4_in[4081]),
   .I2(level4_in[4082]),
   .I3(level4_in[4083]),
   .I4(level4_in[4084]),
   .I5(level4_in[4085])
);

LUT6 #(
   .INIT(64'hf3306e0ef3306e0e)  
) LUT6_inst8457 (
   .O(to_level3[681]),
   .I0(level4_in[4086]),
   .I1(level4_in[4087]),
   .I2(level4_in[4088]),
   .I3(level4_in[4089]),
   .I4(level4_in[4090]),
   .I5(level4_in[4091])
);

LUT6 #(
   .INIT(64'h5a4e4a065a4e4a06)  
) LUT6_inst8458 (
   .O(to_level3[682]),
   .I0(level4_in[4092]),
   .I1(level4_in[4093]),
   .I2(level4_in[4094]),
   .I3(level4_in[4095]),
   .I4(level4_in[4096]),
   .I5(level4_in[4097])
);

LUT6 #(
   .INIT(64'h8360443f8360443f)  
) LUT6_inst8459 (
   .O(to_level3[683]),
   .I0(level4_in[4098]),
   .I1(level4_in[4099]),
   .I2(level4_in[4100]),
   .I3(level4_in[4101]),
   .I4(level4_in[4102]),
   .I5(level4_in[4103])
);

LUT6 #(
   .INIT(64'h0fd6beeb0fd6beeb)  
) LUT6_inst8460 (
   .O(to_level3[684]),
   .I0(level4_in[4104]),
   .I1(level4_in[4105]),
   .I2(level4_in[4106]),
   .I3(level4_in[4107]),
   .I4(level4_in[4108]),
   .I5(level4_in[4109])
);

LUT6 #(
   .INIT(64'h51f1017c51f1017c)  
) LUT6_inst8461 (
   .O(to_level3[685]),
   .I0(level4_in[4110]),
   .I1(level4_in[4111]),
   .I2(level4_in[4112]),
   .I3(level4_in[4113]),
   .I4(level4_in[4114]),
   .I5(level4_in[4115])
);

LUT6 #(
   .INIT(64'h0944ef0d0944ef0d)  
) LUT6_inst8462 (
   .O(to_level3[686]),
   .I0(level4_in[4116]),
   .I1(level4_in[4117]),
   .I2(level4_in[4118]),
   .I3(level4_in[4119]),
   .I4(level4_in[4120]),
   .I5(level4_in[4121])
);

LUT6 #(
   .INIT(64'h19f0221819f02218)  
) LUT6_inst8463 (
   .O(to_level3[687]),
   .I0(level4_in[4122]),
   .I1(level4_in[4123]),
   .I2(level4_in[4124]),
   .I3(level4_in[4125]),
   .I4(level4_in[4126]),
   .I5(level4_in[4127])
);

LUT6 #(
   .INIT(64'h10e7050d10e7050d)  
) LUT6_inst8464 (
   .O(to_level3[688]),
   .I0(level4_in[4128]),
   .I1(level4_in[4129]),
   .I2(level4_in[4130]),
   .I3(level4_in[4131]),
   .I4(level4_in[4132]),
   .I5(level4_in[4133])
);

LUT6 #(
   .INIT(64'h23c89b0123c89b01)  
) LUT6_inst8465 (
   .O(to_level3[689]),
   .I0(level4_in[4134]),
   .I1(level4_in[4135]),
   .I2(level4_in[4136]),
   .I3(level4_in[4137]),
   .I4(level4_in[4138]),
   .I5(level4_in[4139])
);

LUT6 #(
   .INIT(64'hef2d1849ef2d1849)  
) LUT6_inst8466 (
   .O(to_level3[690]),
   .I0(level4_in[4140]),
   .I1(level4_in[4141]),
   .I2(level4_in[4142]),
   .I3(level4_in[4143]),
   .I4(level4_in[4144]),
   .I5(level4_in[4145])
);

LUT6 #(
   .INIT(64'hf68849bbf68849bb)  
) LUT6_inst8467 (
   .O(to_level3[691]),
   .I0(level4_in[4146]),
   .I1(level4_in[4147]),
   .I2(level4_in[4148]),
   .I3(level4_in[4149]),
   .I4(level4_in[4150]),
   .I5(level4_in[4151])
);

LUT6 #(
   .INIT(64'h2353bc8d2353bc8d)  
) LUT6_inst8468 (
   .O(to_level3[692]),
   .I0(level4_in[4152]),
   .I1(level4_in[4153]),
   .I2(level4_in[4154]),
   .I3(level4_in[4155]),
   .I4(level4_in[4156]),
   .I5(level4_in[4157])
);

LUT6 #(
   .INIT(64'h09d3d23a09d3d23a)  
) LUT6_inst8469 (
   .O(to_level3[693]),
   .I0(level4_in[4158]),
   .I1(level4_in[4159]),
   .I2(level4_in[4160]),
   .I3(level4_in[4161]),
   .I4(level4_in[4162]),
   .I5(level4_in[4163])
);

LUT6 #(
   .INIT(64'ha02b8886a02b8886)  
) LUT6_inst8470 (
   .O(to_level3[694]),
   .I0(level4_in[4164]),
   .I1(level4_in[4165]),
   .I2(level4_in[4166]),
   .I3(level4_in[4167]),
   .I4(level4_in[4168]),
   .I5(level4_in[4169])
);

LUT6 #(
   .INIT(64'h0704dd890704dd89)  
) LUT6_inst8471 (
   .O(to_level3[695]),
   .I0(level4_in[4170]),
   .I1(level4_in[4171]),
   .I2(level4_in[4172]),
   .I3(level4_in[4173]),
   .I4(level4_in[4174]),
   .I5(level4_in[4175])
);

LUT6 #(
   .INIT(64'h61a54fa261a54fa2)  
) LUT6_inst8472 (
   .O(to_level3[696]),
   .I0(level4_in[4176]),
   .I1(level4_in[4177]),
   .I2(level4_in[4178]),
   .I3(level4_in[4179]),
   .I4(level4_in[4180]),
   .I5(level4_in[4181])
);

LUT6 #(
   .INIT(64'hfd9d0a79fd9d0a79)  
) LUT6_inst8473 (
   .O(to_level3[697]),
   .I0(level4_in[4182]),
   .I1(level4_in[4183]),
   .I2(level4_in[4184]),
   .I3(level4_in[4185]),
   .I4(level4_in[4186]),
   .I5(level4_in[4187])
);

LUT6 #(
   .INIT(64'hfa3ea196fa3ea196)  
) LUT6_inst8474 (
   .O(to_level3[698]),
   .I0(level4_in[4188]),
   .I1(level4_in[4189]),
   .I2(level4_in[4190]),
   .I3(level4_in[4191]),
   .I4(level4_in[4192]),
   .I5(level4_in[4193])
);

LUT6 #(
   .INIT(64'h32bd52d732bd52d7)  
) LUT6_inst8475 (
   .O(to_level3[699]),
   .I0(level4_in[4194]),
   .I1(level4_in[4195]),
   .I2(level4_in[4196]),
   .I3(level4_in[4197]),
   .I4(level4_in[4198]),
   .I5(level4_in[4199])
);

LUT6 #(
   .INIT(64'h4bd2daa94bd2daa9)  
) LUT6_inst8476 (
   .O(to_level3[700]),
   .I0(level4_in[4200]),
   .I1(level4_in[4201]),
   .I2(level4_in[4202]),
   .I3(level4_in[4203]),
   .I4(level4_in[4204]),
   .I5(level4_in[4205])
);

LUT6 #(
   .INIT(64'he1fc19e6e1fc19e6)  
) LUT6_inst8477 (
   .O(to_level3[701]),
   .I0(level4_in[4206]),
   .I1(level4_in[4207]),
   .I2(level4_in[4208]),
   .I3(level4_in[4209]),
   .I4(level4_in[4210]),
   .I5(level4_in[4211])
);

LUT6 #(
   .INIT(64'hf35166fef35166fe)  
) LUT6_inst8478 (
   .O(to_level3[702]),
   .I0(level4_in[4212]),
   .I1(level4_in[4213]),
   .I2(level4_in[4214]),
   .I3(level4_in[4215]),
   .I4(level4_in[4216]),
   .I5(level4_in[4217])
);

LUT6 #(
   .INIT(64'hb4271efcb4271efc)  
) LUT6_inst8479 (
   .O(to_level3[703]),
   .I0(level4_in[4218]),
   .I1(level4_in[4219]),
   .I2(level4_in[4220]),
   .I3(level4_in[4221]),
   .I4(level4_in[4222]),
   .I5(level4_in[4223])
);

LUT6 #(
   .INIT(64'h4d4d57814d4d5781)  
) LUT6_inst8480 (
   .O(to_level3[704]),
   .I0(level4_in[4224]),
   .I1(level4_in[4225]),
   .I2(level4_in[4226]),
   .I3(level4_in[4227]),
   .I4(level4_in[4228]),
   .I5(level4_in[4229])
);

LUT6 #(
   .INIT(64'h2e74c3db2e74c3db)  
) LUT6_inst8481 (
   .O(to_level3[705]),
   .I0(level4_in[4230]),
   .I1(level4_in[4231]),
   .I2(level4_in[4232]),
   .I3(level4_in[4233]),
   .I4(level4_in[4234]),
   .I5(level4_in[4235])
);

LUT6 #(
   .INIT(64'h992d7c5a992d7c5a)  
) LUT6_inst8482 (
   .O(to_level3[706]),
   .I0(level4_in[4236]),
   .I1(level4_in[4237]),
   .I2(level4_in[4238]),
   .I3(level4_in[4239]),
   .I4(level4_in[4240]),
   .I5(level4_in[4241])
);

LUT6 #(
   .INIT(64'hc47427e8c47427e8)  
) LUT6_inst8483 (
   .O(to_level3[707]),
   .I0(level4_in[4242]),
   .I1(level4_in[4243]),
   .I2(level4_in[4244]),
   .I3(level4_in[4245]),
   .I4(level4_in[4246]),
   .I5(level4_in[4247])
);

LUT6 #(
   .INIT(64'h27b3425f27b3425f)  
) LUT6_inst8484 (
   .O(to_level3[708]),
   .I0(level4_in[4248]),
   .I1(level4_in[4249]),
   .I2(level4_in[4250]),
   .I3(level4_in[4251]),
   .I4(level4_in[4252]),
   .I5(level4_in[4253])
);

LUT6 #(
   .INIT(64'h07a5404907a54049)  
) LUT6_inst8485 (
   .O(to_level3[709]),
   .I0(level4_in[4254]),
   .I1(level4_in[4255]),
   .I2(level4_in[4256]),
   .I3(level4_in[4257]),
   .I4(level4_in[4258]),
   .I5(level4_in[4259])
);

LUT6 #(
   .INIT(64'h42b728f842b728f8)  
) LUT6_inst8486 (
   .O(to_level3[710]),
   .I0(level4_in[4260]),
   .I1(level4_in[4261]),
   .I2(level4_in[4262]),
   .I3(level4_in[4263]),
   .I4(level4_in[4264]),
   .I5(level4_in[4265])
);

LUT6 #(
   .INIT(64'hc01204ccc01204cc)  
) LUT6_inst8487 (
   .O(to_level3[711]),
   .I0(level4_in[4266]),
   .I1(level4_in[4267]),
   .I2(level4_in[4268]),
   .I3(level4_in[4269]),
   .I4(level4_in[4270]),
   .I5(level4_in[4271])
);

LUT6 #(
   .INIT(64'ha650b9fda650b9fd)  
) LUT6_inst8488 (
   .O(to_level3[712]),
   .I0(level4_in[4272]),
   .I1(level4_in[4273]),
   .I2(level4_in[4274]),
   .I3(level4_in[4275]),
   .I4(level4_in[4276]),
   .I5(level4_in[4277])
);

LUT6 #(
   .INIT(64'h17da954317da9543)  
) LUT6_inst8489 (
   .O(to_level3[713]),
   .I0(level4_in[4278]),
   .I1(level4_in[4279]),
   .I2(level4_in[4280]),
   .I3(level4_in[4281]),
   .I4(level4_in[4282]),
   .I5(level4_in[4283])
);

LUT6 #(
   .INIT(64'h6e408c5c6e408c5c)  
) LUT6_inst8490 (
   .O(to_level3[714]),
   .I0(level4_in[4284]),
   .I1(level4_in[4285]),
   .I2(level4_in[4286]),
   .I3(level4_in[4287]),
   .I4(level4_in[4288]),
   .I5(level4_in[4289])
);

LUT6 #(
   .INIT(64'h60db1b8e60db1b8e)  
) LUT6_inst8491 (
   .O(to_level3[715]),
   .I0(level4_in[4290]),
   .I1(level4_in[4291]),
   .I2(level4_in[4292]),
   .I3(level4_in[4293]),
   .I4(level4_in[4294]),
   .I5(level4_in[4295])
);

LUT6 #(
   .INIT(64'hedcc8817edcc8817)  
) LUT6_inst8492 (
   .O(to_level3[716]),
   .I0(level4_in[4296]),
   .I1(level4_in[4297]),
   .I2(level4_in[4298]),
   .I3(level4_in[4299]),
   .I4(level4_in[4300]),
   .I5(level4_in[4301])
);

LUT6 #(
   .INIT(64'he27d4ba4e27d4ba4)  
) LUT6_inst8493 (
   .O(to_level3[717]),
   .I0(level4_in[4302]),
   .I1(level4_in[4303]),
   .I2(level4_in[4304]),
   .I3(level4_in[4305]),
   .I4(level4_in[4306]),
   .I5(level4_in[4307])
);

LUT6 #(
   .INIT(64'h75b710bd75b710bd)  
) LUT6_inst8494 (
   .O(to_level3[718]),
   .I0(level4_in[4308]),
   .I1(level4_in[4309]),
   .I2(level4_in[4310]),
   .I3(level4_in[4311]),
   .I4(level4_in[4312]),
   .I5(level4_in[4313])
);

LUT6 #(
   .INIT(64'h641834fb641834fb)  
) LUT6_inst8495 (
   .O(to_level3[719]),
   .I0(level4_in[4314]),
   .I1(level4_in[4315]),
   .I2(level4_in[4316]),
   .I3(level4_in[4317]),
   .I4(level4_in[4318]),
   .I5(level4_in[4319])
);

LUT6 #(
   .INIT(64'h07fb3d9207fb3d92)  
) LUT6_inst8496 (
   .O(to_level3[720]),
   .I0(level4_in[4320]),
   .I1(level4_in[4321]),
   .I2(level4_in[4322]),
   .I3(level4_in[4323]),
   .I4(level4_in[4324]),
   .I5(level4_in[4325])
);

LUT6 #(
   .INIT(64'h6592994765929947)  
) LUT6_inst8497 (
   .O(to_level3[721]),
   .I0(level4_in[4326]),
   .I1(level4_in[4327]),
   .I2(level4_in[4328]),
   .I3(level4_in[4329]),
   .I4(level4_in[4330]),
   .I5(level4_in[4331])
);

LUT6 #(
   .INIT(64'h5735492957354929)  
) LUT6_inst8498 (
   .O(to_level3[722]),
   .I0(level4_in[4332]),
   .I1(level4_in[4333]),
   .I2(level4_in[4334]),
   .I3(level4_in[4335]),
   .I4(level4_in[4336]),
   .I5(level4_in[4337])
);

LUT6 #(
   .INIT(64'h956ae7e1956ae7e1)  
) LUT6_inst8499 (
   .O(to_level3[723]),
   .I0(level4_in[4338]),
   .I1(level4_in[4339]),
   .I2(level4_in[4340]),
   .I3(level4_in[4341]),
   .I4(level4_in[4342]),
   .I5(level4_in[4343])
);

LUT6 #(
   .INIT(64'h596dc6e2596dc6e2)  
) LUT6_inst8500 (
   .O(to_level3[724]),
   .I0(level4_in[4344]),
   .I1(level4_in[4345]),
   .I2(level4_in[4346]),
   .I3(level4_in[4347]),
   .I4(level4_in[4348]),
   .I5(level4_in[4349])
);

LUT6 #(
   .INIT(64'h839d76d0839d76d0)  
) LUT6_inst8501 (
   .O(to_level3[725]),
   .I0(level4_in[4350]),
   .I1(level4_in[4351]),
   .I2(level4_in[4352]),
   .I3(level4_in[4353]),
   .I4(level4_in[4354]),
   .I5(level4_in[4355])
);

LUT6 #(
   .INIT(64'hec62fdbfec62fdbf)  
) LUT6_inst8502 (
   .O(to_level3[726]),
   .I0(level4_in[4356]),
   .I1(level4_in[4357]),
   .I2(level4_in[4358]),
   .I3(level4_in[4359]),
   .I4(level4_in[4360]),
   .I5(level4_in[4361])
);

LUT6 #(
   .INIT(64'h23e38df523e38df5)  
) LUT6_inst8503 (
   .O(to_level3[727]),
   .I0(level4_in[4362]),
   .I1(level4_in[4363]),
   .I2(level4_in[4364]),
   .I3(level4_in[4365]),
   .I4(level4_in[4366]),
   .I5(level4_in[4367])
);

LUT6 #(
   .INIT(64'h41c022a341c022a3)  
) LUT6_inst8504 (
   .O(to_level3[728]),
   .I0(level4_in[4368]),
   .I1(level4_in[4369]),
   .I2(level4_in[4370]),
   .I3(level4_in[4371]),
   .I4(level4_in[4372]),
   .I5(level4_in[4373])
);

LUT6 #(
   .INIT(64'h7a3a8d047a3a8d04)  
) LUT6_inst8505 (
   .O(to_level3[729]),
   .I0(level4_in[4374]),
   .I1(level4_in[4375]),
   .I2(level4_in[4376]),
   .I3(level4_in[4377]),
   .I4(level4_in[4378]),
   .I5(level4_in[4379])
);

LUT6 #(
   .INIT(64'h2740c3772740c377)  
) LUT6_inst8506 (
   .O(to_level3[730]),
   .I0(level4_in[4380]),
   .I1(level4_in[4381]),
   .I2(level4_in[4382]),
   .I3(level4_in[4383]),
   .I4(level4_in[4384]),
   .I5(level4_in[4385])
);

LUT6 #(
   .INIT(64'h372ffebe372ffebe)  
) LUT6_inst8507 (
   .O(to_level3[731]),
   .I0(level4_in[4386]),
   .I1(level4_in[4387]),
   .I2(level4_in[4388]),
   .I3(level4_in[4389]),
   .I4(level4_in[4390]),
   .I5(level4_in[4391])
);

LUT6 #(
   .INIT(64'h946eaf46946eaf46)  
) LUT6_inst8508 (
   .O(to_level3[732]),
   .I0(level4_in[4392]),
   .I1(level4_in[4393]),
   .I2(level4_in[4394]),
   .I3(level4_in[4395]),
   .I4(level4_in[4396]),
   .I5(level4_in[4397])
);

LUT6 #(
   .INIT(64'h7fa5e63e7fa5e63e)  
) LUT6_inst8509 (
   .O(to_level3[733]),
   .I0(level4_in[4398]),
   .I1(level4_in[4399]),
   .I2(level4_in[4400]),
   .I3(level4_in[4401]),
   .I4(level4_in[4402]),
   .I5(level4_in[4403])
);

LUT6 #(
   .INIT(64'h5041f2395041f239)  
) LUT6_inst8510 (
   .O(to_level3[734]),
   .I0(level4_in[4404]),
   .I1(level4_in[4405]),
   .I2(level4_in[4406]),
   .I3(level4_in[4407]),
   .I4(level4_in[4408]),
   .I5(level4_in[4409])
);

LUT6 #(
   .INIT(64'h34e6b3bc34e6b3bc)  
) LUT6_inst8511 (
   .O(to_level3[735]),
   .I0(level4_in[4410]),
   .I1(level4_in[4411]),
   .I2(level4_in[4412]),
   .I3(level4_in[4413]),
   .I4(level4_in[4414]),
   .I5(level4_in[4415])
);

LUT6 #(
   .INIT(64'hffdc7e0effdc7e0e)  
) LUT6_inst8512 (
   .O(to_level3[736]),
   .I0(level4_in[4416]),
   .I1(level4_in[4417]),
   .I2(level4_in[4418]),
   .I3(level4_in[4419]),
   .I4(level4_in[4420]),
   .I5(level4_in[4421])
);

LUT6 #(
   .INIT(64'h01867afd01867afd)  
) LUT6_inst8513 (
   .O(to_level3[737]),
   .I0(level4_in[4422]),
   .I1(level4_in[4423]),
   .I2(level4_in[4424]),
   .I3(level4_in[4425]),
   .I4(level4_in[4426]),
   .I5(level4_in[4427])
);

LUT6 #(
   .INIT(64'hca2073b4ca2073b4)  
) LUT6_inst8514 (
   .O(to_level3[738]),
   .I0(level4_in[4428]),
   .I1(level4_in[4429]),
   .I2(level4_in[4430]),
   .I3(level4_in[4431]),
   .I4(level4_in[4432]),
   .I5(level4_in[4433])
);

LUT6 #(
   .INIT(64'ha49ff83ea49ff83e)  
) LUT6_inst8515 (
   .O(to_level3[739]),
   .I0(level4_in[4434]),
   .I1(level4_in[4435]),
   .I2(level4_in[4436]),
   .I3(level4_in[4437]),
   .I4(level4_in[4438]),
   .I5(level4_in[4439])
);

LUT6 #(
   .INIT(64'h5a2d4d345a2d4d34)  
) LUT6_inst8516 (
   .O(to_level3[740]),
   .I0(level4_in[4440]),
   .I1(level4_in[4441]),
   .I2(level4_in[4442]),
   .I3(level4_in[4443]),
   .I4(level4_in[4444]),
   .I5(level4_in[4445])
);

LUT6 #(
   .INIT(64'hb7dfd486b7dfd486)  
) LUT6_inst8517 (
   .O(to_level3[741]),
   .I0(level4_in[4446]),
   .I1(level4_in[4447]),
   .I2(level4_in[4448]),
   .I3(level4_in[4449]),
   .I4(level4_in[4450]),
   .I5(level4_in[4451])
);

LUT6 #(
   .INIT(64'h1027edbb1027edbb)  
) LUT6_inst8518 (
   .O(to_level3[742]),
   .I0(level4_in[4452]),
   .I1(level4_in[4453]),
   .I2(level4_in[4454]),
   .I3(level4_in[4455]),
   .I4(level4_in[4456]),
   .I5(level4_in[4457])
);

LUT6 #(
   .INIT(64'h3adcb59b3adcb59b)  
) LUT6_inst8519 (
   .O(to_level3[743]),
   .I0(level4_in[4458]),
   .I1(level4_in[4459]),
   .I2(level4_in[4460]),
   .I3(level4_in[4461]),
   .I4(level4_in[4462]),
   .I5(level4_in[4463])
);

LUT6 #(
   .INIT(64'he3c17fe5e3c17fe5)  
) LUT6_inst8520 (
   .O(to_level3[744]),
   .I0(level4_in[4464]),
   .I1(level4_in[4465]),
   .I2(level4_in[4466]),
   .I3(level4_in[4467]),
   .I4(level4_in[4468]),
   .I5(level4_in[4469])
);

LUT6 #(
   .INIT(64'h5ef13f215ef13f21)  
) LUT6_inst8521 (
   .O(to_level3[745]),
   .I0(level4_in[4470]),
   .I1(level4_in[4471]),
   .I2(level4_in[4472]),
   .I3(level4_in[4473]),
   .I4(level4_in[4474]),
   .I5(level4_in[4475])
);

LUT6 #(
   .INIT(64'he50a69d6e50a69d6)  
) LUT6_inst8522 (
   .O(to_level3[746]),
   .I0(level4_in[4476]),
   .I1(level4_in[4477]),
   .I2(level4_in[4478]),
   .I3(level4_in[4479]),
   .I4(level4_in[4480]),
   .I5(level4_in[4481])
);

LUT6 #(
   .INIT(64'hc0ca570ec0ca570e)  
) LUT6_inst8523 (
   .O(to_level3[747]),
   .I0(level4_in[4482]),
   .I1(level4_in[4483]),
   .I2(level4_in[4484]),
   .I3(level4_in[4485]),
   .I4(level4_in[4486]),
   .I5(level4_in[4487])
);

LUT6 #(
   .INIT(64'he1832433e1832433)  
) LUT6_inst8524 (
   .O(to_level3[748]),
   .I0(level4_in[4488]),
   .I1(level4_in[4489]),
   .I2(level4_in[4490]),
   .I3(level4_in[4491]),
   .I4(level4_in[4492]),
   .I5(level4_in[4493])
);

LUT6 #(
   .INIT(64'hc0da551bc0da551b)  
) LUT6_inst8525 (
   .O(to_level3[749]),
   .I0(level4_in[4494]),
   .I1(level4_in[4495]),
   .I2(level4_in[4496]),
   .I3(level4_in[4497]),
   .I4(level4_in[4498]),
   .I5(level4_in[4499])
);

LUT6 #(
   .INIT(64'h15ace27015ace270)  
) LUT6_inst8526 (
   .O(to_level3[750]),
   .I0(level4_in[4500]),
   .I1(level4_in[4501]),
   .I2(level4_in[4502]),
   .I3(level4_in[4503]),
   .I4(level4_in[4504]),
   .I5(level4_in[4505])
);

LUT6 #(
   .INIT(64'h4cf618954cf61895)  
) LUT6_inst8527 (
   .O(to_level3[751]),
   .I0(level4_in[4506]),
   .I1(level4_in[4507]),
   .I2(level4_in[4508]),
   .I3(level4_in[4509]),
   .I4(level4_in[4510]),
   .I5(level4_in[4511])
);

LUT6 #(
   .INIT(64'ha6ab1d05a6ab1d05)  
) LUT6_inst8528 (
   .O(to_level3[752]),
   .I0(level4_in[4512]),
   .I1(level4_in[4513]),
   .I2(level4_in[4514]),
   .I3(level4_in[4515]),
   .I4(level4_in[4516]),
   .I5(level4_in[4517])
);

LUT6 #(
   .INIT(64'h2c81d3452c81d345)  
) LUT6_inst8529 (
   .O(to_level3[753]),
   .I0(level4_in[4518]),
   .I1(level4_in[4519]),
   .I2(level4_in[4520]),
   .I3(level4_in[4521]),
   .I4(level4_in[4522]),
   .I5(level4_in[4523])
);

LUT6 #(
   .INIT(64'h939bff2b939bff2b)  
) LUT6_inst8530 (
   .O(to_level3[754]),
   .I0(level4_in[4524]),
   .I1(level4_in[4525]),
   .I2(level4_in[4526]),
   .I3(level4_in[4527]),
   .I4(level4_in[4528]),
   .I5(level4_in[4529])
);

LUT6 #(
   .INIT(64'hfa46c555fa46c555)  
) LUT6_inst8531 (
   .O(to_level3[755]),
   .I0(level4_in[4530]),
   .I1(level4_in[4531]),
   .I2(level4_in[4532]),
   .I3(level4_in[4533]),
   .I4(level4_in[4534]),
   .I5(level4_in[4535])
);

LUT6 #(
   .INIT(64'hd9cf8d44d9cf8d44)  
) LUT6_inst8532 (
   .O(to_level3[756]),
   .I0(level4_in[4536]),
   .I1(level4_in[4537]),
   .I2(level4_in[4538]),
   .I3(level4_in[4539]),
   .I4(level4_in[4540]),
   .I5(level4_in[4541])
);

LUT6 #(
   .INIT(64'habbec5b4abbec5b4)  
) LUT6_inst8533 (
   .O(to_level3[757]),
   .I0(level4_in[4542]),
   .I1(level4_in[4543]),
   .I2(level4_in[4544]),
   .I3(level4_in[4545]),
   .I4(level4_in[4546]),
   .I5(level4_in[4547])
);

LUT6 #(
   .INIT(64'h9eb2bd1a9eb2bd1a)  
) LUT6_inst8534 (
   .O(to_level3[758]),
   .I0(level4_in[4548]),
   .I1(level4_in[4549]),
   .I2(level4_in[4550]),
   .I3(level4_in[4551]),
   .I4(level4_in[4552]),
   .I5(level4_in[4553])
);

LUT6 #(
   .INIT(64'h2e1fea262e1fea26)  
) LUT6_inst8535 (
   .O(to_level3[759]),
   .I0(level4_in[4554]),
   .I1(level4_in[4555]),
   .I2(level4_in[4556]),
   .I3(level4_in[4557]),
   .I4(level4_in[4558]),
   .I5(level4_in[4559])
);

LUT6 #(
   .INIT(64'h2c0e96a12c0e96a1)  
) LUT6_inst8536 (
   .O(to_level3[760]),
   .I0(level4_in[4560]),
   .I1(level4_in[4561]),
   .I2(level4_in[4562]),
   .I3(level4_in[4563]),
   .I4(level4_in[4564]),
   .I5(level4_in[4565])
);

LUT6 #(
   .INIT(64'hbe721754be721754)  
) LUT6_inst8537 (
   .O(to_level3[761]),
   .I0(level4_in[4566]),
   .I1(level4_in[4567]),
   .I2(level4_in[4568]),
   .I3(level4_in[4569]),
   .I4(level4_in[4570]),
   .I5(level4_in[4571])
);

LUT6 #(
   .INIT(64'h5a2825885a282588)  
) LUT6_inst8538 (
   .O(to_level3[762]),
   .I0(level4_in[4572]),
   .I1(level4_in[4573]),
   .I2(level4_in[4574]),
   .I3(level4_in[4575]),
   .I4(level4_in[4576]),
   .I5(level4_in[4577])
);

LUT6 #(
   .INIT(64'h351194e4351194e4)  
) LUT6_inst8539 (
   .O(to_level3[763]),
   .I0(level4_in[4578]),
   .I1(level4_in[4579]),
   .I2(level4_in[4580]),
   .I3(level4_in[4581]),
   .I4(level4_in[4582]),
   .I5(level4_in[4583])
);

LUT6 #(
   .INIT(64'h77d7ebdf77d7ebdf)  
) LUT6_inst8540 (
   .O(to_level3[764]),
   .I0(level4_in[4584]),
   .I1(level4_in[4585]),
   .I2(level4_in[4586]),
   .I3(level4_in[4587]),
   .I4(level4_in[4588]),
   .I5(level4_in[4589])
);

LUT6 #(
   .INIT(64'hef3d17c3ef3d17c3)  
) LUT6_inst8541 (
   .O(to_level3[765]),
   .I0(level4_in[4590]),
   .I1(level4_in[4591]),
   .I2(level4_in[4592]),
   .I3(level4_in[4593]),
   .I4(level4_in[4594]),
   .I5(level4_in[4595])
);

LUT6 #(
   .INIT(64'h65b2b39365b2b393)  
) LUT6_inst8542 (
   .O(to_level3[766]),
   .I0(level4_in[4596]),
   .I1(level4_in[4597]),
   .I2(level4_in[4598]),
   .I3(level4_in[4599]),
   .I4(level4_in[4600]),
   .I5(level4_in[4601])
);

LUT6 #(
   .INIT(64'hd67aa03fd67aa03f)  
) LUT6_inst8543 (
   .O(to_level3[767]),
   .I0(level4_in[4602]),
   .I1(level4_in[4603]),
   .I2(level4_in[4604]),
   .I3(level4_in[4605]),
   .I4(level4_in[4606]),
   .I5(level4_in[4607])
);

LUT6 #(
   .INIT(64'hde15e086de15e086)  
) LUT6_inst8544 (
   .O(to_level3[768]),
   .I0(level4_in[4608]),
   .I1(level4_in[4609]),
   .I2(level4_in[4610]),
   .I3(level4_in[4611]),
   .I4(level4_in[4612]),
   .I5(level4_in[4613])
);

LUT6 #(
   .INIT(64'hdfc902d4dfc902d4)  
) LUT6_inst8545 (
   .O(to_level3[769]),
   .I0(level4_in[4614]),
   .I1(level4_in[4615]),
   .I2(level4_in[4616]),
   .I3(level4_in[4617]),
   .I4(level4_in[4618]),
   .I5(level4_in[4619])
);

LUT6 #(
   .INIT(64'h556f835c556f835c)  
) LUT6_inst8546 (
   .O(to_level3[770]),
   .I0(level4_in[4620]),
   .I1(level4_in[4621]),
   .I2(level4_in[4622]),
   .I3(level4_in[4623]),
   .I4(level4_in[4624]),
   .I5(level4_in[4625])
);

LUT6 #(
   .INIT(64'hc0b29ddfc0b29ddf)  
) LUT6_inst8547 (
   .O(to_level3[771]),
   .I0(level4_in[4626]),
   .I1(level4_in[4627]),
   .I2(level4_in[4628]),
   .I3(level4_in[4629]),
   .I4(level4_in[4630]),
   .I5(level4_in[4631])
);

LUT6 #(
   .INIT(64'h7a1d79037a1d7903)  
) LUT6_inst8548 (
   .O(to_level3[772]),
   .I0(level4_in[4632]),
   .I1(level4_in[4633]),
   .I2(level4_in[4634]),
   .I3(level4_in[4635]),
   .I4(level4_in[4636]),
   .I5(level4_in[4637])
);

LUT6 #(
   .INIT(64'h8a7ea7008a7ea700)  
) LUT6_inst8549 (
   .O(to_level3[773]),
   .I0(level4_in[4638]),
   .I1(level4_in[4639]),
   .I2(level4_in[4640]),
   .I3(level4_in[4641]),
   .I4(level4_in[4642]),
   .I5(level4_in[4643])
);

LUT6 #(
   .INIT(64'he8bd72bce8bd72bc)  
) LUT6_inst8550 (
   .O(to_level3[774]),
   .I0(level4_in[4644]),
   .I1(level4_in[4645]),
   .I2(level4_in[4646]),
   .I3(level4_in[4647]),
   .I4(level4_in[4648]),
   .I5(level4_in[4649])
);

LUT6 #(
   .INIT(64'h08e0883d08e0883d)  
) LUT6_inst8551 (
   .O(to_level3[775]),
   .I0(level4_in[4650]),
   .I1(level4_in[4651]),
   .I2(level4_in[4652]),
   .I3(level4_in[4653]),
   .I4(level4_in[4654]),
   .I5(level4_in[4655])
);

LUT6 #(
   .INIT(64'hbe625be7be625be7)  
) LUT6_inst8552 (
   .O(to_level3[776]),
   .I0(level4_in[4656]),
   .I1(level4_in[4657]),
   .I2(level4_in[4658]),
   .I3(level4_in[4659]),
   .I4(level4_in[4660]),
   .I5(level4_in[4661])
);

LUT6 #(
   .INIT(64'hd2e174e2d2e174e2)  
) LUT6_inst8553 (
   .O(to_level3[777]),
   .I0(level4_in[4662]),
   .I1(level4_in[4663]),
   .I2(level4_in[4664]),
   .I3(level4_in[4665]),
   .I4(level4_in[4666]),
   .I5(level4_in[4667])
);

LUT6 #(
   .INIT(64'h17960b8d17960b8d)  
) LUT6_inst8554 (
   .O(to_level3[778]),
   .I0(level4_in[4668]),
   .I1(level4_in[4669]),
   .I2(level4_in[4670]),
   .I3(level4_in[4671]),
   .I4(level4_in[4672]),
   .I5(level4_in[4673])
);

LUT6 #(
   .INIT(64'hbe4722d7be4722d7)  
) LUT6_inst8555 (
   .O(to_level3[779]),
   .I0(level4_in[4674]),
   .I1(level4_in[4675]),
   .I2(level4_in[4676]),
   .I3(level4_in[4677]),
   .I4(level4_in[4678]),
   .I5(level4_in[4679])
);

LUT6 #(
   .INIT(64'h0736ca480736ca48)  
) LUT6_inst8556 (
   .O(to_level3[780]),
   .I0(level4_in[4680]),
   .I1(level4_in[4681]),
   .I2(level4_in[4682]),
   .I3(level4_in[4683]),
   .I4(level4_in[4684]),
   .I5(level4_in[4685])
);

LUT6 #(
   .INIT(64'h042279dc042279dc)  
) LUT6_inst8557 (
   .O(to_level3[781]),
   .I0(level4_in[4686]),
   .I1(level4_in[4687]),
   .I2(level4_in[4688]),
   .I3(level4_in[4689]),
   .I4(level4_in[4690]),
   .I5(level4_in[4691])
);

LUT6 #(
   .INIT(64'hf13e5d80f13e5d80)  
) LUT6_inst8558 (
   .O(to_level3[782]),
   .I0(level4_in[4692]),
   .I1(level4_in[4693]),
   .I2(level4_in[4694]),
   .I3(level4_in[4695]),
   .I4(level4_in[4696]),
   .I5(level4_in[4697])
);

LUT6 #(
   .INIT(64'hfbb5e811fbb5e811)  
) LUT6_inst8559 (
   .O(to_level3[783]),
   .I0(level4_in[4698]),
   .I1(level4_in[4699]),
   .I2(level4_in[4700]),
   .I3(level4_in[4701]),
   .I4(level4_in[4702]),
   .I5(level4_in[4703])
);

LUT6 #(
   .INIT(64'h2703cd812703cd81)  
) LUT6_inst8560 (
   .O(to_level3[784]),
   .I0(level4_in[4704]),
   .I1(level4_in[4705]),
   .I2(level4_in[4706]),
   .I3(level4_in[4707]),
   .I4(level4_in[4708]),
   .I5(level4_in[4709])
);

LUT6 #(
   .INIT(64'h63af742363af7423)  
) LUT6_inst8561 (
   .O(to_level3[785]),
   .I0(level4_in[4710]),
   .I1(level4_in[4711]),
   .I2(level4_in[4712]),
   .I3(level4_in[4713]),
   .I4(level4_in[4714]),
   .I5(level4_in[4715])
);

LUT6 #(
   .INIT(64'hbf592468bf592468)  
) LUT6_inst8562 (
   .O(to_level3[786]),
   .I0(level4_in[4716]),
   .I1(level4_in[4717]),
   .I2(level4_in[4718]),
   .I3(level4_in[4719]),
   .I4(level4_in[4720]),
   .I5(level4_in[4721])
);

LUT6 #(
   .INIT(64'h3f46fc233f46fc23)  
) LUT6_inst8563 (
   .O(to_level3[787]),
   .I0(level4_in[4722]),
   .I1(level4_in[4723]),
   .I2(level4_in[4724]),
   .I3(level4_in[4725]),
   .I4(level4_in[4726]),
   .I5(level4_in[4727])
);

LUT6 #(
   .INIT(64'hddb208afddb208af)  
) LUT6_inst8564 (
   .O(to_level3[788]),
   .I0(level4_in[4728]),
   .I1(level4_in[4729]),
   .I2(level4_in[4730]),
   .I3(level4_in[4731]),
   .I4(level4_in[4732]),
   .I5(level4_in[4733])
);

LUT6 #(
   .INIT(64'h7c51e7f17c51e7f1)  
) LUT6_inst8565 (
   .O(to_level3[789]),
   .I0(level4_in[4734]),
   .I1(level4_in[4735]),
   .I2(level4_in[4736]),
   .I3(level4_in[4737]),
   .I4(level4_in[4738]),
   .I5(level4_in[4739])
);

LUT6 #(
   .INIT(64'hc015f1b0c015f1b0)  
) LUT6_inst8566 (
   .O(to_level3[790]),
   .I0(level4_in[4740]),
   .I1(level4_in[4741]),
   .I2(level4_in[4742]),
   .I3(level4_in[4743]),
   .I4(level4_in[4744]),
   .I5(level4_in[4745])
);

LUT6 #(
   .INIT(64'h2292fe372292fe37)  
) LUT6_inst8567 (
   .O(to_level3[791]),
   .I0(level4_in[4746]),
   .I1(level4_in[4747]),
   .I2(level4_in[4748]),
   .I3(level4_in[4749]),
   .I4(level4_in[4750]),
   .I5(level4_in[4751])
);

LUT6 #(
   .INIT(64'h2b99a4a62b99a4a6)  
) LUT6_inst8568 (
   .O(to_level3[792]),
   .I0(level4_in[4752]),
   .I1(level4_in[4753]),
   .I2(level4_in[4754]),
   .I3(level4_in[4755]),
   .I4(level4_in[4756]),
   .I5(level4_in[4757])
);

LUT6 #(
   .INIT(64'hc480c384c480c384)  
) LUT6_inst8569 (
   .O(to_level3[793]),
   .I0(level4_in[4758]),
   .I1(level4_in[4759]),
   .I2(level4_in[4760]),
   .I3(level4_in[4761]),
   .I4(level4_in[4762]),
   .I5(level4_in[4763])
);

LUT6 #(
   .INIT(64'hcffed1e4cffed1e4)  
) LUT6_inst8570 (
   .O(to_level3[794]),
   .I0(level4_in[4764]),
   .I1(level4_in[4765]),
   .I2(level4_in[4766]),
   .I3(level4_in[4767]),
   .I4(level4_in[4768]),
   .I5(level4_in[4769])
);

LUT6 #(
   .INIT(64'h55ae5e6055ae5e60)  
) LUT6_inst8571 (
   .O(to_level3[795]),
   .I0(level4_in[4770]),
   .I1(level4_in[4771]),
   .I2(level4_in[4772]),
   .I3(level4_in[4773]),
   .I4(level4_in[4774]),
   .I5(level4_in[4775])
);

LUT6 #(
   .INIT(64'h2169b78e2169b78e)  
) LUT6_inst8572 (
   .O(to_level3[796]),
   .I0(level4_in[4776]),
   .I1(level4_in[4777]),
   .I2(level4_in[4778]),
   .I3(level4_in[4779]),
   .I4(level4_in[4780]),
   .I5(level4_in[4781])
);

LUT6 #(
   .INIT(64'h4adde7cf4adde7cf)  
) LUT6_inst8573 (
   .O(to_level3[797]),
   .I0(level4_in[4782]),
   .I1(level4_in[4783]),
   .I2(level4_in[4784]),
   .I3(level4_in[4785]),
   .I4(level4_in[4786]),
   .I5(level4_in[4787])
);

LUT6 #(
   .INIT(64'h5cdca3565cdca356)  
) LUT6_inst8574 (
   .O(to_level3[798]),
   .I0(level4_in[4788]),
   .I1(level4_in[4789]),
   .I2(level4_in[4790]),
   .I3(level4_in[4791]),
   .I4(level4_in[4792]),
   .I5(level4_in[4793])
);

LUT6 #(
   .INIT(64'hc4eb2ea2c4eb2ea2)  
) LUT6_inst8575 (
   .O(to_level3[799]),
   .I0(level4_in[4794]),
   .I1(level4_in[4795]),
   .I2(level4_in[4796]),
   .I3(level4_in[4797]),
   .I4(level4_in[4798]),
   .I5(level4_in[4799])
);

LUT6 #(
   .INIT(64'h2421b8142421b814)  
) LUT6_inst8576 (
   .O(to_level3[800]),
   .I0(level4_in[4800]),
   .I1(level4_in[4801]),
   .I2(level4_in[4802]),
   .I3(level4_in[4803]),
   .I4(level4_in[4804]),
   .I5(level4_in[4805])
);

LUT6 #(
   .INIT(64'hd15797a9d15797a9)  
) LUT6_inst8577 (
   .O(to_level3[801]),
   .I0(level4_in[4806]),
   .I1(level4_in[4807]),
   .I2(level4_in[4808]),
   .I3(level4_in[4809]),
   .I4(level4_in[4810]),
   .I5(level4_in[4811])
);

LUT6 #(
   .INIT(64'h5323a85e5323a85e)  
) LUT6_inst8578 (
   .O(to_level3[802]),
   .I0(level4_in[4812]),
   .I1(level4_in[4813]),
   .I2(level4_in[4814]),
   .I3(level4_in[4815]),
   .I4(level4_in[4816]),
   .I5(level4_in[4817])
);

LUT6 #(
   .INIT(64'h601621d7601621d7)  
) LUT6_inst8579 (
   .O(to_level3[803]),
   .I0(level4_in[4818]),
   .I1(level4_in[4819]),
   .I2(level4_in[4820]),
   .I3(level4_in[4821]),
   .I4(level4_in[4822]),
   .I5(level4_in[4823])
);

LUT6 #(
   .INIT(64'ha38b0007a38b0007)  
) LUT6_inst8580 (
   .O(to_level3[804]),
   .I0(level4_in[4824]),
   .I1(level4_in[4825]),
   .I2(level4_in[4826]),
   .I3(level4_in[4827]),
   .I4(level4_in[4828]),
   .I5(level4_in[4829])
);

LUT6 #(
   .INIT(64'h9bacd30e9bacd30e)  
) LUT6_inst8581 (
   .O(to_level3[805]),
   .I0(level4_in[4830]),
   .I1(level4_in[4831]),
   .I2(level4_in[4832]),
   .I3(level4_in[4833]),
   .I4(level4_in[4834]),
   .I5(level4_in[4835])
);

LUT6 #(
   .INIT(64'hd6751015d6751015)  
) LUT6_inst8582 (
   .O(to_level3[806]),
   .I0(level4_in[4836]),
   .I1(level4_in[4837]),
   .I2(level4_in[4838]),
   .I3(level4_in[4839]),
   .I4(level4_in[4840]),
   .I5(level4_in[4841])
);

LUT6 #(
   .INIT(64'h846997cc846997cc)  
) LUT6_inst8583 (
   .O(to_level3[807]),
   .I0(level4_in[4842]),
   .I1(level4_in[4843]),
   .I2(level4_in[4844]),
   .I3(level4_in[4845]),
   .I4(level4_in[4846]),
   .I5(level4_in[4847])
);

LUT6 #(
   .INIT(64'h246e67fd246e67fd)  
) LUT6_inst8584 (
   .O(to_level3[808]),
   .I0(level4_in[4848]),
   .I1(level4_in[4849]),
   .I2(level4_in[4850]),
   .I3(level4_in[4851]),
   .I4(level4_in[4852]),
   .I5(level4_in[4853])
);

LUT6 #(
   .INIT(64'hcd927090cd927090)  
) LUT6_inst8585 (
   .O(to_level3[809]),
   .I0(level4_in[4854]),
   .I1(level4_in[4855]),
   .I2(level4_in[4856]),
   .I3(level4_in[4857]),
   .I4(level4_in[4858]),
   .I5(level4_in[4859])
);

LUT6 #(
   .INIT(64'h001d9bac001d9bac)  
) LUT6_inst8586 (
   .O(to_level3[810]),
   .I0(level4_in[4860]),
   .I1(level4_in[4861]),
   .I2(level4_in[4862]),
   .I3(level4_in[4863]),
   .I4(level4_in[4864]),
   .I5(level4_in[4865])
);

LUT6 #(
   .INIT(64'h548ba615548ba615)  
) LUT6_inst8587 (
   .O(to_level3[811]),
   .I0(level4_in[4866]),
   .I1(level4_in[4867]),
   .I2(level4_in[4868]),
   .I3(level4_in[4869]),
   .I4(level4_in[4870]),
   .I5(level4_in[4871])
);

LUT6 #(
   .INIT(64'h770e8690770e8690)  
) LUT6_inst8588 (
   .O(to_level3[812]),
   .I0(level4_in[4872]),
   .I1(level4_in[4873]),
   .I2(level4_in[4874]),
   .I3(level4_in[4875]),
   .I4(level4_in[4876]),
   .I5(level4_in[4877])
);

LUT6 #(
   .INIT(64'hd880b011d880b011)  
) LUT6_inst8589 (
   .O(to_level3[813]),
   .I0(level4_in[4878]),
   .I1(level4_in[4879]),
   .I2(level4_in[4880]),
   .I3(level4_in[4881]),
   .I4(level4_in[4882]),
   .I5(level4_in[4883])
);

LUT6 #(
   .INIT(64'h36788c0636788c06)  
) LUT6_inst8590 (
   .O(to_level3[814]),
   .I0(level4_in[4884]),
   .I1(level4_in[4885]),
   .I2(level4_in[4886]),
   .I3(level4_in[4887]),
   .I4(level4_in[4888]),
   .I5(level4_in[4889])
);

LUT6 #(
   .INIT(64'h7b6fdf897b6fdf89)  
) LUT6_inst8591 (
   .O(to_level3[815]),
   .I0(level4_in[4890]),
   .I1(level4_in[4891]),
   .I2(level4_in[4892]),
   .I3(level4_in[4893]),
   .I4(level4_in[4894]),
   .I5(level4_in[4895])
);

LUT6 #(
   .INIT(64'h954b872f954b872f)  
) LUT6_inst8592 (
   .O(to_level3[816]),
   .I0(level4_in[4896]),
   .I1(level4_in[4897]),
   .I2(level4_in[4898]),
   .I3(level4_in[4899]),
   .I4(level4_in[4900]),
   .I5(level4_in[4901])
);

LUT6 #(
   .INIT(64'h5325a6fd5325a6fd)  
) LUT6_inst8593 (
   .O(to_level3[817]),
   .I0(level4_in[4902]),
   .I1(level4_in[4903]),
   .I2(level4_in[4904]),
   .I3(level4_in[4905]),
   .I4(level4_in[4906]),
   .I5(level4_in[4907])
);

LUT6 #(
   .INIT(64'he38a032ce38a032c)  
) LUT6_inst8594 (
   .O(to_level3[818]),
   .I0(level4_in[4908]),
   .I1(level4_in[4909]),
   .I2(level4_in[4910]),
   .I3(level4_in[4911]),
   .I4(level4_in[4912]),
   .I5(level4_in[4913])
);

LUT6 #(
   .INIT(64'h8d7597638d759763)  
) LUT6_inst8595 (
   .O(to_level3[819]),
   .I0(level4_in[4914]),
   .I1(level4_in[4915]),
   .I2(level4_in[4916]),
   .I3(level4_in[4917]),
   .I4(level4_in[4918]),
   .I5(level4_in[4919])
);

LUT6 #(
   .INIT(64'h7d42543b7d42543b)  
) LUT6_inst8596 (
   .O(to_level3[820]),
   .I0(level4_in[4920]),
   .I1(level4_in[4921]),
   .I2(level4_in[4922]),
   .I3(level4_in[4923]),
   .I4(level4_in[4924]),
   .I5(level4_in[4925])
);

LUT6 #(
   .INIT(64'h00a1e8b000a1e8b0)  
) LUT6_inst8597 (
   .O(to_level3[821]),
   .I0(level4_in[4926]),
   .I1(level4_in[4927]),
   .I2(level4_in[4928]),
   .I3(level4_in[4929]),
   .I4(level4_in[4930]),
   .I5(level4_in[4931])
);

LUT6 #(
   .INIT(64'hbcb7c3dbbcb7c3db)  
) LUT6_inst8598 (
   .O(to_level3[822]),
   .I0(level4_in[4932]),
   .I1(level4_in[4933]),
   .I2(level4_in[4934]),
   .I3(level4_in[4935]),
   .I4(level4_in[4936]),
   .I5(level4_in[4937])
);

LUT6 #(
   .INIT(64'h49a7e24349a7e243)  
) LUT6_inst8599 (
   .O(to_level3[823]),
   .I0(level4_in[4938]),
   .I1(level4_in[4939]),
   .I2(level4_in[4940]),
   .I3(level4_in[4941]),
   .I4(level4_in[4942]),
   .I5(level4_in[4943])
);

LUT6 #(
   .INIT(64'h598c78ec598c78ec)  
) LUT6_inst8600 (
   .O(to_level3[824]),
   .I0(level4_in[4944]),
   .I1(level4_in[4945]),
   .I2(level4_in[4946]),
   .I3(level4_in[4947]),
   .I4(level4_in[4948]),
   .I5(level4_in[4949])
);

LUT6 #(
   .INIT(64'hd77cd9bdd77cd9bd)  
) LUT6_inst8601 (
   .O(to_level3[825]),
   .I0(level4_in[4950]),
   .I1(level4_in[4951]),
   .I2(level4_in[4952]),
   .I3(level4_in[4953]),
   .I4(level4_in[4954]),
   .I5(level4_in[4955])
);

LUT6 #(
   .INIT(64'h7ebe00c47ebe00c4)  
) LUT6_inst8602 (
   .O(to_level3[826]),
   .I0(level4_in[4956]),
   .I1(level4_in[4957]),
   .I2(level4_in[4958]),
   .I3(level4_in[4959]),
   .I4(level4_in[4960]),
   .I5(level4_in[4961])
);

LUT6 #(
   .INIT(64'hc210567ec210567e)  
) LUT6_inst8603 (
   .O(to_level3[827]),
   .I0(level4_in[4962]),
   .I1(level4_in[4963]),
   .I2(level4_in[4964]),
   .I3(level4_in[4965]),
   .I4(level4_in[4966]),
   .I5(level4_in[4967])
);

LUT6 #(
   .INIT(64'hbb0e2d6ebb0e2d6e)  
) LUT6_inst8604 (
   .O(to_level3[828]),
   .I0(level4_in[4968]),
   .I1(level4_in[4969]),
   .I2(level4_in[4970]),
   .I3(level4_in[4971]),
   .I4(level4_in[4972]),
   .I5(level4_in[4973])
);

LUT6 #(
   .INIT(64'hc99f604bc99f604b)  
) LUT6_inst8605 (
   .O(to_level3[829]),
   .I0(level4_in[4974]),
   .I1(level4_in[4975]),
   .I2(level4_in[4976]),
   .I3(level4_in[4977]),
   .I4(level4_in[4978]),
   .I5(level4_in[4979])
);

LUT6 #(
   .INIT(64'h30cbec9e30cbec9e)  
) LUT6_inst8606 (
   .O(to_level3[830]),
   .I0(level4_in[4980]),
   .I1(level4_in[4981]),
   .I2(level4_in[4982]),
   .I3(level4_in[4983]),
   .I4(level4_in[4984]),
   .I5(level4_in[4985])
);

LUT6 #(
   .INIT(64'h2864571d2864571d)  
) LUT6_inst8607 (
   .O(to_level3[831]),
   .I0(level4_in[4986]),
   .I1(level4_in[4987]),
   .I2(level4_in[4988]),
   .I3(level4_in[4989]),
   .I4(level4_in[4990]),
   .I5(level4_in[4991])
);

LUT6 #(
   .INIT(64'hfb2b2fd1fb2b2fd1)  
) LUT6_inst8608 (
   .O(to_level3[832]),
   .I0(level4_in[4992]),
   .I1(level4_in[4993]),
   .I2(level4_in[4994]),
   .I3(level4_in[4995]),
   .I4(level4_in[4996]),
   .I5(level4_in[4997])
);

LUT6 #(
   .INIT(64'h025c2186025c2186)  
) LUT6_inst8609 (
   .O(to_level3[833]),
   .I0(level4_in[4998]),
   .I1(level4_in[4999]),
   .I2(level4_in[5000]),
   .I3(level4_in[5001]),
   .I4(level4_in[5002]),
   .I5(level4_in[5003])
);

LUT6 #(
   .INIT(64'hff671bd2ff671bd2)  
) LUT6_inst8610 (
   .O(to_level3[834]),
   .I0(level4_in[5004]),
   .I1(level4_in[5005]),
   .I2(level4_in[5006]),
   .I3(level4_in[5007]),
   .I4(level4_in[5008]),
   .I5(level4_in[5009])
);

LUT6 #(
   .INIT(64'h90b5bd6e90b5bd6e)  
) LUT6_inst8611 (
   .O(to_level3[835]),
   .I0(level4_in[5010]),
   .I1(level4_in[5011]),
   .I2(level4_in[5012]),
   .I3(level4_in[5013]),
   .I4(level4_in[5014]),
   .I5(level4_in[5015])
);

LUT6 #(
   .INIT(64'hfeb2fb3afeb2fb3a)  
) LUT6_inst8612 (
   .O(to_level3[836]),
   .I0(level4_in[5016]),
   .I1(level4_in[5017]),
   .I2(level4_in[5018]),
   .I3(level4_in[5019]),
   .I4(level4_in[5020]),
   .I5(level4_in[5021])
);

LUT6 #(
   .INIT(64'h0483838d0483838d)  
) LUT6_inst8613 (
   .O(to_level3[837]),
   .I0(level4_in[5022]),
   .I1(level4_in[5023]),
   .I2(level4_in[5024]),
   .I3(level4_in[5025]),
   .I4(level4_in[5026]),
   .I5(level4_in[5027])
);

LUT6 #(
   .INIT(64'h0397d1e10397d1e1)  
) LUT6_inst8614 (
   .O(to_level3[838]),
   .I0(level4_in[5028]),
   .I1(level4_in[5029]),
   .I2(level4_in[5030]),
   .I3(level4_in[5031]),
   .I4(level4_in[5032]),
   .I5(level4_in[5033])
);

LUT6 #(
   .INIT(64'ha9802c62a9802c62)  
) LUT6_inst8615 (
   .O(to_level3[839]),
   .I0(level4_in[5034]),
   .I1(level4_in[5035]),
   .I2(level4_in[5036]),
   .I3(level4_in[5037]),
   .I4(level4_in[5038]),
   .I5(level4_in[5039])
);

LUT6 #(
   .INIT(64'h6dcecc516dcecc51)  
) LUT6_inst8616 (
   .O(to_level3[840]),
   .I0(level4_in[5040]),
   .I1(level4_in[5041]),
   .I2(level4_in[5042]),
   .I3(level4_in[5043]),
   .I4(level4_in[5044]),
   .I5(level4_in[5045])
);

LUT6 #(
   .INIT(64'h39405c5439405c54)  
) LUT6_inst8617 (
   .O(to_level3[841]),
   .I0(level4_in[5046]),
   .I1(level4_in[5047]),
   .I2(level4_in[5048]),
   .I3(level4_in[5049]),
   .I4(level4_in[5050]),
   .I5(level4_in[5051])
);

LUT6 #(
   .INIT(64'hcabb244ccabb244c)  
) LUT6_inst8618 (
   .O(to_level3[842]),
   .I0(level4_in[5052]),
   .I1(level4_in[5053]),
   .I2(level4_in[5054]),
   .I3(level4_in[5055]),
   .I4(level4_in[5056]),
   .I5(level4_in[5057])
);

LUT6 #(
   .INIT(64'hdb91fcf1db91fcf1)  
) LUT6_inst8619 (
   .O(to_level3[843]),
   .I0(level4_in[5058]),
   .I1(level4_in[5059]),
   .I2(level4_in[5060]),
   .I3(level4_in[5061]),
   .I4(level4_in[5062]),
   .I5(level4_in[5063])
);

LUT6 #(
   .INIT(64'h6d1571166d157116)  
) LUT6_inst8620 (
   .O(to_level3[844]),
   .I0(level4_in[5064]),
   .I1(level4_in[5065]),
   .I2(level4_in[5066]),
   .I3(level4_in[5067]),
   .I4(level4_in[5068]),
   .I5(level4_in[5069])
);

LUT6 #(
   .INIT(64'h463d34d4463d34d4)  
) LUT6_inst8621 (
   .O(to_level3[845]),
   .I0(level4_in[5070]),
   .I1(level4_in[5071]),
   .I2(level4_in[5072]),
   .I3(level4_in[5073]),
   .I4(level4_in[5074]),
   .I5(level4_in[5075])
);

LUT6 #(
   .INIT(64'hfc92b80dfc92b80d)  
) LUT6_inst8622 (
   .O(to_level3[846]),
   .I0(level4_in[5076]),
   .I1(level4_in[5077]),
   .I2(level4_in[5078]),
   .I3(level4_in[5079]),
   .I4(level4_in[5080]),
   .I5(level4_in[5081])
);

LUT6 #(
   .INIT(64'hf53ef506f53ef506)  
) LUT6_inst8623 (
   .O(to_level3[847]),
   .I0(level4_in[5082]),
   .I1(level4_in[5083]),
   .I2(level4_in[5084]),
   .I3(level4_in[5085]),
   .I4(level4_in[5086]),
   .I5(level4_in[5087])
);

LUT6 #(
   .INIT(64'h188e6619188e6619)  
) LUT6_inst8624 (
   .O(to_level3[848]),
   .I0(level4_in[5088]),
   .I1(level4_in[5089]),
   .I2(level4_in[5090]),
   .I3(level4_in[5091]),
   .I4(level4_in[5092]),
   .I5(level4_in[5093])
);

LUT6 #(
   .INIT(64'h172e73dc172e73dc)  
) LUT6_inst8625 (
   .O(to_level3[849]),
   .I0(level4_in[5094]),
   .I1(level4_in[5095]),
   .I2(level4_in[5096]),
   .I3(level4_in[5097]),
   .I4(level4_in[5098]),
   .I5(level4_in[5099])
);

LUT6 #(
   .INIT(64'h2967b4602967b460)  
) LUT6_inst8626 (
   .O(to_level3[850]),
   .I0(level4_in[5100]),
   .I1(level4_in[5101]),
   .I2(level4_in[5102]),
   .I3(level4_in[5103]),
   .I4(level4_in[5104]),
   .I5(level4_in[5105])
);

LUT6 #(
   .INIT(64'he01bdf50e01bdf50)  
) LUT6_inst8627 (
   .O(to_level3[851]),
   .I0(level4_in[5106]),
   .I1(level4_in[5107]),
   .I2(level4_in[5108]),
   .I3(level4_in[5109]),
   .I4(level4_in[5110]),
   .I5(level4_in[5111])
);

LUT6 #(
   .INIT(64'hc597b902c597b902)  
) LUT6_inst8628 (
   .O(to_level3[852]),
   .I0(level4_in[5112]),
   .I1(level4_in[5113]),
   .I2(level4_in[5114]),
   .I3(level4_in[5115]),
   .I4(level4_in[5116]),
   .I5(level4_in[5117])
);

LUT6 #(
   .INIT(64'h90a5f10b90a5f10b)  
) LUT6_inst8629 (
   .O(to_level3[853]),
   .I0(level4_in[5118]),
   .I1(level4_in[5119]),
   .I2(level4_in[5120]),
   .I3(level4_in[5121]),
   .I4(level4_in[5122]),
   .I5(level4_in[5123])
);

LUT6 #(
   .INIT(64'h6cc03e756cc03e75)  
) LUT6_inst8630 (
   .O(to_level3[854]),
   .I0(level4_in[5124]),
   .I1(level4_in[5125]),
   .I2(level4_in[5126]),
   .I3(level4_in[5127]),
   .I4(level4_in[5128]),
   .I5(level4_in[5129])
);

LUT6 #(
   .INIT(64'hbd58c182bd58c182)  
) LUT6_inst8631 (
   .O(to_level3[855]),
   .I0(level4_in[5130]),
   .I1(level4_in[5131]),
   .I2(level4_in[5132]),
   .I3(level4_in[5133]),
   .I4(level4_in[5134]),
   .I5(level4_in[5135])
);

LUT6 #(
   .INIT(64'he0ff3a6de0ff3a6d)  
) LUT6_inst8632 (
   .O(to_level3[856]),
   .I0(level4_in[5136]),
   .I1(level4_in[5137]),
   .I2(level4_in[5138]),
   .I3(level4_in[5139]),
   .I4(level4_in[5140]),
   .I5(level4_in[5141])
);

LUT6 #(
   .INIT(64'hff61550aff61550a)  
) LUT6_inst8633 (
   .O(to_level3[857]),
   .I0(level4_in[5142]),
   .I1(level4_in[5143]),
   .I2(level4_in[5144]),
   .I3(level4_in[5145]),
   .I4(level4_in[5146]),
   .I5(level4_in[5147])
);

LUT6 #(
   .INIT(64'ha3b0cd23a3b0cd23)  
) LUT6_inst8634 (
   .O(to_level3[858]),
   .I0(level4_in[5148]),
   .I1(level4_in[5149]),
   .I2(level4_in[5150]),
   .I3(level4_in[5151]),
   .I4(level4_in[5152]),
   .I5(level4_in[5153])
);

LUT6 #(
   .INIT(64'ha651b627a651b627)  
) LUT6_inst8635 (
   .O(to_level3[859]),
   .I0(level4_in[5154]),
   .I1(level4_in[5155]),
   .I2(level4_in[5156]),
   .I3(level4_in[5157]),
   .I4(level4_in[5158]),
   .I5(level4_in[5159])
);

LUT6 #(
   .INIT(64'h3eff57973eff5797)  
) LUT6_inst8636 (
   .O(to_level3[860]),
   .I0(level4_in[5160]),
   .I1(level4_in[5161]),
   .I2(level4_in[5162]),
   .I3(level4_in[5163]),
   .I4(level4_in[5164]),
   .I5(level4_in[5165])
);

LUT6 #(
   .INIT(64'h78adbb6378adbb63)  
) LUT6_inst8637 (
   .O(to_level3[861]),
   .I0(level4_in[5166]),
   .I1(level4_in[5167]),
   .I2(level4_in[5168]),
   .I3(level4_in[5169]),
   .I4(level4_in[5170]),
   .I5(level4_in[5171])
);

LUT6 #(
   .INIT(64'h2a98b7632a98b763)  
) LUT6_inst8638 (
   .O(to_level3[862]),
   .I0(level4_in[5172]),
   .I1(level4_in[5173]),
   .I2(level4_in[5174]),
   .I3(level4_in[5175]),
   .I4(level4_in[5176]),
   .I5(level4_in[5177])
);

LUT6 #(
   .INIT(64'h0b1036bb0b1036bb)  
) LUT6_inst8639 (
   .O(to_level3[863]),
   .I0(level4_in[5178]),
   .I1(level4_in[5179]),
   .I2(level4_in[5180]),
   .I3(level4_in[5181]),
   .I4(level4_in[5182]),
   .I5(level4_in[5183])
);

LUT6 #(
   .INIT(64'h7e3d30f77e3d30f7)  
) LUT6_inst8640 (
   .O(to_level3[864]),
   .I0(level4_in[5184]),
   .I1(level4_in[5185]),
   .I2(level4_in[5186]),
   .I3(level4_in[5187]),
   .I4(level4_in[5188]),
   .I5(level4_in[5189])
);

LUT6 #(
   .INIT(64'h9beffb859beffb85)  
) LUT6_inst8641 (
   .O(to_level3[865]),
   .I0(level4_in[5190]),
   .I1(level4_in[5191]),
   .I2(level4_in[5192]),
   .I3(level4_in[5193]),
   .I4(level4_in[5194]),
   .I5(level4_in[5195])
);

LUT6 #(
   .INIT(64'h3354d5e43354d5e4)  
) LUT6_inst8642 (
   .O(to_level3[866]),
   .I0(level4_in[5196]),
   .I1(level4_in[5197]),
   .I2(level4_in[5198]),
   .I3(level4_in[5199]),
   .I4(level4_in[5200]),
   .I5(level4_in[5201])
);

LUT6 #(
   .INIT(64'h78d96baf78d96baf)  
) LUT6_inst8643 (
   .O(to_level3[867]),
   .I0(level4_in[5202]),
   .I1(level4_in[5203]),
   .I2(level4_in[5204]),
   .I3(level4_in[5205]),
   .I4(level4_in[5206]),
   .I5(level4_in[5207])
);

LUT6 #(
   .INIT(64'h85ac85c585ac85c5)  
) LUT6_inst8644 (
   .O(to_level3[868]),
   .I0(level4_in[5208]),
   .I1(level4_in[5209]),
   .I2(level4_in[5210]),
   .I3(level4_in[5211]),
   .I4(level4_in[5212]),
   .I5(level4_in[5213])
);

LUT6 #(
   .INIT(64'hfe4ccfb4fe4ccfb4)  
) LUT6_inst8645 (
   .O(to_level3[869]),
   .I0(level4_in[5214]),
   .I1(level4_in[5215]),
   .I2(level4_in[5216]),
   .I3(level4_in[5217]),
   .I4(level4_in[5218]),
   .I5(level4_in[5219])
);

LUT6 #(
   .INIT(64'h881dd069881dd069)  
) LUT6_inst8646 (
   .O(to_level3[870]),
   .I0(level4_in[5220]),
   .I1(level4_in[5221]),
   .I2(level4_in[5222]),
   .I3(level4_in[5223]),
   .I4(level4_in[5224]),
   .I5(level4_in[5225])
);

LUT6 #(
   .INIT(64'h9040302a9040302a)  
) LUT6_inst8647 (
   .O(to_level3[871]),
   .I0(level4_in[5226]),
   .I1(level4_in[5227]),
   .I2(level4_in[5228]),
   .I3(level4_in[5229]),
   .I4(level4_in[5230]),
   .I5(level4_in[5231])
);

LUT6 #(
   .INIT(64'h94cca61d94cca61d)  
) LUT6_inst8648 (
   .O(to_level3[872]),
   .I0(level4_in[5232]),
   .I1(level4_in[5233]),
   .I2(level4_in[5234]),
   .I3(level4_in[5235]),
   .I4(level4_in[5236]),
   .I5(level4_in[5237])
);

LUT6 #(
   .INIT(64'h4014334940143349)  
) LUT6_inst8649 (
   .O(to_level3[873]),
   .I0(level4_in[5238]),
   .I1(level4_in[5239]),
   .I2(level4_in[5240]),
   .I3(level4_in[5241]),
   .I4(level4_in[5242]),
   .I5(level4_in[5243])
);

LUT6 #(
   .INIT(64'h9d88ef789d88ef78)  
) LUT6_inst8650 (
   .O(to_level3[874]),
   .I0(level4_in[5244]),
   .I1(level4_in[5245]),
   .I2(level4_in[5246]),
   .I3(level4_in[5247]),
   .I4(level4_in[5248]),
   .I5(level4_in[5249])
);

LUT6 #(
   .INIT(64'h4d9320864d932086)  
) LUT6_inst8651 (
   .O(to_level3[875]),
   .I0(level4_in[5250]),
   .I1(level4_in[5251]),
   .I2(level4_in[5252]),
   .I3(level4_in[5253]),
   .I4(level4_in[5254]),
   .I5(level4_in[5255])
);

LUT6 #(
   .INIT(64'hd177c5f2d177c5f2)  
) LUT6_inst8652 (
   .O(to_level3[876]),
   .I0(level4_in[5256]),
   .I1(level4_in[5257]),
   .I2(level4_in[5258]),
   .I3(level4_in[5259]),
   .I4(level4_in[5260]),
   .I5(level4_in[5261])
);

LUT6 #(
   .INIT(64'h8923216f8923216f)  
) LUT6_inst8653 (
   .O(to_level3[877]),
   .I0(level4_in[5262]),
   .I1(level4_in[5263]),
   .I2(level4_in[5264]),
   .I3(level4_in[5265]),
   .I4(level4_in[5266]),
   .I5(level4_in[5267])
);

LUT6 #(
   .INIT(64'h5da8edaf5da8edaf)  
) LUT6_inst8654 (
   .O(to_level3[878]),
   .I0(level4_in[5268]),
   .I1(level4_in[5269]),
   .I2(level4_in[5270]),
   .I3(level4_in[5271]),
   .I4(level4_in[5272]),
   .I5(level4_in[5273])
);

LUT6 #(
   .INIT(64'h844c66c3844c66c3)  
) LUT6_inst8655 (
   .O(to_level3[879]),
   .I0(level4_in[5274]),
   .I1(level4_in[5275]),
   .I2(level4_in[5276]),
   .I3(level4_in[5277]),
   .I4(level4_in[5278]),
   .I5(level4_in[5279])
);

LUT6 #(
   .INIT(64'hcce5737acce5737a)  
) LUT6_inst8656 (
   .O(to_level3[880]),
   .I0(level4_in[5280]),
   .I1(level4_in[5281]),
   .I2(level4_in[5282]),
   .I3(level4_in[5283]),
   .I4(level4_in[5284]),
   .I5(level4_in[5285])
);

LUT6 #(
   .INIT(64'hc8c315fac8c315fa)  
) LUT6_inst8657 (
   .O(to_level3[881]),
   .I0(level4_in[5286]),
   .I1(level4_in[5287]),
   .I2(level4_in[5288]),
   .I3(level4_in[5289]),
   .I4(level4_in[5290]),
   .I5(level4_in[5291])
);

LUT6 #(
   .INIT(64'hcdfa535ecdfa535e)  
) LUT6_inst8658 (
   .O(to_level3[882]),
   .I0(level4_in[5292]),
   .I1(level4_in[5293]),
   .I2(level4_in[5294]),
   .I3(level4_in[5295]),
   .I4(level4_in[5296]),
   .I5(level4_in[5297])
);

LUT6 #(
   .INIT(64'h8134def38134def3)  
) LUT6_inst8659 (
   .O(to_level3[883]),
   .I0(level4_in[5298]),
   .I1(level4_in[5299]),
   .I2(level4_in[5300]),
   .I3(level4_in[5301]),
   .I4(level4_in[5302]),
   .I5(level4_in[5303])
);

LUT6 #(
   .INIT(64'hefbd3250efbd3250)  
) LUT6_inst8660 (
   .O(to_level3[884]),
   .I0(level4_in[5304]),
   .I1(level4_in[5305]),
   .I2(level4_in[5306]),
   .I3(level4_in[5307]),
   .I4(level4_in[5308]),
   .I5(level4_in[5309])
);

LUT6 #(
   .INIT(64'h379a3b2e379a3b2e)  
) LUT6_inst8661 (
   .O(to_level3[885]),
   .I0(level4_in[5310]),
   .I1(level4_in[5311]),
   .I2(level4_in[5312]),
   .I3(level4_in[5313]),
   .I4(level4_in[5314]),
   .I5(level4_in[5315])
);

LUT6 #(
   .INIT(64'hf94a8bc9f94a8bc9)  
) LUT6_inst8662 (
   .O(to_level3[886]),
   .I0(level4_in[5316]),
   .I1(level4_in[5317]),
   .I2(level4_in[5318]),
   .I3(level4_in[5319]),
   .I4(level4_in[5320]),
   .I5(level4_in[5321])
);

LUT6 #(
   .INIT(64'h89cdd5f089cdd5f0)  
) LUT6_inst8663 (
   .O(to_level3[887]),
   .I0(level4_in[5322]),
   .I1(level4_in[5323]),
   .I2(level4_in[5324]),
   .I3(level4_in[5325]),
   .I4(level4_in[5326]),
   .I5(level4_in[5327])
);

LUT6 #(
   .INIT(64'h091ef662091ef662)  
) LUT6_inst8664 (
   .O(to_level3[888]),
   .I0(level4_in[5328]),
   .I1(level4_in[5329]),
   .I2(level4_in[5330]),
   .I3(level4_in[5331]),
   .I4(level4_in[5332]),
   .I5(level4_in[5333])
);

LUT6 #(
   .INIT(64'h478a51a5478a51a5)  
) LUT6_inst8665 (
   .O(to_level3[889]),
   .I0(level4_in[5334]),
   .I1(level4_in[5335]),
   .I2(level4_in[5336]),
   .I3(level4_in[5337]),
   .I4(level4_in[5338]),
   .I5(level4_in[5339])
);

LUT6 #(
   .INIT(64'h57ef414b57ef414b)  
) LUT6_inst8666 (
   .O(to_level3[890]),
   .I0(level4_in[5340]),
   .I1(level4_in[5341]),
   .I2(level4_in[5342]),
   .I3(level4_in[5343]),
   .I4(level4_in[5344]),
   .I5(level4_in[5345])
);

LUT6 #(
   .INIT(64'h0aaaa8950aaaa895)  
) LUT6_inst8667 (
   .O(to_level3[891]),
   .I0(level4_in[5346]),
   .I1(level4_in[5347]),
   .I2(level4_in[5348]),
   .I3(level4_in[5349]),
   .I4(level4_in[5350]),
   .I5(level4_in[5351])
);

LUT6 #(
   .INIT(64'he5578045e5578045)  
) LUT6_inst8668 (
   .O(to_level3[892]),
   .I0(level4_in[5352]),
   .I1(level4_in[5353]),
   .I2(level4_in[5354]),
   .I3(level4_in[5355]),
   .I4(level4_in[5356]),
   .I5(level4_in[5357])
);

LUT6 #(
   .INIT(64'h8012f3508012f350)  
) LUT6_inst8669 (
   .O(to_level3[893]),
   .I0(level4_in[5358]),
   .I1(level4_in[5359]),
   .I2(level4_in[5360]),
   .I3(level4_in[5361]),
   .I4(level4_in[5362]),
   .I5(level4_in[5363])
);

LUT6 #(
   .INIT(64'h457d1fe0457d1fe0)  
) LUT6_inst8670 (
   .O(to_level3[894]),
   .I0(level4_in[5364]),
   .I1(level4_in[5365]),
   .I2(level4_in[5366]),
   .I3(level4_in[5367]),
   .I4(level4_in[5368]),
   .I5(level4_in[5369])
);

LUT6 #(
   .INIT(64'ha80703a5a80703a5)  
) LUT6_inst8671 (
   .O(to_level3[895]),
   .I0(level4_in[5370]),
   .I1(level4_in[5371]),
   .I2(level4_in[5372]),
   .I3(level4_in[5373]),
   .I4(level4_in[5374]),
   .I5(level4_in[5375])
);

LUT6 #(
   .INIT(64'hb5611491b5611491)  
) LUT6_inst8672 (
   .O(to_level3[896]),
   .I0(level4_in[5376]),
   .I1(level4_in[5377]),
   .I2(level4_in[5378]),
   .I3(level4_in[5379]),
   .I4(level4_in[5380]),
   .I5(level4_in[5381])
);

LUT6 #(
   .INIT(64'ha72d2ed0a72d2ed0)  
) LUT6_inst8673 (
   .O(to_level3[897]),
   .I0(level4_in[5382]),
   .I1(level4_in[5383]),
   .I2(level4_in[5384]),
   .I3(level4_in[5385]),
   .I4(level4_in[5386]),
   .I5(level4_in[5387])
);

LUT6 #(
   .INIT(64'h691422bd691422bd)  
) LUT6_inst8674 (
   .O(to_level3[898]),
   .I0(level4_in[5388]),
   .I1(level4_in[5389]),
   .I2(level4_in[5390]),
   .I3(level4_in[5391]),
   .I4(level4_in[5392]),
   .I5(level4_in[5393])
);

LUT6 #(
   .INIT(64'h247d66a4247d66a4)  
) LUT6_inst8675 (
   .O(to_level3[899]),
   .I0(level4_in[5394]),
   .I1(level4_in[5395]),
   .I2(level4_in[5396]),
   .I3(level4_in[5397]),
   .I4(level4_in[5398]),
   .I5(level4_in[5399])
);

LUT6 #(
   .INIT(64'h8394b8c28394b8c2)  
) LUT6_inst8676 (
   .O(to_level3[900]),
   .I0(level4_in[5400]),
   .I1(level4_in[5401]),
   .I2(level4_in[5402]),
   .I3(level4_in[5403]),
   .I4(level4_in[5404]),
   .I5(level4_in[5405])
);

LUT6 #(
   .INIT(64'h84e2b2bf84e2b2bf)  
) LUT6_inst8677 (
   .O(to_level3[901]),
   .I0(level4_in[5406]),
   .I1(level4_in[5407]),
   .I2(level4_in[5408]),
   .I3(level4_in[5409]),
   .I4(level4_in[5410]),
   .I5(level4_in[5411])
);

LUT6 #(
   .INIT(64'h7122469771224697)  
) LUT6_inst8678 (
   .O(to_level3[902]),
   .I0(level4_in[5412]),
   .I1(level4_in[5413]),
   .I2(level4_in[5414]),
   .I3(level4_in[5415]),
   .I4(level4_in[5416]),
   .I5(level4_in[5417])
);

LUT6 #(
   .INIT(64'h83e2fe4c83e2fe4c)  
) LUT6_inst8679 (
   .O(to_level3[903]),
   .I0(level4_in[5418]),
   .I1(level4_in[5419]),
   .I2(level4_in[5420]),
   .I3(level4_in[5421]),
   .I4(level4_in[5422]),
   .I5(level4_in[5423])
);

LUT6 #(
   .INIT(64'hd2821e5bd2821e5b)  
) LUT6_inst8680 (
   .O(to_level3[904]),
   .I0(level4_in[5424]),
   .I1(level4_in[5425]),
   .I2(level4_in[5426]),
   .I3(level4_in[5427]),
   .I4(level4_in[5428]),
   .I5(level4_in[5429])
);

LUT6 #(
   .INIT(64'h2c072d982c072d98)  
) LUT6_inst8681 (
   .O(to_level3[905]),
   .I0(level4_in[5430]),
   .I1(level4_in[5431]),
   .I2(level4_in[5432]),
   .I3(level4_in[5433]),
   .I4(level4_in[5434]),
   .I5(level4_in[5435])
);

LUT6 #(
   .INIT(64'h84afe78a84afe78a)  
) LUT6_inst8682 (
   .O(to_level3[906]),
   .I0(level4_in[5436]),
   .I1(level4_in[5437]),
   .I2(level4_in[5438]),
   .I3(level4_in[5439]),
   .I4(level4_in[5440]),
   .I5(level4_in[5441])
);

LUT6 #(
   .INIT(64'hd5ba7aedd5ba7aed)  
) LUT6_inst8683 (
   .O(to_level3[907]),
   .I0(level4_in[5442]),
   .I1(level4_in[5443]),
   .I2(level4_in[5444]),
   .I3(level4_in[5445]),
   .I4(level4_in[5446]),
   .I5(level4_in[5447])
);

LUT6 #(
   .INIT(64'h0d5b8c600d5b8c60)  
) LUT6_inst8684 (
   .O(to_level3[908]),
   .I0(level4_in[5448]),
   .I1(level4_in[5449]),
   .I2(level4_in[5450]),
   .I3(level4_in[5451]),
   .I4(level4_in[5452]),
   .I5(level4_in[5453])
);

LUT6 #(
   .INIT(64'hb9ac8ebcb9ac8ebc)  
) LUT6_inst8685 (
   .O(to_level3[909]),
   .I0(level4_in[5454]),
   .I1(level4_in[5455]),
   .I2(level4_in[5456]),
   .I3(level4_in[5457]),
   .I4(level4_in[5458]),
   .I5(level4_in[5459])
);

LUT6 #(
   .INIT(64'h84d3341684d33416)  
) LUT6_inst8686 (
   .O(to_level3[910]),
   .I0(level4_in[5460]),
   .I1(level4_in[5461]),
   .I2(level4_in[5462]),
   .I3(level4_in[5463]),
   .I4(level4_in[5464]),
   .I5(level4_in[5465])
);

LUT6 #(
   .INIT(64'h62a35bd962a35bd9)  
) LUT6_inst8687 (
   .O(to_level3[911]),
   .I0(level4_in[5466]),
   .I1(level4_in[5467]),
   .I2(level4_in[5468]),
   .I3(level4_in[5469]),
   .I4(level4_in[5470]),
   .I5(level4_in[5471])
);

LUT6 #(
   .INIT(64'hda7ce95bda7ce95b)  
) LUT6_inst8688 (
   .O(to_level3[912]),
   .I0(level4_in[5472]),
   .I1(level4_in[5473]),
   .I2(level4_in[5474]),
   .I3(level4_in[5475]),
   .I4(level4_in[5476]),
   .I5(level4_in[5477])
);

LUT6 #(
   .INIT(64'h812f9571812f9571)  
) LUT6_inst8689 (
   .O(to_level3[913]),
   .I0(level4_in[5478]),
   .I1(level4_in[5479]),
   .I2(level4_in[5480]),
   .I3(level4_in[5481]),
   .I4(level4_in[5482]),
   .I5(level4_in[5483])
);

LUT6 #(
   .INIT(64'hc76e1900c76e1900)  
) LUT6_inst8690 (
   .O(to_level3[914]),
   .I0(level4_in[5484]),
   .I1(level4_in[5485]),
   .I2(level4_in[5486]),
   .I3(level4_in[5487]),
   .I4(level4_in[5488]),
   .I5(level4_in[5489])
);

LUT6 #(
   .INIT(64'h8ae8af688ae8af68)  
) LUT6_inst8691 (
   .O(to_level3[915]),
   .I0(level4_in[5490]),
   .I1(level4_in[5491]),
   .I2(level4_in[5492]),
   .I3(level4_in[5493]),
   .I4(level4_in[5494]),
   .I5(level4_in[5495])
);

LUT6 #(
   .INIT(64'h03ecf92c03ecf92c)  
) LUT6_inst8692 (
   .O(to_level3[916]),
   .I0(level4_in[5496]),
   .I1(level4_in[5497]),
   .I2(level4_in[5498]),
   .I3(level4_in[5499]),
   .I4(level4_in[5500]),
   .I5(level4_in[5501])
);

LUT6 #(
   .INIT(64'h0f78b2100f78b210)  
) LUT6_inst8693 (
   .O(to_level3[917]),
   .I0(level4_in[5502]),
   .I1(level4_in[5503]),
   .I2(level4_in[5504]),
   .I3(level4_in[5505]),
   .I4(level4_in[5506]),
   .I5(level4_in[5507])
);

LUT6 #(
   .INIT(64'haf70d5e0af70d5e0)  
) LUT6_inst8694 (
   .O(to_level3[918]),
   .I0(level4_in[5508]),
   .I1(level4_in[5509]),
   .I2(level4_in[5510]),
   .I3(level4_in[5511]),
   .I4(level4_in[5512]),
   .I5(level4_in[5513])
);

LUT6 #(
   .INIT(64'hd61318c6d61318c6)  
) LUT6_inst8695 (
   .O(to_level3[919]),
   .I0(level4_in[5514]),
   .I1(level4_in[5515]),
   .I2(level4_in[5516]),
   .I3(level4_in[5517]),
   .I4(level4_in[5518]),
   .I5(level4_in[5519])
);

LUT6 #(
   .INIT(64'hafe2e4e6afe2e4e6)  
) LUT6_inst8696 (
   .O(to_level3[920]),
   .I0(level4_in[5520]),
   .I1(level4_in[5521]),
   .I2(level4_in[5522]),
   .I3(level4_in[5523]),
   .I4(level4_in[5524]),
   .I5(level4_in[5525])
);

LUT6 #(
   .INIT(64'hf8ef0598f8ef0598)  
) LUT6_inst8697 (
   .O(to_level3[921]),
   .I0(level4_in[5526]),
   .I1(level4_in[5527]),
   .I2(level4_in[5528]),
   .I3(level4_in[5529]),
   .I4(level4_in[5530]),
   .I5(level4_in[5531])
);

LUT6 #(
   .INIT(64'hb5859734b5859734)  
) LUT6_inst8698 (
   .O(to_level3[922]),
   .I0(level4_in[5532]),
   .I1(level4_in[5533]),
   .I2(level4_in[5534]),
   .I3(level4_in[5535]),
   .I4(level4_in[5536]),
   .I5(level4_in[5537])
);

LUT6 #(
   .INIT(64'h081625e3081625e3)  
) LUT6_inst8699 (
   .O(to_level3[923]),
   .I0(level4_in[5538]),
   .I1(level4_in[5539]),
   .I2(level4_in[5540]),
   .I3(level4_in[5541]),
   .I4(level4_in[5542]),
   .I5(level4_in[5543])
);

LUT6 #(
   .INIT(64'hda3fa181da3fa181)  
) LUT6_inst8700 (
   .O(to_level3[924]),
   .I0(level4_in[5544]),
   .I1(level4_in[5545]),
   .I2(level4_in[5546]),
   .I3(level4_in[5547]),
   .I4(level4_in[5548]),
   .I5(level4_in[5549])
);

LUT6 #(
   .INIT(64'h1c17412b1c17412b)  
) LUT6_inst8701 (
   .O(to_level3[925]),
   .I0(level4_in[5550]),
   .I1(level4_in[5551]),
   .I2(level4_in[5552]),
   .I3(level4_in[5553]),
   .I4(level4_in[5554]),
   .I5(level4_in[5555])
);

LUT6 #(
   .INIT(64'hba843f4fba843f4f)  
) LUT6_inst8702 (
   .O(to_level3[926]),
   .I0(level4_in[5556]),
   .I1(level4_in[5557]),
   .I2(level4_in[5558]),
   .I3(level4_in[5559]),
   .I4(level4_in[5560]),
   .I5(level4_in[5561])
);

LUT6 #(
   .INIT(64'h0964dae60964dae6)  
) LUT6_inst8703 (
   .O(to_level3[927]),
   .I0(level4_in[5562]),
   .I1(level4_in[5563]),
   .I2(level4_in[5564]),
   .I3(level4_in[5565]),
   .I4(level4_in[5566]),
   .I5(level4_in[5567])
);

LUT6 #(
   .INIT(64'hdbe0e6c8dbe0e6c8)  
) LUT6_inst8704 (
   .O(to_level3[928]),
   .I0(level4_in[5568]),
   .I1(level4_in[5569]),
   .I2(level4_in[5570]),
   .I3(level4_in[5571]),
   .I4(level4_in[5572]),
   .I5(level4_in[5573])
);

LUT6 #(
   .INIT(64'h5f2dc6825f2dc682)  
) LUT6_inst8705 (
   .O(to_level3[929]),
   .I0(level4_in[5574]),
   .I1(level4_in[5575]),
   .I2(level4_in[5576]),
   .I3(level4_in[5577]),
   .I4(level4_in[5578]),
   .I5(level4_in[5579])
);

LUT6 #(
   .INIT(64'h7ac20b567ac20b56)  
) LUT6_inst8706 (
   .O(to_level3[930]),
   .I0(level4_in[5580]),
   .I1(level4_in[5581]),
   .I2(level4_in[5582]),
   .I3(level4_in[5583]),
   .I4(level4_in[5584]),
   .I5(level4_in[5585])
);

LUT6 #(
   .INIT(64'hccd9d7a6ccd9d7a6)  
) LUT6_inst8707 (
   .O(to_level3[931]),
   .I0(level4_in[5586]),
   .I1(level4_in[5587]),
   .I2(level4_in[5588]),
   .I3(level4_in[5589]),
   .I4(level4_in[5590]),
   .I5(level4_in[5591])
);

LUT6 #(
   .INIT(64'h1182cd7d1182cd7d)  
) LUT6_inst8708 (
   .O(to_level3[932]),
   .I0(level4_in[5592]),
   .I1(level4_in[5593]),
   .I2(level4_in[5594]),
   .I3(level4_in[5595]),
   .I4(level4_in[5596]),
   .I5(level4_in[5597])
);

LUT6 #(
   .INIT(64'he09f97a8e09f97a8)  
) LUT6_inst8709 (
   .O(to_level3[933]),
   .I0(level4_in[5598]),
   .I1(level4_in[5599]),
   .I2(level4_in[5600]),
   .I3(level4_in[5601]),
   .I4(level4_in[5602]),
   .I5(level4_in[5603])
);

LUT6 #(
   .INIT(64'h16f02db516f02db5)  
) LUT6_inst8710 (
   .O(to_level3[934]),
   .I0(level4_in[5604]),
   .I1(level4_in[5605]),
   .I2(level4_in[5606]),
   .I3(level4_in[5607]),
   .I4(level4_in[5608]),
   .I5(level4_in[5609])
);

LUT6 #(
   .INIT(64'h8c7180d48c7180d4)  
) LUT6_inst8711 (
   .O(to_level3[935]),
   .I0(level4_in[5610]),
   .I1(level4_in[5611]),
   .I2(level4_in[5612]),
   .I3(level4_in[5613]),
   .I4(level4_in[5614]),
   .I5(level4_in[5615])
);

LUT6 #(
   .INIT(64'h320a4e24320a4e24)  
) LUT6_inst8712 (
   .O(to_level3[936]),
   .I0(level4_in[5616]),
   .I1(level4_in[5617]),
   .I2(level4_in[5618]),
   .I3(level4_in[5619]),
   .I4(level4_in[5620]),
   .I5(level4_in[5621])
);

LUT6 #(
   .INIT(64'he655664ce655664c)  
) LUT6_inst8713 (
   .O(to_level3[937]),
   .I0(level4_in[5622]),
   .I1(level4_in[5623]),
   .I2(level4_in[5624]),
   .I3(level4_in[5625]),
   .I4(level4_in[5626]),
   .I5(level4_in[5627])
);

LUT6 #(
   .INIT(64'haa4b566aaa4b566a)  
) LUT6_inst8714 (
   .O(to_level3[938]),
   .I0(level4_in[5628]),
   .I1(level4_in[5629]),
   .I2(level4_in[5630]),
   .I3(level4_in[5631]),
   .I4(level4_in[5632]),
   .I5(level4_in[5633])
);

LUT6 #(
   .INIT(64'hac11f630ac11f630)  
) LUT6_inst8715 (
   .O(to_level3[939]),
   .I0(level4_in[5634]),
   .I1(level4_in[5635]),
   .I2(level4_in[5636]),
   .I3(level4_in[5637]),
   .I4(level4_in[5638]),
   .I5(level4_in[5639])
);

LUT6 #(
   .INIT(64'h0dcde1880dcde188)  
) LUT6_inst8716 (
   .O(to_level3[940]),
   .I0(level4_in[5640]),
   .I1(level4_in[5641]),
   .I2(level4_in[5642]),
   .I3(level4_in[5643]),
   .I4(level4_in[5644]),
   .I5(level4_in[5645])
);

LUT6 #(
   .INIT(64'he2b39805e2b39805)  
) LUT6_inst8717 (
   .O(to_level3[941]),
   .I0(level4_in[5646]),
   .I1(level4_in[5647]),
   .I2(level4_in[5648]),
   .I3(level4_in[5649]),
   .I4(level4_in[5650]),
   .I5(level4_in[5651])
);

LUT6 #(
   .INIT(64'h8a4ce66b8a4ce66b)  
) LUT6_inst8718 (
   .O(to_level3[942]),
   .I0(level4_in[5652]),
   .I1(level4_in[5653]),
   .I2(level4_in[5654]),
   .I3(level4_in[5655]),
   .I4(level4_in[5656]),
   .I5(level4_in[5657])
);

LUT6 #(
   .INIT(64'h989dde63989dde63)  
) LUT6_inst8719 (
   .O(to_level3[943]),
   .I0(level4_in[5658]),
   .I1(level4_in[5659]),
   .I2(level4_in[5660]),
   .I3(level4_in[5661]),
   .I4(level4_in[5662]),
   .I5(level4_in[5663])
);

LUT6 #(
   .INIT(64'h5b7bd1e75b7bd1e7)  
) LUT6_inst8720 (
   .O(to_level3[944]),
   .I0(level4_in[5664]),
   .I1(level4_in[5665]),
   .I2(level4_in[5666]),
   .I3(level4_in[5667]),
   .I4(level4_in[5668]),
   .I5(level4_in[5669])
);

LUT6 #(
   .INIT(64'h6a6b1e7b6a6b1e7b)  
) LUT6_inst8721 (
   .O(to_level3[945]),
   .I0(level4_in[5670]),
   .I1(level4_in[5671]),
   .I2(level4_in[5672]),
   .I3(level4_in[5673]),
   .I4(level4_in[5674]),
   .I5(level4_in[5675])
);

LUT6 #(
   .INIT(64'h42dcf0af42dcf0af)  
) LUT6_inst8722 (
   .O(to_level3[946]),
   .I0(level4_in[5676]),
   .I1(level4_in[5677]),
   .I2(level4_in[5678]),
   .I3(level4_in[5679]),
   .I4(level4_in[5680]),
   .I5(level4_in[5681])
);

LUT6 #(
   .INIT(64'h05636be705636be7)  
) LUT6_inst8723 (
   .O(to_level3[947]),
   .I0(level4_in[5682]),
   .I1(level4_in[5683]),
   .I2(level4_in[5684]),
   .I3(level4_in[5685]),
   .I4(level4_in[5686]),
   .I5(level4_in[5687])
);

LUT6 #(
   .INIT(64'h4d3018a34d3018a3)  
) LUT6_inst8724 (
   .O(to_level3[948]),
   .I0(level4_in[5688]),
   .I1(level4_in[5689]),
   .I2(level4_in[5690]),
   .I3(level4_in[5691]),
   .I4(level4_in[5692]),
   .I5(level4_in[5693])
);

LUT6 #(
   .INIT(64'h318baf0d318baf0d)  
) LUT6_inst8725 (
   .O(to_level3[949]),
   .I0(level4_in[5694]),
   .I1(level4_in[5695]),
   .I2(level4_in[5696]),
   .I3(level4_in[5697]),
   .I4(level4_in[5698]),
   .I5(level4_in[5699])
);

LUT6 #(
   .INIT(64'h776c25f4776c25f4)  
) LUT6_inst8726 (
   .O(to_level3[950]),
   .I0(level4_in[5700]),
   .I1(level4_in[5701]),
   .I2(level4_in[5702]),
   .I3(level4_in[5703]),
   .I4(level4_in[5704]),
   .I5(level4_in[5705])
);

LUT6 #(
   .INIT(64'hce61b31dce61b31d)  
) LUT6_inst8727 (
   .O(to_level3[951]),
   .I0(level4_in[5706]),
   .I1(level4_in[5707]),
   .I2(level4_in[5708]),
   .I3(level4_in[5709]),
   .I4(level4_in[5710]),
   .I5(level4_in[5711])
);

LUT6 #(
   .INIT(64'h1ba510241ba51024)  
) LUT6_inst8728 (
   .O(to_level3[952]),
   .I0(level4_in[5712]),
   .I1(level4_in[5713]),
   .I2(level4_in[5714]),
   .I3(level4_in[5715]),
   .I4(level4_in[5716]),
   .I5(level4_in[5717])
);

LUT6 #(
   .INIT(64'h1eac9d1c1eac9d1c)  
) LUT6_inst8729 (
   .O(to_level3[953]),
   .I0(level4_in[5718]),
   .I1(level4_in[5719]),
   .I2(level4_in[5720]),
   .I3(level4_in[5721]),
   .I4(level4_in[5722]),
   .I5(level4_in[5723])
);

LUT6 #(
   .INIT(64'he5bce91be5bce91b)  
) LUT6_inst8730 (
   .O(to_level3[954]),
   .I0(level4_in[5724]),
   .I1(level4_in[5725]),
   .I2(level4_in[5726]),
   .I3(level4_in[5727]),
   .I4(level4_in[5728]),
   .I5(level4_in[5729])
);

LUT6 #(
   .INIT(64'hdbdf694adbdf694a)  
) LUT6_inst8731 (
   .O(to_level3[955]),
   .I0(level4_in[5730]),
   .I1(level4_in[5731]),
   .I2(level4_in[5732]),
   .I3(level4_in[5733]),
   .I4(level4_in[5734]),
   .I5(level4_in[5735])
);

LUT6 #(
   .INIT(64'h27c1047527c10475)  
) LUT6_inst8732 (
   .O(to_level3[956]),
   .I0(level4_in[5736]),
   .I1(level4_in[5737]),
   .I2(level4_in[5738]),
   .I3(level4_in[5739]),
   .I4(level4_in[5740]),
   .I5(level4_in[5741])
);

LUT6 #(
   .INIT(64'h44b6c0f044b6c0f0)  
) LUT6_inst8733 (
   .O(to_level3[957]),
   .I0(level4_in[5742]),
   .I1(level4_in[5743]),
   .I2(level4_in[5744]),
   .I3(level4_in[5745]),
   .I4(level4_in[5746]),
   .I5(level4_in[5747])
);

LUT6 #(
   .INIT(64'ha4d73f9aa4d73f9a)  
) LUT6_inst8734 (
   .O(to_level3[958]),
   .I0(level4_in[5748]),
   .I1(level4_in[5749]),
   .I2(level4_in[5750]),
   .I3(level4_in[5751]),
   .I4(level4_in[5752]),
   .I5(level4_in[5753])
);

LUT6 #(
   .INIT(64'h4851c4c74851c4c7)  
) LUT6_inst8735 (
   .O(to_level3[959]),
   .I0(level4_in[5754]),
   .I1(level4_in[5755]),
   .I2(level4_in[5756]),
   .I3(level4_in[5757]),
   .I4(level4_in[5758]),
   .I5(level4_in[5759])
);

LUT6 #(
   .INIT(64'hfbd6cfb7fbd6cfb7)  
) LUT6_inst8736 (
   .O(to_level3[960]),
   .I0(level4_in[5760]),
   .I1(level4_in[5761]),
   .I2(level4_in[5762]),
   .I3(level4_in[5763]),
   .I4(level4_in[5764]),
   .I5(level4_in[5765])
);

LUT6 #(
   .INIT(64'hcd1cfbc4cd1cfbc4)  
) LUT6_inst8737 (
   .O(to_level3[961]),
   .I0(level4_in[5766]),
   .I1(level4_in[5767]),
   .I2(level4_in[5768]),
   .I3(level4_in[5769]),
   .I4(level4_in[5770]),
   .I5(level4_in[5771])
);

LUT6 #(
   .INIT(64'hb177aafbb177aafb)  
) LUT6_inst8738 (
   .O(to_level3[962]),
   .I0(level4_in[5772]),
   .I1(level4_in[5773]),
   .I2(level4_in[5774]),
   .I3(level4_in[5775]),
   .I4(level4_in[5776]),
   .I5(level4_in[5777])
);

LUT6 #(
   .INIT(64'h7cf9c9a17cf9c9a1)  
) LUT6_inst8739 (
   .O(to_level3[963]),
   .I0(level4_in[5778]),
   .I1(level4_in[5779]),
   .I2(level4_in[5780]),
   .I3(level4_in[5781]),
   .I4(level4_in[5782]),
   .I5(level4_in[5783])
);

LUT6 #(
   .INIT(64'h49b1cfde49b1cfde)  
) LUT6_inst8740 (
   .O(to_level3[964]),
   .I0(level4_in[5784]),
   .I1(level4_in[5785]),
   .I2(level4_in[5786]),
   .I3(level4_in[5787]),
   .I4(level4_in[5788]),
   .I5(level4_in[5789])
);

LUT6 #(
   .INIT(64'h1b8d66a71b8d66a7)  
) LUT6_inst8741 (
   .O(to_level3[965]),
   .I0(level4_in[5790]),
   .I1(level4_in[5791]),
   .I2(level4_in[5792]),
   .I3(level4_in[5793]),
   .I4(level4_in[5794]),
   .I5(level4_in[5795])
);

LUT6 #(
   .INIT(64'h6290b0cd6290b0cd)  
) LUT6_inst8742 (
   .O(to_level3[966]),
   .I0(level4_in[5796]),
   .I1(level4_in[5797]),
   .I2(level4_in[5798]),
   .I3(level4_in[5799]),
   .I4(level4_in[5800]),
   .I5(level4_in[5801])
);

LUT6 #(
   .INIT(64'hb6260ffab6260ffa)  
) LUT6_inst8743 (
   .O(to_level3[967]),
   .I0(level4_in[5802]),
   .I1(level4_in[5803]),
   .I2(level4_in[5804]),
   .I3(level4_in[5805]),
   .I4(level4_in[5806]),
   .I5(level4_in[5807])
);

LUT6 #(
   .INIT(64'hed8f3fc4ed8f3fc4)  
) LUT6_inst8744 (
   .O(to_level3[968]),
   .I0(level4_in[5808]),
   .I1(level4_in[5809]),
   .I2(level4_in[5810]),
   .I3(level4_in[5811]),
   .I4(level4_in[5812]),
   .I5(level4_in[5813])
);

LUT6 #(
   .INIT(64'hba17f89fba17f89f)  
) LUT6_inst8745 (
   .O(to_level3[969]),
   .I0(level4_in[5814]),
   .I1(level4_in[5815]),
   .I2(level4_in[5816]),
   .I3(level4_in[5817]),
   .I4(level4_in[5818]),
   .I5(level4_in[5819])
);

LUT6 #(
   .INIT(64'h2873454528734545)  
) LUT6_inst8746 (
   .O(to_level3[970]),
   .I0(level4_in[5820]),
   .I1(level4_in[5821]),
   .I2(level4_in[5822]),
   .I3(level4_in[5823]),
   .I4(level4_in[5824]),
   .I5(level4_in[5825])
);

LUT6 #(
   .INIT(64'hcdb2cca9cdb2cca9)  
) LUT6_inst8747 (
   .O(to_level3[971]),
   .I0(level4_in[5826]),
   .I1(level4_in[5827]),
   .I2(level4_in[5828]),
   .I3(level4_in[5829]),
   .I4(level4_in[5830]),
   .I5(level4_in[5831])
);

LUT6 #(
   .INIT(64'heae7fd56eae7fd56)  
) LUT6_inst8748 (
   .O(to_level3[972]),
   .I0(level4_in[5832]),
   .I1(level4_in[5833]),
   .I2(level4_in[5834]),
   .I3(level4_in[5835]),
   .I4(level4_in[5836]),
   .I5(level4_in[5837])
);

LUT6 #(
   .INIT(64'h4c7156644c715664)  
) LUT6_inst8749 (
   .O(to_level3[973]),
   .I0(level4_in[5838]),
   .I1(level4_in[5839]),
   .I2(level4_in[5840]),
   .I3(level4_in[5841]),
   .I4(level4_in[5842]),
   .I5(level4_in[5843])
);

LUT6 #(
   .INIT(64'h9a0ffec99a0ffec9)  
) LUT6_inst8750 (
   .O(to_level3[974]),
   .I0(level4_in[5844]),
   .I1(level4_in[5845]),
   .I2(level4_in[5846]),
   .I3(level4_in[5847]),
   .I4(level4_in[5848]),
   .I5(level4_in[5849])
);

LUT6 #(
   .INIT(64'h4203098a4203098a)  
) LUT6_inst8751 (
   .O(to_level3[975]),
   .I0(level4_in[5850]),
   .I1(level4_in[5851]),
   .I2(level4_in[5852]),
   .I3(level4_in[5853]),
   .I4(level4_in[5854]),
   .I5(level4_in[5855])
);

LUT6 #(
   .INIT(64'h6bec66376bec6637)  
) LUT6_inst8752 (
   .O(to_level3[976]),
   .I0(level4_in[5856]),
   .I1(level4_in[5857]),
   .I2(level4_in[5858]),
   .I3(level4_in[5859]),
   .I4(level4_in[5860]),
   .I5(level4_in[5861])
);

LUT6 #(
   .INIT(64'ha092ca03a092ca03)  
) LUT6_inst8753 (
   .O(to_level3[977]),
   .I0(level4_in[5862]),
   .I1(level4_in[5863]),
   .I2(level4_in[5864]),
   .I3(level4_in[5865]),
   .I4(level4_in[5866]),
   .I5(level4_in[5867])
);

LUT6 #(
   .INIT(64'h676e2157676e2157)  
) LUT6_inst8754 (
   .O(to_level3[978]),
   .I0(level4_in[5868]),
   .I1(level4_in[5869]),
   .I2(level4_in[5870]),
   .I3(level4_in[5871]),
   .I4(level4_in[5872]),
   .I5(level4_in[5873])
);

LUT6 #(
   .INIT(64'h2cbe4d7b2cbe4d7b)  
) LUT6_inst8755 (
   .O(to_level3[979]),
   .I0(level4_in[5874]),
   .I1(level4_in[5875]),
   .I2(level4_in[5876]),
   .I3(level4_in[5877]),
   .I4(level4_in[5878]),
   .I5(level4_in[5879])
);

LUT6 #(
   .INIT(64'hb6c1b8fdb6c1b8fd)  
) LUT6_inst8756 (
   .O(to_level3[980]),
   .I0(level4_in[5880]),
   .I1(level4_in[5881]),
   .I2(level4_in[5882]),
   .I3(level4_in[5883]),
   .I4(level4_in[5884]),
   .I5(level4_in[5885])
);

LUT6 #(
   .INIT(64'hc8db2b1ec8db2b1e)  
) LUT6_inst8757 (
   .O(to_level3[981]),
   .I0(level4_in[5886]),
   .I1(level4_in[5887]),
   .I2(level4_in[5888]),
   .I3(level4_in[5889]),
   .I4(level4_in[5890]),
   .I5(level4_in[5891])
);

LUT6 #(
   .INIT(64'h8a37b5108a37b510)  
) LUT6_inst8758 (
   .O(to_level3[982]),
   .I0(level4_in[5892]),
   .I1(level4_in[5893]),
   .I2(level4_in[5894]),
   .I3(level4_in[5895]),
   .I4(level4_in[5896]),
   .I5(level4_in[5897])
);

LUT6 #(
   .INIT(64'h8ce3d1018ce3d101)  
) LUT6_inst8759 (
   .O(to_level3[983]),
   .I0(level4_in[5898]),
   .I1(level4_in[5899]),
   .I2(level4_in[5900]),
   .I3(level4_in[5901]),
   .I4(level4_in[5902]),
   .I5(level4_in[5903])
);

LUT6 #(
   .INIT(64'h6862a2246862a224)  
) LUT6_inst8760 (
   .O(to_level3[984]),
   .I0(level4_in[5904]),
   .I1(level4_in[5905]),
   .I2(level4_in[5906]),
   .I3(level4_in[5907]),
   .I4(level4_in[5908]),
   .I5(level4_in[5909])
);

LUT6 #(
   .INIT(64'hd2f9033cd2f9033c)  
) LUT6_inst8761 (
   .O(to_level3[985]),
   .I0(level4_in[5910]),
   .I1(level4_in[5911]),
   .I2(level4_in[5912]),
   .I3(level4_in[5913]),
   .I4(level4_in[5914]),
   .I5(level4_in[5915])
);

LUT6 #(
   .INIT(64'h037d4008037d4008)  
) LUT6_inst8762 (
   .O(to_level3[986]),
   .I0(level4_in[5916]),
   .I1(level4_in[5917]),
   .I2(level4_in[5918]),
   .I3(level4_in[5919]),
   .I4(level4_in[5920]),
   .I5(level4_in[5921])
);

LUT6 #(
   .INIT(64'h8cfe8dc58cfe8dc5)  
) LUT6_inst8763 (
   .O(to_level3[987]),
   .I0(level4_in[5922]),
   .I1(level4_in[5923]),
   .I2(level4_in[5924]),
   .I3(level4_in[5925]),
   .I4(level4_in[5926]),
   .I5(level4_in[5927])
);

LUT6 #(
   .INIT(64'hf618a33bf618a33b)  
) LUT6_inst8764 (
   .O(to_level3[988]),
   .I0(level4_in[5928]),
   .I1(level4_in[5929]),
   .I2(level4_in[5930]),
   .I3(level4_in[5931]),
   .I4(level4_in[5932]),
   .I5(level4_in[5933])
);

LUT6 #(
   .INIT(64'h1429a9f81429a9f8)  
) LUT6_inst8765 (
   .O(to_level3[989]),
   .I0(level4_in[5934]),
   .I1(level4_in[5935]),
   .I2(level4_in[5936]),
   .I3(level4_in[5937]),
   .I4(level4_in[5938]),
   .I5(level4_in[5939])
);

LUT6 #(
   .INIT(64'h1c902afa1c902afa)  
) LUT6_inst8766 (
   .O(to_level3[990]),
   .I0(level4_in[5940]),
   .I1(level4_in[5941]),
   .I2(level4_in[5942]),
   .I3(level4_in[5943]),
   .I4(level4_in[5944]),
   .I5(level4_in[5945])
);

LUT6 #(
   .INIT(64'haef8fb43aef8fb43)  
) LUT6_inst8767 (
   .O(to_level3[991]),
   .I0(level4_in[5946]),
   .I1(level4_in[5947]),
   .I2(level4_in[5948]),
   .I3(level4_in[5949]),
   .I4(level4_in[5950]),
   .I5(level4_in[5951])
);

LUT6 #(
   .INIT(64'h4e5aca774e5aca77)  
) LUT6_inst8768 (
   .O(to_level3[992]),
   .I0(level4_in[5952]),
   .I1(level4_in[5953]),
   .I2(level4_in[5954]),
   .I3(level4_in[5955]),
   .I4(level4_in[5956]),
   .I5(level4_in[5957])
);

LUT6 #(
   .INIT(64'h1c11e9b01c11e9b0)  
) LUT6_inst8769 (
   .O(to_level3[993]),
   .I0(level4_in[5958]),
   .I1(level4_in[5959]),
   .I2(level4_in[5960]),
   .I3(level4_in[5961]),
   .I4(level4_in[5962]),
   .I5(level4_in[5963])
);

LUT6 #(
   .INIT(64'h176d3ab4176d3ab4)  
) LUT6_inst8770 (
   .O(to_level3[994]),
   .I0(level4_in[5964]),
   .I1(level4_in[5965]),
   .I2(level4_in[5966]),
   .I3(level4_in[5967]),
   .I4(level4_in[5968]),
   .I5(level4_in[5969])
);

LUT6 #(
   .INIT(64'h5d0665cd5d0665cd)  
) LUT6_inst8771 (
   .O(to_level3[995]),
   .I0(level4_in[5970]),
   .I1(level4_in[5971]),
   .I2(level4_in[5972]),
   .I3(level4_in[5973]),
   .I4(level4_in[5974]),
   .I5(level4_in[5975])
);

LUT6 #(
   .INIT(64'h462bd810462bd810)  
) LUT6_inst8772 (
   .O(to_level3[996]),
   .I0(level4_in[5976]),
   .I1(level4_in[5977]),
   .I2(level4_in[5978]),
   .I3(level4_in[5979]),
   .I4(level4_in[5980]),
   .I5(level4_in[5981])
);

LUT6 #(
   .INIT(64'h50b64bd950b64bd9)  
) LUT6_inst8773 (
   .O(to_level3[997]),
   .I0(level4_in[5982]),
   .I1(level4_in[5983]),
   .I2(level4_in[5984]),
   .I3(level4_in[5985]),
   .I4(level4_in[5986]),
   .I5(level4_in[5987])
);

LUT6 #(
   .INIT(64'h902d09fa902d09fa)  
) LUT6_inst8774 (
   .O(to_level3[998]),
   .I0(level4_in[5988]),
   .I1(level4_in[5989]),
   .I2(level4_in[5990]),
   .I3(level4_in[5991]),
   .I4(level4_in[5992]),
   .I5(level4_in[5993])
);

LUT6 #(
   .INIT(64'h4afb86ba4afb86ba)  
) LUT6_inst8775 (
   .O(to_level3[999]),
   .I0(level4_in[5994]),
   .I1(level4_in[5995]),
   .I2(level4_in[5996]),
   .I3(level4_in[5997]),
   .I4(level4_in[5998]),
   .I5(level4_in[5999])
);

LUT6 #(
   .INIT(64'h1e1a3d431e1a3d43)  
) LUT6_inst8776 (
   .O(to_level3[1000]),
   .I0(level4_in[6000]),
   .I1(level4_in[6001]),
   .I2(level4_in[6002]),
   .I3(level4_in[6003]),
   .I4(level4_in[6004]),
   .I5(level4_in[6005])
);

LUT6 #(
   .INIT(64'ha0771b8ba0771b8b)  
) LUT6_inst8777 (
   .O(to_level3[1001]),
   .I0(level4_in[6006]),
   .I1(level4_in[6007]),
   .I2(level4_in[6008]),
   .I3(level4_in[6009]),
   .I4(level4_in[6010]),
   .I5(level4_in[6011])
);

LUT6 #(
   .INIT(64'h3864df533864df53)  
) LUT6_inst8778 (
   .O(to_level3[1002]),
   .I0(level4_in[6012]),
   .I1(level4_in[6013]),
   .I2(level4_in[6014]),
   .I3(level4_in[6015]),
   .I4(level4_in[6016]),
   .I5(level4_in[6017])
);

LUT6 #(
   .INIT(64'h52e6083352e60833)  
) LUT6_inst8779 (
   .O(to_level3[1003]),
   .I0(level4_in[6018]),
   .I1(level4_in[6019]),
   .I2(level4_in[6020]),
   .I3(level4_in[6021]),
   .I4(level4_in[6022]),
   .I5(level4_in[6023])
);

LUT6 #(
   .INIT(64'hedf2ea13edf2ea13)  
) LUT6_inst8780 (
   .O(to_level3[1004]),
   .I0(level4_in[6024]),
   .I1(level4_in[6025]),
   .I2(level4_in[6026]),
   .I3(level4_in[6027]),
   .I4(level4_in[6028]),
   .I5(level4_in[6029])
);

LUT6 #(
   .INIT(64'he3110503e3110503)  
) LUT6_inst8781 (
   .O(to_level3[1005]),
   .I0(level4_in[6030]),
   .I1(level4_in[6031]),
   .I2(level4_in[6032]),
   .I3(level4_in[6033]),
   .I4(level4_in[6034]),
   .I5(level4_in[6035])
);

LUT6 #(
   .INIT(64'hcd45964acd45964a)  
) LUT6_inst8782 (
   .O(to_level3[1006]),
   .I0(level4_in[6036]),
   .I1(level4_in[6037]),
   .I2(level4_in[6038]),
   .I3(level4_in[6039]),
   .I4(level4_in[6040]),
   .I5(level4_in[6041])
);

LUT6 #(
   .INIT(64'h9841076998410769)  
) LUT6_inst8783 (
   .O(to_level3[1007]),
   .I0(level4_in[6042]),
   .I1(level4_in[6043]),
   .I2(level4_in[6044]),
   .I3(level4_in[6045]),
   .I4(level4_in[6046]),
   .I5(level4_in[6047])
);

LUT6 #(
   .INIT(64'h33ebb17533ebb175)  
) LUT6_inst8784 (
   .O(to_level3[1008]),
   .I0(level4_in[6048]),
   .I1(level4_in[6049]),
   .I2(level4_in[6050]),
   .I3(level4_in[6051]),
   .I4(level4_in[6052]),
   .I5(level4_in[6053])
);

LUT6 #(
   .INIT(64'h4aedb3524aedb352)  
) LUT6_inst8785 (
   .O(to_level3[1009]),
   .I0(level4_in[6054]),
   .I1(level4_in[6055]),
   .I2(level4_in[6056]),
   .I3(level4_in[6057]),
   .I4(level4_in[6058]),
   .I5(level4_in[6059])
);

LUT6 #(
   .INIT(64'h523fc931523fc931)  
) LUT6_inst8786 (
   .O(to_level3[1010]),
   .I0(level4_in[6060]),
   .I1(level4_in[6061]),
   .I2(level4_in[6062]),
   .I3(level4_in[6063]),
   .I4(level4_in[6064]),
   .I5(level4_in[6065])
);

LUT6 #(
   .INIT(64'h09146e3e09146e3e)  
) LUT6_inst8787 (
   .O(to_level3[1011]),
   .I0(level4_in[6066]),
   .I1(level4_in[6067]),
   .I2(level4_in[6068]),
   .I3(level4_in[6069]),
   .I4(level4_in[6070]),
   .I5(level4_in[6071])
);

LUT6 #(
   .INIT(64'h89bbf43589bbf435)  
) LUT6_inst8788 (
   .O(to_level3[1012]),
   .I0(level4_in[6072]),
   .I1(level4_in[6073]),
   .I2(level4_in[6074]),
   .I3(level4_in[6075]),
   .I4(level4_in[6076]),
   .I5(level4_in[6077])
);

LUT6 #(
   .INIT(64'hed72426eed72426e)  
) LUT6_inst8789 (
   .O(to_level3[1013]),
   .I0(level4_in[6078]),
   .I1(level4_in[6079]),
   .I2(level4_in[6080]),
   .I3(level4_in[6081]),
   .I4(level4_in[6082]),
   .I5(level4_in[6083])
);

LUT6 #(
   .INIT(64'h140c906c140c906c)  
) LUT6_inst8790 (
   .O(to_level3[1014]),
   .I0(level4_in[6084]),
   .I1(level4_in[6085]),
   .I2(level4_in[6086]),
   .I3(level4_in[6087]),
   .I4(level4_in[6088]),
   .I5(level4_in[6089])
);

LUT6 #(
   .INIT(64'h29a29bab29a29bab)  
) LUT6_inst8791 (
   .O(to_level3[1015]),
   .I0(level4_in[6090]),
   .I1(level4_in[6091]),
   .I2(level4_in[6092]),
   .I3(level4_in[6093]),
   .I4(level4_in[6094]),
   .I5(level4_in[6095])
);

LUT6 #(
   .INIT(64'ha052b521a052b521)  
) LUT6_inst8792 (
   .O(to_level3[1016]),
   .I0(level4_in[6096]),
   .I1(level4_in[6097]),
   .I2(level4_in[6098]),
   .I3(level4_in[6099]),
   .I4(level4_in[6100]),
   .I5(level4_in[6101])
);

LUT6 #(
   .INIT(64'h4de28f124de28f12)  
) LUT6_inst8793 (
   .O(to_level3[1017]),
   .I0(level4_in[6102]),
   .I1(level4_in[6103]),
   .I2(level4_in[6104]),
   .I3(level4_in[6105]),
   .I4(level4_in[6106]),
   .I5(level4_in[6107])
);

LUT6 #(
   .INIT(64'h3804e7353804e735)  
) LUT6_inst8794 (
   .O(to_level3[1018]),
   .I0(level4_in[6108]),
   .I1(level4_in[6109]),
   .I2(level4_in[6110]),
   .I3(level4_in[6111]),
   .I4(level4_in[6112]),
   .I5(level4_in[6113])
);

LUT6 #(
   .INIT(64'h46aeba8c46aeba8c)  
) LUT6_inst8795 (
   .O(to_level3[1019]),
   .I0(level4_in[6114]),
   .I1(level4_in[6115]),
   .I2(level4_in[6116]),
   .I3(level4_in[6117]),
   .I4(level4_in[6118]),
   .I5(level4_in[6119])
);

LUT6 #(
   .INIT(64'h604ea8fd604ea8fd)  
) LUT6_inst8796 (
   .O(to_level3[1020]),
   .I0(level4_in[6120]),
   .I1(level4_in[6121]),
   .I2(level4_in[6122]),
   .I3(level4_in[6123]),
   .I4(level4_in[6124]),
   .I5(level4_in[6125])
);

LUT6 #(
   .INIT(64'hd48bf73cd48bf73c)  
) LUT6_inst8797 (
   .O(to_level3[1021]),
   .I0(level4_in[6126]),
   .I1(level4_in[6127]),
   .I2(level4_in[6128]),
   .I3(level4_in[6129]),
   .I4(level4_in[6130]),
   .I5(level4_in[6131])
);

LUT6 #(
   .INIT(64'h4dea3a9a4dea3a9a)  
) LUT6_inst8798 (
   .O(to_level3[1022]),
   .I0(level4_in[6132]),
   .I1(level4_in[6133]),
   .I2(level4_in[6134]),
   .I3(level4_in[6135]),
   .I4(level4_in[6136]),
   .I5(level4_in[6137])
);

LUT6 #(
   .INIT(64'h2752998327529983)  
) LUT6_inst8799 (
   .O(to_level3[1023]),
   .I0(level4_in[6138]),
   .I1(level4_in[6139]),
   .I2(level4_in[6140]),
   .I3(level4_in[6141]),
   .I4(level4_in[6142]),
   .I5(level4_in[6143])
);

LUT6 #(
   .INIT(64'hdd792022dd792022)  
) LUT6_inst8800 (
   .O(to_level3[1024]),
   .I0(level4_in[6144]),
   .I1(level4_in[6145]),
   .I2(level4_in[6146]),
   .I3(level4_in[6147]),
   .I4(level4_in[6148]),
   .I5(level4_in[6149])
);

LUT6 #(
   .INIT(64'h5549a7605549a760)  
) LUT6_inst8801 (
   .O(to_level3[1025]),
   .I0(level4_in[6150]),
   .I1(level4_in[6151]),
   .I2(level4_in[6152]),
   .I3(level4_in[6153]),
   .I4(level4_in[6154]),
   .I5(level4_in[6155])
);

LUT6 #(
   .INIT(64'hd8afb3bdd8afb3bd)  
) LUT6_inst8802 (
   .O(to_level3[1026]),
   .I0(level4_in[6156]),
   .I1(level4_in[6157]),
   .I2(level4_in[6158]),
   .I3(level4_in[6159]),
   .I4(level4_in[6160]),
   .I5(level4_in[6161])
);

LUT6 #(
   .INIT(64'h882ac645882ac645)  
) LUT6_inst8803 (
   .O(to_level3[1027]),
   .I0(level4_in[6162]),
   .I1(level4_in[6163]),
   .I2(level4_in[6164]),
   .I3(level4_in[6165]),
   .I4(level4_in[6166]),
   .I5(level4_in[6167])
);

LUT6 #(
   .INIT(64'h211a125c211a125c)  
) LUT6_inst8804 (
   .O(to_level3[1028]),
   .I0(level4_in[6168]),
   .I1(level4_in[6169]),
   .I2(level4_in[6170]),
   .I3(level4_in[6171]),
   .I4(level4_in[6172]),
   .I5(level4_in[6173])
);

LUT6 #(
   .INIT(64'hb9637f45b9637f45)  
) LUT6_inst8805 (
   .O(to_level3[1029]),
   .I0(level4_in[6174]),
   .I1(level4_in[6175]),
   .I2(level4_in[6176]),
   .I3(level4_in[6177]),
   .I4(level4_in[6178]),
   .I5(level4_in[6179])
);

LUT6 #(
   .INIT(64'hb8c03065b8c03065)  
) LUT6_inst8806 (
   .O(to_level3[1030]),
   .I0(level4_in[6180]),
   .I1(level4_in[6181]),
   .I2(level4_in[6182]),
   .I3(level4_in[6183]),
   .I4(level4_in[6184]),
   .I5(level4_in[6185])
);

LUT6 #(
   .INIT(64'h422b4e5c422b4e5c)  
) LUT6_inst8807 (
   .O(to_level3[1031]),
   .I0(level4_in[6186]),
   .I1(level4_in[6187]),
   .I2(level4_in[6188]),
   .I3(level4_in[6189]),
   .I4(level4_in[6190]),
   .I5(level4_in[6191])
);

LUT6 #(
   .INIT(64'hbee531ccbee531cc)  
) LUT6_inst8808 (
   .O(to_level3[1032]),
   .I0(level4_in[6192]),
   .I1(level4_in[6193]),
   .I2(level4_in[6194]),
   .I3(level4_in[6195]),
   .I4(level4_in[6196]),
   .I5(level4_in[6197])
);

LUT6 #(
   .INIT(64'hd38ecb59d38ecb59)  
) LUT6_inst8809 (
   .O(to_level3[1033]),
   .I0(level4_in[6198]),
   .I1(level4_in[6199]),
   .I2(level4_in[6200]),
   .I3(level4_in[6201]),
   .I4(level4_in[6202]),
   .I5(level4_in[6203])
);

LUT6 #(
   .INIT(64'hd5273daed5273dae)  
) LUT6_inst8810 (
   .O(to_level3[1034]),
   .I0(level4_in[6204]),
   .I1(level4_in[6205]),
   .I2(level4_in[6206]),
   .I3(level4_in[6207]),
   .I4(level4_in[6208]),
   .I5(level4_in[6209])
);

LUT6 #(
   .INIT(64'h8498e2278498e227)  
) LUT6_inst8811 (
   .O(to_level3[1035]),
   .I0(level4_in[6210]),
   .I1(level4_in[6211]),
   .I2(level4_in[6212]),
   .I3(level4_in[6213]),
   .I4(level4_in[6214]),
   .I5(level4_in[6215])
);

LUT6 #(
   .INIT(64'h11e8d3d911e8d3d9)  
) LUT6_inst8812 (
   .O(to_level3[1036]),
   .I0(level4_in[6216]),
   .I1(level4_in[6217]),
   .I2(level4_in[6218]),
   .I3(level4_in[6219]),
   .I4(level4_in[6220]),
   .I5(level4_in[6221])
);

LUT6 #(
   .INIT(64'h00bbbdfb00bbbdfb)  
) LUT6_inst8813 (
   .O(to_level3[1037]),
   .I0(level4_in[6222]),
   .I1(level4_in[6223]),
   .I2(level4_in[6224]),
   .I3(level4_in[6225]),
   .I4(level4_in[6226]),
   .I5(level4_in[6227])
);

LUT6 #(
   .INIT(64'h3d29e8083d29e808)  
) LUT6_inst8814 (
   .O(to_level3[1038]),
   .I0(level4_in[6228]),
   .I1(level4_in[6229]),
   .I2(level4_in[6230]),
   .I3(level4_in[6231]),
   .I4(level4_in[6232]),
   .I5(level4_in[6233])
);

LUT6 #(
   .INIT(64'h955f0019955f0019)  
) LUT6_inst8815 (
   .O(to_level3[1039]),
   .I0(level4_in[6234]),
   .I1(level4_in[6235]),
   .I2(level4_in[6236]),
   .I3(level4_in[6237]),
   .I4(level4_in[6238]),
   .I5(level4_in[6239])
);

LUT6 #(
   .INIT(64'hddb0edbcddb0edbc)  
) LUT6_inst8816 (
   .O(to_level3[1040]),
   .I0(level4_in[6240]),
   .I1(level4_in[6241]),
   .I2(level4_in[6242]),
   .I3(level4_in[6243]),
   .I4(level4_in[6244]),
   .I5(level4_in[6245])
);

LUT6 #(
   .INIT(64'h7477137274771372)  
) LUT6_inst8817 (
   .O(to_level3[1041]),
   .I0(level4_in[6246]),
   .I1(level4_in[6247]),
   .I2(level4_in[6248]),
   .I3(level4_in[6249]),
   .I4(level4_in[6250]),
   .I5(level4_in[6251])
);

LUT6 #(
   .INIT(64'h3b68ff573b68ff57)  
) LUT6_inst8818 (
   .O(to_level3[1042]),
   .I0(level4_in[6252]),
   .I1(level4_in[6253]),
   .I2(level4_in[6254]),
   .I3(level4_in[6255]),
   .I4(level4_in[6256]),
   .I5(level4_in[6257])
);

LUT6 #(
   .INIT(64'hd58dd96ad58dd96a)  
) LUT6_inst8819 (
   .O(to_level3[1043]),
   .I0(level4_in[6258]),
   .I1(level4_in[6259]),
   .I2(level4_in[6260]),
   .I3(level4_in[6261]),
   .I4(level4_in[6262]),
   .I5(level4_in[6263])
);

LUT6 #(
   .INIT(64'hdf260674df260674)  
) LUT6_inst8820 (
   .O(to_level3[1044]),
   .I0(level4_in[6264]),
   .I1(level4_in[6265]),
   .I2(level4_in[6266]),
   .I3(level4_in[6267]),
   .I4(level4_in[6268]),
   .I5(level4_in[6269])
);

LUT6 #(
   .INIT(64'hcbac3d06cbac3d06)  
) LUT6_inst8821 (
   .O(to_level3[1045]),
   .I0(level4_in[6270]),
   .I1(level4_in[6271]),
   .I2(level4_in[6272]),
   .I3(level4_in[6273]),
   .I4(level4_in[6274]),
   .I5(level4_in[6275])
);

LUT6 #(
   .INIT(64'h2d04ef042d04ef04)  
) LUT6_inst8822 (
   .O(to_level3[1046]),
   .I0(level4_in[6276]),
   .I1(level4_in[6277]),
   .I2(level4_in[6278]),
   .I3(level4_in[6279]),
   .I4(level4_in[6280]),
   .I5(level4_in[6281])
);

LUT6 #(
   .INIT(64'hcfc90c35cfc90c35)  
) LUT6_inst8823 (
   .O(to_level3[1047]),
   .I0(level4_in[6282]),
   .I1(level4_in[6283]),
   .I2(level4_in[6284]),
   .I3(level4_in[6285]),
   .I4(level4_in[6286]),
   .I5(level4_in[6287])
);

LUT6 #(
   .INIT(64'h0c8f74350c8f7435)  
) LUT6_inst8824 (
   .O(to_level3[1048]),
   .I0(level4_in[6288]),
   .I1(level4_in[6289]),
   .I2(level4_in[6290]),
   .I3(level4_in[6291]),
   .I4(level4_in[6292]),
   .I5(level4_in[6293])
);

LUT6 #(
   .INIT(64'h8b9f3dd78b9f3dd7)  
) LUT6_inst8825 (
   .O(to_level3[1049]),
   .I0(level4_in[6294]),
   .I1(level4_in[6295]),
   .I2(level4_in[6296]),
   .I3(level4_in[6297]),
   .I4(level4_in[6298]),
   .I5(level4_in[6299])
);

LUT6 #(
   .INIT(64'h9e89d8ad9e89d8ad)  
) LUT6_inst8826 (
   .O(to_level3[1050]),
   .I0(level4_in[6300]),
   .I1(level4_in[6301]),
   .I2(level4_in[6302]),
   .I3(level4_in[6303]),
   .I4(level4_in[6304]),
   .I5(level4_in[6305])
);

LUT6 #(
   .INIT(64'h33f8fcab33f8fcab)  
) LUT6_inst8827 (
   .O(to_level3[1051]),
   .I0(level4_in[6306]),
   .I1(level4_in[6307]),
   .I2(level4_in[6308]),
   .I3(level4_in[6309]),
   .I4(level4_in[6310]),
   .I5(level4_in[6311])
);

LUT6 #(
   .INIT(64'h918c4ec6918c4ec6)  
) LUT6_inst8828 (
   .O(to_level3[1052]),
   .I0(level4_in[6312]),
   .I1(level4_in[6313]),
   .I2(level4_in[6314]),
   .I3(level4_in[6315]),
   .I4(level4_in[6316]),
   .I5(level4_in[6317])
);

LUT6 #(
   .INIT(64'h80e5c4d780e5c4d7)  
) LUT6_inst8829 (
   .O(to_level3[1053]),
   .I0(level4_in[6318]),
   .I1(level4_in[6319]),
   .I2(level4_in[6320]),
   .I3(level4_in[6321]),
   .I4(level4_in[6322]),
   .I5(level4_in[6323])
);

LUT6 #(
   .INIT(64'h40dd889440dd8894)  
) LUT6_inst8830 (
   .O(to_level3[1054]),
   .I0(level4_in[6324]),
   .I1(level4_in[6325]),
   .I2(level4_in[6326]),
   .I3(level4_in[6327]),
   .I4(level4_in[6328]),
   .I5(level4_in[6329])
);

LUT6 #(
   .INIT(64'hfbabb9b2fbabb9b2)  
) LUT6_inst8831 (
   .O(to_level3[1055]),
   .I0(level4_in[6330]),
   .I1(level4_in[6331]),
   .I2(level4_in[6332]),
   .I3(level4_in[6333]),
   .I4(level4_in[6334]),
   .I5(level4_in[6335])
);

LUT6 #(
   .INIT(64'hc46bec03c46bec03)  
) LUT6_inst8832 (
   .O(to_level3[1056]),
   .I0(level4_in[6336]),
   .I1(level4_in[6337]),
   .I2(level4_in[6338]),
   .I3(level4_in[6339]),
   .I4(level4_in[6340]),
   .I5(level4_in[6341])
);

LUT6 #(
   .INIT(64'hc2cc620ec2cc620e)  
) LUT6_inst8833 (
   .O(to_level3[1057]),
   .I0(level4_in[6342]),
   .I1(level4_in[6343]),
   .I2(level4_in[6344]),
   .I3(level4_in[6345]),
   .I4(level4_in[6346]),
   .I5(level4_in[6347])
);

LUT6 #(
   .INIT(64'h1c46510e1c46510e)  
) LUT6_inst8834 (
   .O(to_level3[1058]),
   .I0(level4_in[6348]),
   .I1(level4_in[6349]),
   .I2(level4_in[6350]),
   .I3(level4_in[6351]),
   .I4(level4_in[6352]),
   .I5(level4_in[6353])
);

LUT6 #(
   .INIT(64'h197f0523197f0523)  
) LUT6_inst8835 (
   .O(to_level3[1059]),
   .I0(level4_in[6354]),
   .I1(level4_in[6355]),
   .I2(level4_in[6356]),
   .I3(level4_in[6357]),
   .I4(level4_in[6358]),
   .I5(level4_in[6359])
);

LUT6 #(
   .INIT(64'h1498a6ad1498a6ad)  
) LUT6_inst8836 (
   .O(to_level3[1060]),
   .I0(level4_in[6360]),
   .I1(level4_in[6361]),
   .I2(level4_in[6362]),
   .I3(level4_in[6363]),
   .I4(level4_in[6364]),
   .I5(level4_in[6365])
);

LUT6 #(
   .INIT(64'h5f9ffb285f9ffb28)  
) LUT6_inst8837 (
   .O(to_level3[1061]),
   .I0(level4_in[6366]),
   .I1(level4_in[6367]),
   .I2(level4_in[6368]),
   .I3(level4_in[6369]),
   .I4(level4_in[6370]),
   .I5(level4_in[6371])
);

LUT6 #(
   .INIT(64'hf5947148f5947148)  
) LUT6_inst8838 (
   .O(to_level3[1062]),
   .I0(level4_in[6372]),
   .I1(level4_in[6373]),
   .I2(level4_in[6374]),
   .I3(level4_in[6375]),
   .I4(level4_in[6376]),
   .I5(level4_in[6377])
);

LUT6 #(
   .INIT(64'hd9cf43ecd9cf43ec)  
) LUT6_inst8839 (
   .O(to_level3[1063]),
   .I0(level4_in[6378]),
   .I1(level4_in[6379]),
   .I2(level4_in[6380]),
   .I3(level4_in[6381]),
   .I4(level4_in[6382]),
   .I5(level4_in[6383])
);

LUT6 #(
   .INIT(64'h19fa746919fa7469)  
) LUT6_inst8840 (
   .O(to_level3[1064]),
   .I0(level4_in[6384]),
   .I1(level4_in[6385]),
   .I2(level4_in[6386]),
   .I3(level4_in[6387]),
   .I4(level4_in[6388]),
   .I5(level4_in[6389])
);

LUT6 #(
   .INIT(64'h7d6832147d683214)  
) LUT6_inst8841 (
   .O(to_level3[1065]),
   .I0(level4_in[6390]),
   .I1(level4_in[6391]),
   .I2(level4_in[6392]),
   .I3(level4_in[6393]),
   .I4(level4_in[6394]),
   .I5(level4_in[6395])
);

LUT6 #(
   .INIT(64'h37e58b4137e58b41)  
) LUT6_inst8842 (
   .O(to_level3[1066]),
   .I0(level4_in[6396]),
   .I1(level4_in[6397]),
   .I2(level4_in[6398]),
   .I3(level4_in[6399]),
   .I4(level4_in[6400]),
   .I5(level4_in[6401])
);

LUT6 #(
   .INIT(64'h7d1165807d116580)  
) LUT6_inst8843 (
   .O(to_level3[1067]),
   .I0(level4_in[6402]),
   .I1(level4_in[6403]),
   .I2(level4_in[6404]),
   .I3(level4_in[6405]),
   .I4(level4_in[6406]),
   .I5(level4_in[6407])
);

LUT6 #(
   .INIT(64'h90f4d0b290f4d0b2)  
) LUT6_inst8844 (
   .O(to_level3[1068]),
   .I0(level4_in[6408]),
   .I1(level4_in[6409]),
   .I2(level4_in[6410]),
   .I3(level4_in[6411]),
   .I4(level4_in[6412]),
   .I5(level4_in[6413])
);

LUT6 #(
   .INIT(64'h9e6b88589e6b8858)  
) LUT6_inst8845 (
   .O(to_level3[1069]),
   .I0(level4_in[6414]),
   .I1(level4_in[6415]),
   .I2(level4_in[6416]),
   .I3(level4_in[6417]),
   .I4(level4_in[6418]),
   .I5(level4_in[6419])
);

LUT6 #(
   .INIT(64'h15b3fe3c15b3fe3c)  
) LUT6_inst8846 (
   .O(to_level3[1070]),
   .I0(level4_in[6420]),
   .I1(level4_in[6421]),
   .I2(level4_in[6422]),
   .I3(level4_in[6423]),
   .I4(level4_in[6424]),
   .I5(level4_in[6425])
);

LUT6 #(
   .INIT(64'h726910c5726910c5)  
) LUT6_inst8847 (
   .O(to_level3[1071]),
   .I0(level4_in[6426]),
   .I1(level4_in[6427]),
   .I2(level4_in[6428]),
   .I3(level4_in[6429]),
   .I4(level4_in[6430]),
   .I5(level4_in[6431])
);

LUT6 #(
   .INIT(64'h6356032563560325)  
) LUT6_inst8848 (
   .O(to_level3[1072]),
   .I0(level4_in[6432]),
   .I1(level4_in[6433]),
   .I2(level4_in[6434]),
   .I3(level4_in[6435]),
   .I4(level4_in[6436]),
   .I5(level4_in[6437])
);

LUT6 #(
   .INIT(64'h586af39d586af39d)  
) LUT6_inst8849 (
   .O(to_level3[1073]),
   .I0(level4_in[6438]),
   .I1(level4_in[6439]),
   .I2(level4_in[6440]),
   .I3(level4_in[6441]),
   .I4(level4_in[6442]),
   .I5(level4_in[6443])
);

LUT6 #(
   .INIT(64'h1c04ded31c04ded3)  
) LUT6_inst8850 (
   .O(to_level3[1074]),
   .I0(level4_in[6444]),
   .I1(level4_in[6445]),
   .I2(level4_in[6446]),
   .I3(level4_in[6447]),
   .I4(level4_in[6448]),
   .I5(level4_in[6449])
);

LUT6 #(
   .INIT(64'h9c45c7089c45c708)  
) LUT6_inst8851 (
   .O(to_level3[1075]),
   .I0(level4_in[6450]),
   .I1(level4_in[6451]),
   .I2(level4_in[6452]),
   .I3(level4_in[6453]),
   .I4(level4_in[6454]),
   .I5(level4_in[6455])
);

LUT6 #(
   .INIT(64'ha22de7f5a22de7f5)  
) LUT6_inst8852 (
   .O(to_level3[1076]),
   .I0(level4_in[6456]),
   .I1(level4_in[6457]),
   .I2(level4_in[6458]),
   .I3(level4_in[6459]),
   .I4(level4_in[6460]),
   .I5(level4_in[6461])
);

LUT6 #(
   .INIT(64'h7c7106317c710631)  
) LUT6_inst8853 (
   .O(to_level3[1077]),
   .I0(level4_in[6462]),
   .I1(level4_in[6463]),
   .I2(level4_in[6464]),
   .I3(level4_in[6465]),
   .I4(level4_in[6466]),
   .I5(level4_in[6467])
);

LUT6 #(
   .INIT(64'he13bcc11e13bcc11)  
) LUT6_inst8854 (
   .O(to_level3[1078]),
   .I0(level4_in[6468]),
   .I1(level4_in[6469]),
   .I2(level4_in[6470]),
   .I3(level4_in[6471]),
   .I4(level4_in[6472]),
   .I5(level4_in[6473])
);

LUT6 #(
   .INIT(64'h88615ec988615ec9)  
) LUT6_inst8855 (
   .O(to_level3[1079]),
   .I0(level4_in[6474]),
   .I1(level4_in[6475]),
   .I2(level4_in[6476]),
   .I3(level4_in[6477]),
   .I4(level4_in[6478]),
   .I5(level4_in[6479])
);

LUT6 #(
   .INIT(64'ha613076aa613076a)  
) LUT6_inst8856 (
   .O(to_level3[1080]),
   .I0(level4_in[6480]),
   .I1(level4_in[6481]),
   .I2(level4_in[6482]),
   .I3(level4_in[6483]),
   .I4(level4_in[6484]),
   .I5(level4_in[6485])
);

LUT6 #(
   .INIT(64'hc43c3696c43c3696)  
) LUT6_inst8857 (
   .O(to_level3[1081]),
   .I0(level4_in[6486]),
   .I1(level4_in[6487]),
   .I2(level4_in[6488]),
   .I3(level4_in[6489]),
   .I4(level4_in[6490]),
   .I5(level4_in[6491])
);

LUT6 #(
   .INIT(64'h40073c9940073c99)  
) LUT6_inst8858 (
   .O(to_level3[1082]),
   .I0(level4_in[6492]),
   .I1(level4_in[6493]),
   .I2(level4_in[6494]),
   .I3(level4_in[6495]),
   .I4(level4_in[6496]),
   .I5(level4_in[6497])
);

LUT6 #(
   .INIT(64'h6c177b5c6c177b5c)  
) LUT6_inst8859 (
   .O(to_level3[1083]),
   .I0(level4_in[6498]),
   .I1(level4_in[6499]),
   .I2(level4_in[6500]),
   .I3(level4_in[6501]),
   .I4(level4_in[6502]),
   .I5(level4_in[6503])
);

LUT6 #(
   .INIT(64'ha1fc7ecea1fc7ece)  
) LUT6_inst8860 (
   .O(to_level3[1084]),
   .I0(level4_in[6504]),
   .I1(level4_in[6505]),
   .I2(level4_in[6506]),
   .I3(level4_in[6507]),
   .I4(level4_in[6508]),
   .I5(level4_in[6509])
);

LUT6 #(
   .INIT(64'h5171690451716904)  
) LUT6_inst8861 (
   .O(to_level3[1085]),
   .I0(level4_in[6510]),
   .I1(level4_in[6511]),
   .I2(level4_in[6512]),
   .I3(level4_in[6513]),
   .I4(level4_in[6514]),
   .I5(level4_in[6515])
);

LUT6 #(
   .INIT(64'h3f9520f13f9520f1)  
) LUT6_inst8862 (
   .O(to_level3[1086]),
   .I0(level4_in[6516]),
   .I1(level4_in[6517]),
   .I2(level4_in[6518]),
   .I3(level4_in[6519]),
   .I4(level4_in[6520]),
   .I5(level4_in[6521])
);

LUT6 #(
   .INIT(64'h35fc83ea35fc83ea)  
) LUT6_inst8863 (
   .O(to_level3[1087]),
   .I0(level4_in[6522]),
   .I1(level4_in[6523]),
   .I2(level4_in[6524]),
   .I3(level4_in[6525]),
   .I4(level4_in[6526]),
   .I5(level4_in[6527])
);

LUT6 #(
   .INIT(64'h4c4b37134c4b3713)  
) LUT6_inst8864 (
   .O(to_level3[1088]),
   .I0(level4_in[6528]),
   .I1(level4_in[6529]),
   .I2(level4_in[6530]),
   .I3(level4_in[6531]),
   .I4(level4_in[6532]),
   .I5(level4_in[6533])
);

LUT6 #(
   .INIT(64'h6ea423a56ea423a5)  
) LUT6_inst8865 (
   .O(to_level3[1089]),
   .I0(level4_in[6534]),
   .I1(level4_in[6535]),
   .I2(level4_in[6536]),
   .I3(level4_in[6537]),
   .I4(level4_in[6538]),
   .I5(level4_in[6539])
);

LUT6 #(
   .INIT(64'hee7c3cd3ee7c3cd3)  
) LUT6_inst8866 (
   .O(to_level3[1090]),
   .I0(level4_in[6540]),
   .I1(level4_in[6541]),
   .I2(level4_in[6542]),
   .I3(level4_in[6543]),
   .I4(level4_in[6544]),
   .I5(level4_in[6545])
);

LUT6 #(
   .INIT(64'h49105c9149105c91)  
) LUT6_inst8867 (
   .O(to_level3[1091]),
   .I0(level4_in[6546]),
   .I1(level4_in[6547]),
   .I2(level4_in[6548]),
   .I3(level4_in[6549]),
   .I4(level4_in[6550]),
   .I5(level4_in[6551])
);

LUT6 #(
   .INIT(64'h3ab0af4c3ab0af4c)  
) LUT6_inst8868 (
   .O(to_level3[1092]),
   .I0(level4_in[6552]),
   .I1(level4_in[6553]),
   .I2(level4_in[6554]),
   .I3(level4_in[6555]),
   .I4(level4_in[6556]),
   .I5(level4_in[6557])
);

LUT6 #(
   .INIT(64'h5d84eb995d84eb99)  
) LUT6_inst8869 (
   .O(to_level3[1093]),
   .I0(level4_in[6558]),
   .I1(level4_in[6559]),
   .I2(level4_in[6560]),
   .I3(level4_in[6561]),
   .I4(level4_in[6562]),
   .I5(level4_in[6563])
);

LUT6 #(
   .INIT(64'h71b3c58e71b3c58e)  
) LUT6_inst8870 (
   .O(to_level3[1094]),
   .I0(level4_in[6564]),
   .I1(level4_in[6565]),
   .I2(level4_in[6566]),
   .I3(level4_in[6567]),
   .I4(level4_in[6568]),
   .I5(level4_in[6569])
);

LUT6 #(
   .INIT(64'h18f2ac7318f2ac73)  
) LUT6_inst8871 (
   .O(to_level3[1095]),
   .I0(level4_in[6570]),
   .I1(level4_in[6571]),
   .I2(level4_in[6572]),
   .I3(level4_in[6573]),
   .I4(level4_in[6574]),
   .I5(level4_in[6575])
);

LUT6 #(
   .INIT(64'h4684024446840244)  
) LUT6_inst8872 (
   .O(to_level3[1096]),
   .I0(level4_in[6576]),
   .I1(level4_in[6577]),
   .I2(level4_in[6578]),
   .I3(level4_in[6579]),
   .I4(level4_in[6580]),
   .I5(level4_in[6581])
);

LUT6 #(
   .INIT(64'h983e88e6983e88e6)  
) LUT6_inst8873 (
   .O(to_level3[1097]),
   .I0(level4_in[6582]),
   .I1(level4_in[6583]),
   .I2(level4_in[6584]),
   .I3(level4_in[6585]),
   .I4(level4_in[6586]),
   .I5(level4_in[6587])
);

LUT6 #(
   .INIT(64'h7aa9d0857aa9d085)  
) LUT6_inst8874 (
   .O(to_level3[1098]),
   .I0(level4_in[6588]),
   .I1(level4_in[6589]),
   .I2(level4_in[6590]),
   .I3(level4_in[6591]),
   .I4(level4_in[6592]),
   .I5(level4_in[6593])
);

LUT6 #(
   .INIT(64'h385dbb87385dbb87)  
) LUT6_inst8875 (
   .O(to_level3[1099]),
   .I0(level4_in[6594]),
   .I1(level4_in[6595]),
   .I2(level4_in[6596]),
   .I3(level4_in[6597]),
   .I4(level4_in[6598]),
   .I5(level4_in[6599])
);

LUT6 #(
   .INIT(64'h844f1de8844f1de8)  
) LUT6_inst8876 (
   .O(to_level3[1100]),
   .I0(level4_in[6600]),
   .I1(level4_in[6601]),
   .I2(level4_in[6602]),
   .I3(level4_in[6603]),
   .I4(level4_in[6604]),
   .I5(level4_in[6605])
);

LUT6 #(
   .INIT(64'he55aa152e55aa152)  
) LUT6_inst8877 (
   .O(to_level3[1101]),
   .I0(level4_in[6606]),
   .I1(level4_in[6607]),
   .I2(level4_in[6608]),
   .I3(level4_in[6609]),
   .I4(level4_in[6610]),
   .I5(level4_in[6611])
);

LUT6 #(
   .INIT(64'h6f2ef2e16f2ef2e1)  
) LUT6_inst8878 (
   .O(to_level3[1102]),
   .I0(level4_in[6612]),
   .I1(level4_in[6613]),
   .I2(level4_in[6614]),
   .I3(level4_in[6615]),
   .I4(level4_in[6616]),
   .I5(level4_in[6617])
);

LUT6 #(
   .INIT(64'h5b9750875b975087)  
) LUT6_inst8879 (
   .O(to_level3[1103]),
   .I0(level4_in[6618]),
   .I1(level4_in[6619]),
   .I2(level4_in[6620]),
   .I3(level4_in[6621]),
   .I4(level4_in[6622]),
   .I5(level4_in[6623])
);

LUT6 #(
   .INIT(64'h1ff74edb1ff74edb)  
) LUT6_inst8880 (
   .O(to_level3[1104]),
   .I0(level4_in[6624]),
   .I1(level4_in[6625]),
   .I2(level4_in[6626]),
   .I3(level4_in[6627]),
   .I4(level4_in[6628]),
   .I5(level4_in[6629])
);

LUT6 #(
   .INIT(64'h0edf7ecd0edf7ecd)  
) LUT6_inst8881 (
   .O(to_level3[1105]),
   .I0(level4_in[6630]),
   .I1(level4_in[6631]),
   .I2(level4_in[6632]),
   .I3(level4_in[6633]),
   .I4(level4_in[6634]),
   .I5(level4_in[6635])
);

LUT6 #(
   .INIT(64'h115b80ff115b80ff)  
) LUT6_inst8882 (
   .O(to_level3[1106]),
   .I0(level4_in[6636]),
   .I1(level4_in[6637]),
   .I2(level4_in[6638]),
   .I3(level4_in[6639]),
   .I4(level4_in[6640]),
   .I5(level4_in[6641])
);

LUT6 #(
   .INIT(64'h7754424477544244)  
) LUT6_inst8883 (
   .O(to_level3[1107]),
   .I0(level4_in[6642]),
   .I1(level4_in[6643]),
   .I2(level4_in[6644]),
   .I3(level4_in[6645]),
   .I4(level4_in[6646]),
   .I5(level4_in[6647])
);

LUT6 #(
   .INIT(64'h4dfbd3b24dfbd3b2)  
) LUT6_inst8884 (
   .O(to_level3[1108]),
   .I0(level4_in[6648]),
   .I1(level4_in[6649]),
   .I2(level4_in[6650]),
   .I3(level4_in[6651]),
   .I4(level4_in[6652]),
   .I5(level4_in[6653])
);

LUT6 #(
   .INIT(64'h190cf7f8190cf7f8)  
) LUT6_inst8885 (
   .O(to_level3[1109]),
   .I0(level4_in[6654]),
   .I1(level4_in[6655]),
   .I2(level4_in[6656]),
   .I3(level4_in[6657]),
   .I4(level4_in[6658]),
   .I5(level4_in[6659])
);

LUT6 #(
   .INIT(64'h68d862be68d862be)  
) LUT6_inst8886 (
   .O(to_level3[1110]),
   .I0(level4_in[6660]),
   .I1(level4_in[6661]),
   .I2(level4_in[6662]),
   .I3(level4_in[6663]),
   .I4(level4_in[6664]),
   .I5(level4_in[6665])
);

LUT6 #(
   .INIT(64'h9fa5ab719fa5ab71)  
) LUT6_inst8887 (
   .O(to_level3[1111]),
   .I0(level4_in[6666]),
   .I1(level4_in[6667]),
   .I2(level4_in[6668]),
   .I3(level4_in[6669]),
   .I4(level4_in[6670]),
   .I5(level4_in[6671])
);

LUT6 #(
   .INIT(64'h9a286af99a286af9)  
) LUT6_inst8888 (
   .O(to_level3[1112]),
   .I0(level4_in[6672]),
   .I1(level4_in[6673]),
   .I2(level4_in[6674]),
   .I3(level4_in[6675]),
   .I4(level4_in[6676]),
   .I5(level4_in[6677])
);

LUT6 #(
   .INIT(64'h13d2a57913d2a579)  
) LUT6_inst8889 (
   .O(to_level3[1113]),
   .I0(level4_in[6678]),
   .I1(level4_in[6679]),
   .I2(level4_in[6680]),
   .I3(level4_in[6681]),
   .I4(level4_in[6682]),
   .I5(level4_in[6683])
);

LUT6 #(
   .INIT(64'h66a83d1466a83d14)  
) LUT6_inst8890 (
   .O(to_level3[1114]),
   .I0(level4_in[6684]),
   .I1(level4_in[6685]),
   .I2(level4_in[6686]),
   .I3(level4_in[6687]),
   .I4(level4_in[6688]),
   .I5(level4_in[6689])
);

LUT6 #(
   .INIT(64'hfb1562a7fb1562a7)  
) LUT6_inst8891 (
   .O(to_level3[1115]),
   .I0(level4_in[6690]),
   .I1(level4_in[6691]),
   .I2(level4_in[6692]),
   .I3(level4_in[6693]),
   .I4(level4_in[6694]),
   .I5(level4_in[6695])
);

LUT6 #(
   .INIT(64'hbba98221bba98221)  
) LUT6_inst8892 (
   .O(to_level3[1116]),
   .I0(level4_in[6696]),
   .I1(level4_in[6697]),
   .I2(level4_in[6698]),
   .I3(level4_in[6699]),
   .I4(level4_in[6700]),
   .I5(level4_in[6701])
);

LUT6 #(
   .INIT(64'h514ac0db514ac0db)  
) LUT6_inst8893 (
   .O(to_level3[1117]),
   .I0(level4_in[6702]),
   .I1(level4_in[6703]),
   .I2(level4_in[6704]),
   .I3(level4_in[6705]),
   .I4(level4_in[6706]),
   .I5(level4_in[6707])
);

LUT6 #(
   .INIT(64'h453a4a0c453a4a0c)  
) LUT6_inst8894 (
   .O(to_level3[1118]),
   .I0(level4_in[6708]),
   .I1(level4_in[6709]),
   .I2(level4_in[6710]),
   .I3(level4_in[6711]),
   .I4(level4_in[6712]),
   .I5(level4_in[6713])
);

LUT6 #(
   .INIT(64'hfe7e0334fe7e0334)  
) LUT6_inst8895 (
   .O(to_level3[1119]),
   .I0(level4_in[6714]),
   .I1(level4_in[6715]),
   .I2(level4_in[6716]),
   .I3(level4_in[6717]),
   .I4(level4_in[6718]),
   .I5(level4_in[6719])
);

LUT6 #(
   .INIT(64'h6f233c7c6f233c7c)  
) LUT6_inst8896 (
   .O(to_level3[1120]),
   .I0(level4_in[6720]),
   .I1(level4_in[6721]),
   .I2(level4_in[6722]),
   .I3(level4_in[6723]),
   .I4(level4_in[6724]),
   .I5(level4_in[6725])
);

LUT6 #(
   .INIT(64'h622c337e622c337e)  
) LUT6_inst8897 (
   .O(to_level3[1121]),
   .I0(level4_in[6726]),
   .I1(level4_in[6727]),
   .I2(level4_in[6728]),
   .I3(level4_in[6729]),
   .I4(level4_in[6730]),
   .I5(level4_in[6731])
);

LUT6 #(
   .INIT(64'h675c8035675c8035)  
) LUT6_inst8898 (
   .O(to_level3[1122]),
   .I0(level4_in[6732]),
   .I1(level4_in[6733]),
   .I2(level4_in[6734]),
   .I3(level4_in[6735]),
   .I4(level4_in[6736]),
   .I5(level4_in[6737])
);

LUT6 #(
   .INIT(64'h2125d6b82125d6b8)  
) LUT6_inst8899 (
   .O(to_level3[1123]),
   .I0(level4_in[6738]),
   .I1(level4_in[6739]),
   .I2(level4_in[6740]),
   .I3(level4_in[6741]),
   .I4(level4_in[6742]),
   .I5(level4_in[6743])
);

LUT6 #(
   .INIT(64'h9cba47359cba4735)  
) LUT6_inst8900 (
   .O(to_level3[1124]),
   .I0(level4_in[6744]),
   .I1(level4_in[6745]),
   .I2(level4_in[6746]),
   .I3(level4_in[6747]),
   .I4(level4_in[6748]),
   .I5(level4_in[6749])
);

LUT6 #(
   .INIT(64'hdc4c88b4dc4c88b4)  
) LUT6_inst8901 (
   .O(to_level3[1125]),
   .I0(level4_in[6750]),
   .I1(level4_in[6751]),
   .I2(level4_in[6752]),
   .I3(level4_in[6753]),
   .I4(level4_in[6754]),
   .I5(level4_in[6755])
);

LUT6 #(
   .INIT(64'h5656677056566770)  
) LUT6_inst8902 (
   .O(to_level3[1126]),
   .I0(level4_in[6756]),
   .I1(level4_in[6757]),
   .I2(level4_in[6758]),
   .I3(level4_in[6759]),
   .I4(level4_in[6760]),
   .I5(level4_in[6761])
);

LUT6 #(
   .INIT(64'h39dda64b39dda64b)  
) LUT6_inst8903 (
   .O(to_level3[1127]),
   .I0(level4_in[6762]),
   .I1(level4_in[6763]),
   .I2(level4_in[6764]),
   .I3(level4_in[6765]),
   .I4(level4_in[6766]),
   .I5(level4_in[6767])
);

LUT6 #(
   .INIT(64'h52ab048752ab0487)  
) LUT6_inst8904 (
   .O(to_level3[1128]),
   .I0(level4_in[6768]),
   .I1(level4_in[6769]),
   .I2(level4_in[6770]),
   .I3(level4_in[6771]),
   .I4(level4_in[6772]),
   .I5(level4_in[6773])
);

LUT6 #(
   .INIT(64'h5e2ad9e85e2ad9e8)  
) LUT6_inst8905 (
   .O(to_level3[1129]),
   .I0(level4_in[6774]),
   .I1(level4_in[6775]),
   .I2(level4_in[6776]),
   .I3(level4_in[6777]),
   .I4(level4_in[6778]),
   .I5(level4_in[6779])
);

LUT6 #(
   .INIT(64'hb7be4855b7be4855)  
) LUT6_inst8906 (
   .O(to_level3[1130]),
   .I0(level4_in[6780]),
   .I1(level4_in[6781]),
   .I2(level4_in[6782]),
   .I3(level4_in[6783]),
   .I4(level4_in[6784]),
   .I5(level4_in[6785])
);

LUT6 #(
   .INIT(64'hef94fe26ef94fe26)  
) LUT6_inst8907 (
   .O(to_level3[1131]),
   .I0(level4_in[6786]),
   .I1(level4_in[6787]),
   .I2(level4_in[6788]),
   .I3(level4_in[6789]),
   .I4(level4_in[6790]),
   .I5(level4_in[6791])
);

LUT6 #(
   .INIT(64'h07e4a37607e4a376)  
) LUT6_inst8908 (
   .O(to_level3[1132]),
   .I0(level4_in[6792]),
   .I1(level4_in[6793]),
   .I2(level4_in[6794]),
   .I3(level4_in[6795]),
   .I4(level4_in[6796]),
   .I5(level4_in[6797])
);

LUT6 #(
   .INIT(64'hf0931205f0931205)  
) LUT6_inst8909 (
   .O(to_level3[1133]),
   .I0(level4_in[6798]),
   .I1(level4_in[6799]),
   .I2(level4_in[6800]),
   .I3(level4_in[6801]),
   .I4(level4_in[6802]),
   .I5(level4_in[6803])
);

LUT6 #(
   .INIT(64'h64850d4164850d41)  
) LUT6_inst8910 (
   .O(to_level3[1134]),
   .I0(level4_in[6804]),
   .I1(level4_in[6805]),
   .I2(level4_in[6806]),
   .I3(level4_in[6807]),
   .I4(level4_in[6808]),
   .I5(level4_in[6809])
);

LUT6 #(
   .INIT(64'h58f4fa8858f4fa88)  
) LUT6_inst8911 (
   .O(to_level3[1135]),
   .I0(level4_in[6810]),
   .I1(level4_in[6811]),
   .I2(level4_in[6812]),
   .I3(level4_in[6813]),
   .I4(level4_in[6814]),
   .I5(level4_in[6815])
);

LUT6 #(
   .INIT(64'hecbcc7f7ecbcc7f7)  
) LUT6_inst8912 (
   .O(to_level3[1136]),
   .I0(level4_in[6816]),
   .I1(level4_in[6817]),
   .I2(level4_in[6818]),
   .I3(level4_in[6819]),
   .I4(level4_in[6820]),
   .I5(level4_in[6821])
);

LUT6 #(
   .INIT(64'ha3d0ce3da3d0ce3d)  
) LUT6_inst8913 (
   .O(to_level3[1137]),
   .I0(level4_in[6822]),
   .I1(level4_in[6823]),
   .I2(level4_in[6824]),
   .I3(level4_in[6825]),
   .I4(level4_in[6826]),
   .I5(level4_in[6827])
);

LUT6 #(
   .INIT(64'h625a20b4625a20b4)  
) LUT6_inst8914 (
   .O(to_level3[1138]),
   .I0(level4_in[6828]),
   .I1(level4_in[6829]),
   .I2(level4_in[6830]),
   .I3(level4_in[6831]),
   .I4(level4_in[6832]),
   .I5(level4_in[6833])
);

LUT6 #(
   .INIT(64'h90e6854690e68546)  
) LUT6_inst8915 (
   .O(to_level3[1139]),
   .I0(level4_in[6834]),
   .I1(level4_in[6835]),
   .I2(level4_in[6836]),
   .I3(level4_in[6837]),
   .I4(level4_in[6838]),
   .I5(level4_in[6839])
);

LUT6 #(
   .INIT(64'hb9a8d2d4b9a8d2d4)  
) LUT6_inst8916 (
   .O(to_level3[1140]),
   .I0(level4_in[6840]),
   .I1(level4_in[6841]),
   .I2(level4_in[6842]),
   .I3(level4_in[6843]),
   .I4(level4_in[6844]),
   .I5(level4_in[6845])
);

LUT6 #(
   .INIT(64'hbe770a76be770a76)  
) LUT6_inst8917 (
   .O(to_level3[1141]),
   .I0(level4_in[6846]),
   .I1(level4_in[6847]),
   .I2(level4_in[6848]),
   .I3(level4_in[6849]),
   .I4(level4_in[6850]),
   .I5(level4_in[6851])
);

LUT6 #(
   .INIT(64'hddf7daf3ddf7daf3)  
) LUT6_inst8918 (
   .O(to_level3[1142]),
   .I0(level4_in[6852]),
   .I1(level4_in[6853]),
   .I2(level4_in[6854]),
   .I3(level4_in[6855]),
   .I4(level4_in[6856]),
   .I5(level4_in[6857])
);

LUT6 #(
   .INIT(64'h0dbe1c670dbe1c67)  
) LUT6_inst8919 (
   .O(to_level3[1143]),
   .I0(level4_in[6858]),
   .I1(level4_in[6859]),
   .I2(level4_in[6860]),
   .I3(level4_in[6861]),
   .I4(level4_in[6862]),
   .I5(level4_in[6863])
);

LUT6 #(
   .INIT(64'h1fd9d5fe1fd9d5fe)  
) LUT6_inst8920 (
   .O(to_level3[1144]),
   .I0(level4_in[6864]),
   .I1(level4_in[6865]),
   .I2(level4_in[6866]),
   .I3(level4_in[6867]),
   .I4(level4_in[6868]),
   .I5(level4_in[6869])
);

LUT6 #(
   .INIT(64'h929a9299929a9299)  
) LUT6_inst8921 (
   .O(to_level3[1145]),
   .I0(level4_in[6870]),
   .I1(level4_in[6871]),
   .I2(level4_in[6872]),
   .I3(level4_in[6873]),
   .I4(level4_in[6874]),
   .I5(level4_in[6875])
);

LUT6 #(
   .INIT(64'h1c96f7481c96f748)  
) LUT6_inst8922 (
   .O(to_level3[1146]),
   .I0(level4_in[6876]),
   .I1(level4_in[6877]),
   .I2(level4_in[6878]),
   .I3(level4_in[6879]),
   .I4(level4_in[6880]),
   .I5(level4_in[6881])
);

LUT6 #(
   .INIT(64'h1b2cccb81b2cccb8)  
) LUT6_inst8923 (
   .O(to_level3[1147]),
   .I0(level4_in[6882]),
   .I1(level4_in[6883]),
   .I2(level4_in[6884]),
   .I3(level4_in[6885]),
   .I4(level4_in[6886]),
   .I5(level4_in[6887])
);

LUT6 #(
   .INIT(64'hf9cc75e7f9cc75e7)  
) LUT6_inst8924 (
   .O(to_level3[1148]),
   .I0(level4_in[6888]),
   .I1(level4_in[6889]),
   .I2(level4_in[6890]),
   .I3(level4_in[6891]),
   .I4(level4_in[6892]),
   .I5(level4_in[6893])
);

LUT6 #(
   .INIT(64'hbb891467bb891467)  
) LUT6_inst8925 (
   .O(to_level3[1149]),
   .I0(level4_in[6894]),
   .I1(level4_in[6895]),
   .I2(level4_in[6896]),
   .I3(level4_in[6897]),
   .I4(level4_in[6898]),
   .I5(level4_in[6899])
);

LUT6 #(
   .INIT(64'h7ce801bf7ce801bf)  
) LUT6_inst8926 (
   .O(to_level3[1150]),
   .I0(level4_in[6900]),
   .I1(level4_in[6901]),
   .I2(level4_in[6902]),
   .I3(level4_in[6903]),
   .I4(level4_in[6904]),
   .I5(level4_in[6905])
);

LUT6 #(
   .INIT(64'h714c72eb714c72eb)  
) LUT6_inst8927 (
   .O(to_level3[1151]),
   .I0(level4_in[6906]),
   .I1(level4_in[6907]),
   .I2(level4_in[6908]),
   .I3(level4_in[6909]),
   .I4(level4_in[6910]),
   .I5(level4_in[6911])
);

LUT6 #(
   .INIT(64'h474d0459474d0459)  
) LUT6_inst8928 (
   .O(to_level3[1152]),
   .I0(level4_in[6912]),
   .I1(level4_in[6913]),
   .I2(level4_in[6914]),
   .I3(level4_in[6915]),
   .I4(level4_in[6916]),
   .I5(level4_in[6917])
);

LUT6 #(
   .INIT(64'he94e9d92e94e9d92)  
) LUT6_inst8929 (
   .O(to_level3[1153]),
   .I0(level4_in[6918]),
   .I1(level4_in[6919]),
   .I2(level4_in[6920]),
   .I3(level4_in[6921]),
   .I4(level4_in[6922]),
   .I5(level4_in[6923])
);

LUT6 #(
   .INIT(64'hc20f466dc20f466d)  
) LUT6_inst8930 (
   .O(to_level3[1154]),
   .I0(level4_in[6924]),
   .I1(level4_in[6925]),
   .I2(level4_in[6926]),
   .I3(level4_in[6927]),
   .I4(level4_in[6928]),
   .I5(level4_in[6929])
);

LUT6 #(
   .INIT(64'hddca9c94ddca9c94)  
) LUT6_inst8931 (
   .O(to_level3[1155]),
   .I0(level4_in[6930]),
   .I1(level4_in[6931]),
   .I2(level4_in[6932]),
   .I3(level4_in[6933]),
   .I4(level4_in[6934]),
   .I5(level4_in[6935])
);

LUT6 #(
   .INIT(64'h559188af559188af)  
) LUT6_inst8932 (
   .O(to_level3[1156]),
   .I0(level4_in[6936]),
   .I1(level4_in[6937]),
   .I2(level4_in[6938]),
   .I3(level4_in[6939]),
   .I4(level4_in[6940]),
   .I5(level4_in[6941])
);

LUT6 #(
   .INIT(64'hf7f1dca3f7f1dca3)  
) LUT6_inst8933 (
   .O(to_level3[1157]),
   .I0(level4_in[6942]),
   .I1(level4_in[6943]),
   .I2(level4_in[6944]),
   .I3(level4_in[6945]),
   .I4(level4_in[6946]),
   .I5(level4_in[6947])
);

LUT6 #(
   .INIT(64'haf786028af786028)  
) LUT6_inst8934 (
   .O(to_level3[1158]),
   .I0(level4_in[6948]),
   .I1(level4_in[6949]),
   .I2(level4_in[6950]),
   .I3(level4_in[6951]),
   .I4(level4_in[6952]),
   .I5(level4_in[6953])
);

LUT6 #(
   .INIT(64'h368a496e368a496e)  
) LUT6_inst8935 (
   .O(to_level3[1159]),
   .I0(level4_in[6954]),
   .I1(level4_in[6955]),
   .I2(level4_in[6956]),
   .I3(level4_in[6957]),
   .I4(level4_in[6958]),
   .I5(level4_in[6959])
);

LUT6 #(
   .INIT(64'h748ba34c748ba34c)  
) LUT6_inst8936 (
   .O(to_level3[1160]),
   .I0(level4_in[6960]),
   .I1(level4_in[6961]),
   .I2(level4_in[6962]),
   .I3(level4_in[6963]),
   .I4(level4_in[6964]),
   .I5(level4_in[6965])
);

LUT6 #(
   .INIT(64'he9464e35e9464e35)  
) LUT6_inst8937 (
   .O(to_level3[1161]),
   .I0(level4_in[6966]),
   .I1(level4_in[6967]),
   .I2(level4_in[6968]),
   .I3(level4_in[6969]),
   .I4(level4_in[6970]),
   .I5(level4_in[6971])
);

LUT6 #(
   .INIT(64'h180b0deb180b0deb)  
) LUT6_inst8938 (
   .O(to_level3[1162]),
   .I0(level4_in[6972]),
   .I1(level4_in[6973]),
   .I2(level4_in[6974]),
   .I3(level4_in[6975]),
   .I4(level4_in[6976]),
   .I5(level4_in[6977])
);

LUT6 #(
   .INIT(64'hbbf048a7bbf048a7)  
) LUT6_inst8939 (
   .O(to_level3[1163]),
   .I0(level4_in[6978]),
   .I1(level4_in[6979]),
   .I2(level4_in[6980]),
   .I3(level4_in[6981]),
   .I4(level4_in[6982]),
   .I5(level4_in[6983])
);

LUT6 #(
   .INIT(64'h320cbd84320cbd84)  
) LUT6_inst8940 (
   .O(to_level3[1164]),
   .I0(level4_in[6984]),
   .I1(level4_in[6985]),
   .I2(level4_in[6986]),
   .I3(level4_in[6987]),
   .I4(level4_in[6988]),
   .I5(level4_in[6989])
);

LUT6 #(
   .INIT(64'hea5f1489ea5f1489)  
) LUT6_inst8941 (
   .O(to_level3[1165]),
   .I0(level4_in[6990]),
   .I1(level4_in[6991]),
   .I2(level4_in[6992]),
   .I3(level4_in[6993]),
   .I4(level4_in[6994]),
   .I5(level4_in[6995])
);

LUT6 #(
   .INIT(64'h2e103b662e103b66)  
) LUT6_inst8942 (
   .O(to_level3[1166]),
   .I0(level4_in[6996]),
   .I1(level4_in[6997]),
   .I2(level4_in[6998]),
   .I3(level4_in[6999]),
   .I4(level4_in[7000]),
   .I5(level4_in[7001])
);

LUT6 #(
   .INIT(64'h84ba08d384ba08d3)  
) LUT6_inst8943 (
   .O(to_level3[1167]),
   .I0(level4_in[7002]),
   .I1(level4_in[7003]),
   .I2(level4_in[7004]),
   .I3(level4_in[7005]),
   .I4(level4_in[7006]),
   .I5(level4_in[7007])
);

LUT6 #(
   .INIT(64'h22a0a99322a0a993)  
) LUT6_inst8944 (
   .O(to_level3[1168]),
   .I0(level4_in[7008]),
   .I1(level4_in[7009]),
   .I2(level4_in[7010]),
   .I3(level4_in[7011]),
   .I4(level4_in[7012]),
   .I5(level4_in[7013])
);

LUT6 #(
   .INIT(64'h5e98fd065e98fd06)  
) LUT6_inst8945 (
   .O(to_level3[1169]),
   .I0(level4_in[7014]),
   .I1(level4_in[7015]),
   .I2(level4_in[7016]),
   .I3(level4_in[7017]),
   .I4(level4_in[7018]),
   .I5(level4_in[7019])
);

LUT6 #(
   .INIT(64'h1a38c74e1a38c74e)  
) LUT6_inst8946 (
   .O(to_level3[1170]),
   .I0(level4_in[7020]),
   .I1(level4_in[7021]),
   .I2(level4_in[7022]),
   .I3(level4_in[7023]),
   .I4(level4_in[7024]),
   .I5(level4_in[7025])
);

LUT6 #(
   .INIT(64'h1114992911149929)  
) LUT6_inst8947 (
   .O(to_level3[1171]),
   .I0(level4_in[7026]),
   .I1(level4_in[7027]),
   .I2(level4_in[7028]),
   .I3(level4_in[7029]),
   .I4(level4_in[7030]),
   .I5(level4_in[7031])
);

LUT6 #(
   .INIT(64'h205f2e96205f2e96)  
) LUT6_inst8948 (
   .O(to_level3[1172]),
   .I0(level4_in[7032]),
   .I1(level4_in[7033]),
   .I2(level4_in[7034]),
   .I3(level4_in[7035]),
   .I4(level4_in[7036]),
   .I5(level4_in[7037])
);

LUT6 #(
   .INIT(64'ha2fc59d4a2fc59d4)  
) LUT6_inst8949 (
   .O(to_level3[1173]),
   .I0(level4_in[7038]),
   .I1(level4_in[7039]),
   .I2(level4_in[7040]),
   .I3(level4_in[7041]),
   .I4(level4_in[7042]),
   .I5(level4_in[7043])
);

LUT6 #(
   .INIT(64'h5ba23e1c5ba23e1c)  
) LUT6_inst8950 (
   .O(to_level3[1174]),
   .I0(level4_in[7044]),
   .I1(level4_in[7045]),
   .I2(level4_in[7046]),
   .I3(level4_in[7047]),
   .I4(level4_in[7048]),
   .I5(level4_in[7049])
);

LUT6 #(
   .INIT(64'hfca6bcb5fca6bcb5)  
) LUT6_inst8951 (
   .O(to_level3[1175]),
   .I0(level4_in[7050]),
   .I1(level4_in[7051]),
   .I2(level4_in[7052]),
   .I3(level4_in[7053]),
   .I4(level4_in[7054]),
   .I5(level4_in[7055])
);

LUT6 #(
   .INIT(64'h225e6381225e6381)  
) LUT6_inst8952 (
   .O(to_level3[1176]),
   .I0(level4_in[7056]),
   .I1(level4_in[7057]),
   .I2(level4_in[7058]),
   .I3(level4_in[7059]),
   .I4(level4_in[7060]),
   .I5(level4_in[7061])
);

LUT6 #(
   .INIT(64'h7b904a227b904a22)  
) LUT6_inst8953 (
   .O(to_level3[1177]),
   .I0(level4_in[7062]),
   .I1(level4_in[7063]),
   .I2(level4_in[7064]),
   .I3(level4_in[7065]),
   .I4(level4_in[7066]),
   .I5(level4_in[7067])
);

LUT6 #(
   .INIT(64'h6bea824e6bea824e)  
) LUT6_inst8954 (
   .O(to_level3[1178]),
   .I0(level4_in[7068]),
   .I1(level4_in[7069]),
   .I2(level4_in[7070]),
   .I3(level4_in[7071]),
   .I4(level4_in[7072]),
   .I5(level4_in[7073])
);

LUT6 #(
   .INIT(64'he655d1a9e655d1a9)  
) LUT6_inst8955 (
   .O(to_level3[1179]),
   .I0(level4_in[7074]),
   .I1(level4_in[7075]),
   .I2(level4_in[7076]),
   .I3(level4_in[7077]),
   .I4(level4_in[7078]),
   .I5(level4_in[7079])
);

LUT6 #(
   .INIT(64'h6460605c6460605c)  
) LUT6_inst8956 (
   .O(to_level3[1180]),
   .I0(level4_in[7080]),
   .I1(level4_in[7081]),
   .I2(level4_in[7082]),
   .I3(level4_in[7083]),
   .I4(level4_in[7084]),
   .I5(level4_in[7085])
);

LUT6 #(
   .INIT(64'h97587fe297587fe2)  
) LUT6_inst8957 (
   .O(to_level3[1181]),
   .I0(level4_in[7086]),
   .I1(level4_in[7087]),
   .I2(level4_in[7088]),
   .I3(level4_in[7089]),
   .I4(level4_in[7090]),
   .I5(level4_in[7091])
);

LUT6 #(
   .INIT(64'h0dc88f440dc88f44)  
) LUT6_inst8958 (
   .O(to_level3[1182]),
   .I0(level4_in[7092]),
   .I1(level4_in[7093]),
   .I2(level4_in[7094]),
   .I3(level4_in[7095]),
   .I4(level4_in[7096]),
   .I5(level4_in[7097])
);

LUT6 #(
   .INIT(64'hb881fae8b881fae8)  
) LUT6_inst8959 (
   .O(to_level3[1183]),
   .I0(level4_in[7098]),
   .I1(level4_in[7099]),
   .I2(level4_in[7100]),
   .I3(level4_in[7101]),
   .I4(level4_in[7102]),
   .I5(level4_in[7103])
);

LUT6 #(
   .INIT(64'h1ea2bac31ea2bac3)  
) LUT6_inst8960 (
   .O(to_level3[1184]),
   .I0(level4_in[7104]),
   .I1(level4_in[7105]),
   .I2(level4_in[7106]),
   .I3(level4_in[7107]),
   .I4(level4_in[7108]),
   .I5(level4_in[7109])
);

LUT6 #(
   .INIT(64'h0c336b1e0c336b1e)  
) LUT6_inst8961 (
   .O(to_level3[1185]),
   .I0(level4_in[7110]),
   .I1(level4_in[7111]),
   .I2(level4_in[7112]),
   .I3(level4_in[7113]),
   .I4(level4_in[7114]),
   .I5(level4_in[7115])
);

LUT6 #(
   .INIT(64'h19a0a85719a0a857)  
) LUT6_inst8962 (
   .O(to_level3[1186]),
   .I0(level4_in[7116]),
   .I1(level4_in[7117]),
   .I2(level4_in[7118]),
   .I3(level4_in[7119]),
   .I4(level4_in[7120]),
   .I5(level4_in[7121])
);

LUT6 #(
   .INIT(64'h7618c96d7618c96d)  
) LUT6_inst8963 (
   .O(to_level3[1187]),
   .I0(level4_in[7122]),
   .I1(level4_in[7123]),
   .I2(level4_in[7124]),
   .I3(level4_in[7125]),
   .I4(level4_in[7126]),
   .I5(level4_in[7127])
);

LUT6 #(
   .INIT(64'had9f9bb7ad9f9bb7)  
) LUT6_inst8964 (
   .O(to_level3[1188]),
   .I0(level4_in[7128]),
   .I1(level4_in[7129]),
   .I2(level4_in[7130]),
   .I3(level4_in[7131]),
   .I4(level4_in[7132]),
   .I5(level4_in[7133])
);

LUT6 #(
   .INIT(64'hd8bcf18fd8bcf18f)  
) LUT6_inst8965 (
   .O(to_level3[1189]),
   .I0(level4_in[7134]),
   .I1(level4_in[7135]),
   .I2(level4_in[7136]),
   .I3(level4_in[7137]),
   .I4(level4_in[7138]),
   .I5(level4_in[7139])
);

LUT6 #(
   .INIT(64'h9452fab09452fab0)  
) LUT6_inst8966 (
   .O(to_level3[1190]),
   .I0(level4_in[7140]),
   .I1(level4_in[7141]),
   .I2(level4_in[7142]),
   .I3(level4_in[7143]),
   .I4(level4_in[7144]),
   .I5(level4_in[7145])
);

LUT6 #(
   .INIT(64'h5934b0e65934b0e6)  
) LUT6_inst8967 (
   .O(to_level3[1191]),
   .I0(level4_in[7146]),
   .I1(level4_in[7147]),
   .I2(level4_in[7148]),
   .I3(level4_in[7149]),
   .I4(level4_in[7150]),
   .I5(level4_in[7151])
);

LUT6 #(
   .INIT(64'hc92dfbadc92dfbad)  
) LUT6_inst8968 (
   .O(to_level3[1192]),
   .I0(level4_in[7152]),
   .I1(level4_in[7153]),
   .I2(level4_in[7154]),
   .I3(level4_in[7155]),
   .I4(level4_in[7156]),
   .I5(level4_in[7157])
);

LUT6 #(
   .INIT(64'h53ccf2f753ccf2f7)  
) LUT6_inst8969 (
   .O(to_level3[1193]),
   .I0(level4_in[7158]),
   .I1(level4_in[7159]),
   .I2(level4_in[7160]),
   .I3(level4_in[7161]),
   .I4(level4_in[7162]),
   .I5(level4_in[7163])
);

LUT6 #(
   .INIT(64'hb7dd3960b7dd3960)  
) LUT6_inst8970 (
   .O(to_level3[1194]),
   .I0(level4_in[7164]),
   .I1(level4_in[7165]),
   .I2(level4_in[7166]),
   .I3(level4_in[7167]),
   .I4(level4_in[7168]),
   .I5(level4_in[7169])
);

LUT6 #(
   .INIT(64'hb68cc315b68cc315)  
) LUT6_inst8971 (
   .O(to_level3[1195]),
   .I0(level4_in[7170]),
   .I1(level4_in[7171]),
   .I2(level4_in[7172]),
   .I3(level4_in[7173]),
   .I4(level4_in[7174]),
   .I5(level4_in[7175])
);

LUT6 #(
   .INIT(64'h31b2634e31b2634e)  
) LUT6_inst8972 (
   .O(to_level3[1196]),
   .I0(level4_in[7176]),
   .I1(level4_in[7177]),
   .I2(level4_in[7178]),
   .I3(level4_in[7179]),
   .I4(level4_in[7180]),
   .I5(level4_in[7181])
);

LUT6 #(
   .INIT(64'hecb8b20aecb8b20a)  
) LUT6_inst8973 (
   .O(to_level3[1197]),
   .I0(level4_in[7182]),
   .I1(level4_in[7183]),
   .I2(level4_in[7184]),
   .I3(level4_in[7185]),
   .I4(level4_in[7186]),
   .I5(level4_in[7187])
);

LUT6 #(
   .INIT(64'hc8cbc469c8cbc469)  
) LUT6_inst8974 (
   .O(to_level3[1198]),
   .I0(level4_in[7188]),
   .I1(level4_in[7189]),
   .I2(level4_in[7190]),
   .I3(level4_in[7191]),
   .I4(level4_in[7192]),
   .I5(level4_in[7193])
);

LUT6 #(
   .INIT(64'h19f3a5a119f3a5a1)  
) LUT6_inst8975 (
   .O(to_level3[1199]),
   .I0(level4_in[7194]),
   .I1(level4_in[7195]),
   .I2(level4_in[7196]),
   .I3(level4_in[7197]),
   .I4(level4_in[7198]),
   .I5(level4_in[7199])
);

LUT6 #(
   .INIT(64'hccfd0de9ccfd0de9)  
) LUT6_inst8976 (
   .O(to_level3[1200]),
   .I0(level4_in[7200]),
   .I1(level4_in[7201]),
   .I2(level4_in[7202]),
   .I3(level4_in[7203]),
   .I4(level4_in[7204]),
   .I5(level4_in[7205])
);

LUT6 #(
   .INIT(64'h2b4135422b413542)  
) LUT6_inst8977 (
   .O(to_level3[1201]),
   .I0(level4_in[7206]),
   .I1(level4_in[7207]),
   .I2(level4_in[7208]),
   .I3(level4_in[7209]),
   .I4(level4_in[7210]),
   .I5(level4_in[7211])
);

LUT6 #(
   .INIT(64'h5221aeb65221aeb6)  
) LUT6_inst8978 (
   .O(to_level3[1202]),
   .I0(level4_in[7212]),
   .I1(level4_in[7213]),
   .I2(level4_in[7214]),
   .I3(level4_in[7215]),
   .I4(level4_in[7216]),
   .I5(level4_in[7217])
);

LUT6 #(
   .INIT(64'h1408a9f71408a9f7)  
) LUT6_inst8979 (
   .O(to_level3[1203]),
   .I0(level4_in[7218]),
   .I1(level4_in[7219]),
   .I2(level4_in[7220]),
   .I3(level4_in[7221]),
   .I4(level4_in[7222]),
   .I5(level4_in[7223])
);

LUT6 #(
   .INIT(64'had2ad3f1ad2ad3f1)  
) LUT6_inst8980 (
   .O(to_level3[1204]),
   .I0(level4_in[7224]),
   .I1(level4_in[7225]),
   .I2(level4_in[7226]),
   .I3(level4_in[7227]),
   .I4(level4_in[7228]),
   .I5(level4_in[7229])
);

LUT6 #(
   .INIT(64'hd2841e3cd2841e3c)  
) LUT6_inst8981 (
   .O(to_level3[1205]),
   .I0(level4_in[7230]),
   .I1(level4_in[7231]),
   .I2(level4_in[7232]),
   .I3(level4_in[7233]),
   .I4(level4_in[7234]),
   .I5(level4_in[7235])
);

LUT6 #(
   .INIT(64'h0a23a9120a23a912)  
) LUT6_inst8982 (
   .O(to_level3[1206]),
   .I0(level4_in[7236]),
   .I1(level4_in[7237]),
   .I2(level4_in[7238]),
   .I3(level4_in[7239]),
   .I4(level4_in[7240]),
   .I5(level4_in[7241])
);

LUT6 #(
   .INIT(64'h8798b4868798b486)  
) LUT6_inst8983 (
   .O(to_level3[1207]),
   .I0(level4_in[7242]),
   .I1(level4_in[7243]),
   .I2(level4_in[7244]),
   .I3(level4_in[7245]),
   .I4(level4_in[7246]),
   .I5(level4_in[7247])
);

LUT6 #(
   .INIT(64'hfbb44fcdfbb44fcd)  
) LUT6_inst8984 (
   .O(to_level3[1208]),
   .I0(level4_in[7248]),
   .I1(level4_in[7249]),
   .I2(level4_in[7250]),
   .I3(level4_in[7251]),
   .I4(level4_in[7252]),
   .I5(level4_in[7253])
);

LUT6 #(
   .INIT(64'hc80db42bc80db42b)  
) LUT6_inst8985 (
   .O(to_level3[1209]),
   .I0(level4_in[7254]),
   .I1(level4_in[7255]),
   .I2(level4_in[7256]),
   .I3(level4_in[7257]),
   .I4(level4_in[7258]),
   .I5(level4_in[7259])
);

LUT6 #(
   .INIT(64'h9db008409db00840)  
) LUT6_inst8986 (
   .O(to_level3[1210]),
   .I0(level4_in[7260]),
   .I1(level4_in[7261]),
   .I2(level4_in[7262]),
   .I3(level4_in[7263]),
   .I4(level4_in[7264]),
   .I5(level4_in[7265])
);

LUT6 #(
   .INIT(64'h65ca9c9265ca9c92)  
) LUT6_inst8987 (
   .O(to_level3[1211]),
   .I0(level4_in[7266]),
   .I1(level4_in[7267]),
   .I2(level4_in[7268]),
   .I3(level4_in[7269]),
   .I4(level4_in[7270]),
   .I5(level4_in[7271])
);

LUT6 #(
   .INIT(64'h38be8c6938be8c69)  
) LUT6_inst8988 (
   .O(to_level3[1212]),
   .I0(level4_in[7272]),
   .I1(level4_in[7273]),
   .I2(level4_in[7274]),
   .I3(level4_in[7275]),
   .I4(level4_in[7276]),
   .I5(level4_in[7277])
);

LUT6 #(
   .INIT(64'h01c11a6701c11a67)  
) LUT6_inst8989 (
   .O(to_level3[1213]),
   .I0(level4_in[7278]),
   .I1(level4_in[7279]),
   .I2(level4_in[7280]),
   .I3(level4_in[7281]),
   .I4(level4_in[7282]),
   .I5(level4_in[7283])
);

LUT6 #(
   .INIT(64'h02e4ded502e4ded5)  
) LUT6_inst8990 (
   .O(to_level3[1214]),
   .I0(level4_in[7284]),
   .I1(level4_in[7285]),
   .I2(level4_in[7286]),
   .I3(level4_in[7287]),
   .I4(level4_in[7288]),
   .I5(level4_in[7289])
);

LUT6 #(
   .INIT(64'hdd458576dd458576)  
) LUT6_inst8991 (
   .O(to_level3[1215]),
   .I0(level4_in[7290]),
   .I1(level4_in[7291]),
   .I2(level4_in[7292]),
   .I3(level4_in[7293]),
   .I4(level4_in[7294]),
   .I5(level4_in[7295])
);

LUT6 #(
   .INIT(64'hee7d87f5ee7d87f5)  
) LUT6_inst8992 (
   .O(to_level3[1216]),
   .I0(level4_in[7296]),
   .I1(level4_in[7297]),
   .I2(level4_in[7298]),
   .I3(level4_in[7299]),
   .I4(level4_in[7300]),
   .I5(level4_in[7301])
);

LUT6 #(
   .INIT(64'he505c729e505c729)  
) LUT6_inst8993 (
   .O(to_level3[1217]),
   .I0(level4_in[7302]),
   .I1(level4_in[7303]),
   .I2(level4_in[7304]),
   .I3(level4_in[7305]),
   .I4(level4_in[7306]),
   .I5(level4_in[7307])
);

LUT6 #(
   .INIT(64'h8657c05b8657c05b)  
) LUT6_inst8994 (
   .O(to_level3[1218]),
   .I0(level4_in[7308]),
   .I1(level4_in[7309]),
   .I2(level4_in[7310]),
   .I3(level4_in[7311]),
   .I4(level4_in[7312]),
   .I5(level4_in[7313])
);

LUT6 #(
   .INIT(64'h2639764e2639764e)  
) LUT6_inst8995 (
   .O(to_level3[1219]),
   .I0(level4_in[7314]),
   .I1(level4_in[7315]),
   .I2(level4_in[7316]),
   .I3(level4_in[7317]),
   .I4(level4_in[7318]),
   .I5(level4_in[7319])
);

LUT6 #(
   .INIT(64'ha0ceab75a0ceab75)  
) LUT6_inst8996 (
   .O(to_level3[1220]),
   .I0(level4_in[7320]),
   .I1(level4_in[7321]),
   .I2(level4_in[7322]),
   .I3(level4_in[7323]),
   .I4(level4_in[7324]),
   .I5(level4_in[7325])
);

LUT6 #(
   .INIT(64'ha8a81072a8a81072)  
) LUT6_inst8997 (
   .O(to_level3[1221]),
   .I0(level4_in[7326]),
   .I1(level4_in[7327]),
   .I2(level4_in[7328]),
   .I3(level4_in[7329]),
   .I4(level4_in[7330]),
   .I5(level4_in[7331])
);

LUT6 #(
   .INIT(64'h300f1033300f1033)  
) LUT6_inst8998 (
   .O(to_level3[1222]),
   .I0(level4_in[7332]),
   .I1(level4_in[7333]),
   .I2(level4_in[7334]),
   .I3(level4_in[7335]),
   .I4(level4_in[7336]),
   .I5(level4_in[7337])
);

LUT6 #(
   .INIT(64'hadf5150dadf5150d)  
) LUT6_inst8999 (
   .O(to_level3[1223]),
   .I0(level4_in[7338]),
   .I1(level4_in[7339]),
   .I2(level4_in[7340]),
   .I3(level4_in[7341]),
   .I4(level4_in[7342]),
   .I5(level4_in[7343])
);

LUT6 #(
   .INIT(64'h69cc25d369cc25d3)  
) LUT6_inst9000 (
   .O(to_level3[1224]),
   .I0(level4_in[7344]),
   .I1(level4_in[7345]),
   .I2(level4_in[7346]),
   .I3(level4_in[7347]),
   .I4(level4_in[7348]),
   .I5(level4_in[7349])
);

LUT6 #(
   .INIT(64'hd5b60d47d5b60d47)  
) LUT6_inst9001 (
   .O(to_level3[1225]),
   .I0(level4_in[7350]),
   .I1(level4_in[7351]),
   .I2(level4_in[7352]),
   .I3(level4_in[7353]),
   .I4(level4_in[7354]),
   .I5(level4_in[7355])
);

LUT6 #(
   .INIT(64'hbf4de5eebf4de5ee)  
) LUT6_inst9002 (
   .O(to_level3[1226]),
   .I0(level4_in[7356]),
   .I1(level4_in[7357]),
   .I2(level4_in[7358]),
   .I3(level4_in[7359]),
   .I4(level4_in[7360]),
   .I5(level4_in[7361])
);

LUT6 #(
   .INIT(64'h1b6299a91b6299a9)  
) LUT6_inst9003 (
   .O(to_level3[1227]),
   .I0(level4_in[7362]),
   .I1(level4_in[7363]),
   .I2(level4_in[7364]),
   .I3(level4_in[7365]),
   .I4(level4_in[7366]),
   .I5(level4_in[7367])
);

LUT6 #(
   .INIT(64'h2c2fc1cd2c2fc1cd)  
) LUT6_inst9004 (
   .O(to_level3[1228]),
   .I0(level4_in[7368]),
   .I1(level4_in[7369]),
   .I2(level4_in[7370]),
   .I3(level4_in[7371]),
   .I4(level4_in[7372]),
   .I5(level4_in[7373])
);

LUT6 #(
   .INIT(64'h10c8159010c81590)  
) LUT6_inst9005 (
   .O(to_level3[1229]),
   .I0(level4_in[7374]),
   .I1(level4_in[7375]),
   .I2(level4_in[7376]),
   .I3(level4_in[7377]),
   .I4(level4_in[7378]),
   .I5(level4_in[7379])
);

LUT6 #(
   .INIT(64'h6beea3766beea376)  
) LUT6_inst9006 (
   .O(to_level3[1230]),
   .I0(level4_in[7380]),
   .I1(level4_in[7381]),
   .I2(level4_in[7382]),
   .I3(level4_in[7383]),
   .I4(level4_in[7384]),
   .I5(level4_in[7385])
);

LUT6 #(
   .INIT(64'h20d9f90d20d9f90d)  
) LUT6_inst9007 (
   .O(to_level3[1231]),
   .I0(level4_in[7386]),
   .I1(level4_in[7387]),
   .I2(level4_in[7388]),
   .I3(level4_in[7389]),
   .I4(level4_in[7390]),
   .I5(level4_in[7391])
);

LUT6 #(
   .INIT(64'h05cc0e0405cc0e04)  
) LUT6_inst9008 (
   .O(to_level3[1232]),
   .I0(level4_in[7392]),
   .I1(level4_in[7393]),
   .I2(level4_in[7394]),
   .I3(level4_in[7395]),
   .I4(level4_in[7396]),
   .I5(level4_in[7397])
);

LUT6 #(
   .INIT(64'h53e49f2b53e49f2b)  
) LUT6_inst9009 (
   .O(to_level3[1233]),
   .I0(level4_in[7398]),
   .I1(level4_in[7399]),
   .I2(level4_in[7400]),
   .I3(level4_in[7401]),
   .I4(level4_in[7402]),
   .I5(level4_in[7403])
);

LUT6 #(
   .INIT(64'h352ed136352ed136)  
) LUT6_inst9010 (
   .O(to_level3[1234]),
   .I0(level4_in[7404]),
   .I1(level4_in[7405]),
   .I2(level4_in[7406]),
   .I3(level4_in[7407]),
   .I4(level4_in[7408]),
   .I5(level4_in[7409])
);

LUT6 #(
   .INIT(64'hb3ddcee9b3ddcee9)  
) LUT6_inst9011 (
   .O(to_level3[1235]),
   .I0(level4_in[7410]),
   .I1(level4_in[7411]),
   .I2(level4_in[7412]),
   .I3(level4_in[7413]),
   .I4(level4_in[7414]),
   .I5(level4_in[7415])
);

LUT6 #(
   .INIT(64'h6933093169330931)  
) LUT6_inst9012 (
   .O(to_level3[1236]),
   .I0(level4_in[7416]),
   .I1(level4_in[7417]),
   .I2(level4_in[7418]),
   .I3(level4_in[7419]),
   .I4(level4_in[7420]),
   .I5(level4_in[7421])
);

LUT6 #(
   .INIT(64'h765a64b9765a64b9)  
) LUT6_inst9013 (
   .O(to_level3[1237]),
   .I0(level4_in[7422]),
   .I1(level4_in[7423]),
   .I2(level4_in[7424]),
   .I3(level4_in[7425]),
   .I4(level4_in[7426]),
   .I5(level4_in[7427])
);

LUT6 #(
   .INIT(64'hf5934420f5934420)  
) LUT6_inst9014 (
   .O(to_level3[1238]),
   .I0(level4_in[7428]),
   .I1(level4_in[7429]),
   .I2(level4_in[7430]),
   .I3(level4_in[7431]),
   .I4(level4_in[7432]),
   .I5(level4_in[7433])
);

LUT6 #(
   .INIT(64'he6ad3fe2e6ad3fe2)  
) LUT6_inst9015 (
   .O(to_level3[1239]),
   .I0(level4_in[7434]),
   .I1(level4_in[7435]),
   .I2(level4_in[7436]),
   .I3(level4_in[7437]),
   .I4(level4_in[7438]),
   .I5(level4_in[7439])
);

LUT6 #(
   .INIT(64'ha41281dda41281dd)  
) LUT6_inst9016 (
   .O(to_level3[1240]),
   .I0(level4_in[7440]),
   .I1(level4_in[7441]),
   .I2(level4_in[7442]),
   .I3(level4_in[7443]),
   .I4(level4_in[7444]),
   .I5(level4_in[7445])
);

LUT6 #(
   .INIT(64'ha3fb2cd1a3fb2cd1)  
) LUT6_inst9017 (
   .O(to_level3[1241]),
   .I0(level4_in[7446]),
   .I1(level4_in[7447]),
   .I2(level4_in[7448]),
   .I3(level4_in[7449]),
   .I4(level4_in[7450]),
   .I5(level4_in[7451])
);

LUT6 #(
   .INIT(64'had30a449ad30a449)  
) LUT6_inst9018 (
   .O(to_level3[1242]),
   .I0(level4_in[7452]),
   .I1(level4_in[7453]),
   .I2(level4_in[7454]),
   .I3(level4_in[7455]),
   .I4(level4_in[7456]),
   .I5(level4_in[7457])
);

LUT6 #(
   .INIT(64'he3a747bfe3a747bf)  
) LUT6_inst9019 (
   .O(to_level3[1243]),
   .I0(level4_in[7458]),
   .I1(level4_in[7459]),
   .I2(level4_in[7460]),
   .I3(level4_in[7461]),
   .I4(level4_in[7462]),
   .I5(level4_in[7463])
);

LUT6 #(
   .INIT(64'h9dc1f6589dc1f658)  
) LUT6_inst9020 (
   .O(to_level3[1244]),
   .I0(level4_in[7464]),
   .I1(level4_in[7465]),
   .I2(level4_in[7466]),
   .I3(level4_in[7467]),
   .I4(level4_in[7468]),
   .I5(level4_in[7469])
);

LUT6 #(
   .INIT(64'h310f001e310f001e)  
) LUT6_inst9021 (
   .O(to_level3[1245]),
   .I0(level4_in[7470]),
   .I1(level4_in[7471]),
   .I2(level4_in[7472]),
   .I3(level4_in[7473]),
   .I4(level4_in[7474]),
   .I5(level4_in[7475])
);

LUT6 #(
   .INIT(64'h9676287b9676287b)  
) LUT6_inst9022 (
   .O(to_level3[1246]),
   .I0(level4_in[7476]),
   .I1(level4_in[7477]),
   .I2(level4_in[7478]),
   .I3(level4_in[7479]),
   .I4(level4_in[7480]),
   .I5(level4_in[7481])
);

LUT6 #(
   .INIT(64'h1ac36ebe1ac36ebe)  
) LUT6_inst9023 (
   .O(to_level3[1247]),
   .I0(level4_in[7482]),
   .I1(level4_in[7483]),
   .I2(level4_in[7484]),
   .I3(level4_in[7485]),
   .I4(level4_in[7486]),
   .I5(level4_in[7487])
);

LUT6 #(
   .INIT(64'hd2d77608d2d77608)  
) LUT6_inst9024 (
   .O(to_level3[1248]),
   .I0(level4_in[7488]),
   .I1(level4_in[7489]),
   .I2(level4_in[7490]),
   .I3(level4_in[7491]),
   .I4(level4_in[7492]),
   .I5(level4_in[7493])
);

LUT6 #(
   .INIT(64'h9fffeade9fffeade)  
) LUT6_inst9025 (
   .O(to_level3[1249]),
   .I0(level4_in[7494]),
   .I1(level4_in[7495]),
   .I2(level4_in[7496]),
   .I3(level4_in[7497]),
   .I4(level4_in[7498]),
   .I5(level4_in[7499])
);

LUT6 #(
   .INIT(64'h2230c8652230c865)  
) LUT6_inst9026 (
   .O(to_level3[1250]),
   .I0(level4_in[7500]),
   .I1(level4_in[7501]),
   .I2(level4_in[7502]),
   .I3(level4_in[7503]),
   .I4(level4_in[7504]),
   .I5(level4_in[7505])
);

LUT6 #(
   .INIT(64'h0747de510747de51)  
) LUT6_inst9027 (
   .O(to_level3[1251]),
   .I0(level4_in[7506]),
   .I1(level4_in[7507]),
   .I2(level4_in[7508]),
   .I3(level4_in[7509]),
   .I4(level4_in[7510]),
   .I5(level4_in[7511])
);

LUT6 #(
   .INIT(64'h6837c2246837c224)  
) LUT6_inst9028 (
   .O(to_level3[1252]),
   .I0(level4_in[7512]),
   .I1(level4_in[7513]),
   .I2(level4_in[7514]),
   .I3(level4_in[7515]),
   .I4(level4_in[7516]),
   .I5(level4_in[7517])
);

LUT6 #(
   .INIT(64'h62ef558762ef5587)  
) LUT6_inst9029 (
   .O(to_level3[1253]),
   .I0(level4_in[7518]),
   .I1(level4_in[7519]),
   .I2(level4_in[7520]),
   .I3(level4_in[7521]),
   .I4(level4_in[7522]),
   .I5(level4_in[7523])
);

LUT6 #(
   .INIT(64'hcda90be9cda90be9)  
) LUT6_inst9030 (
   .O(to_level3[1254]),
   .I0(level4_in[7524]),
   .I1(level4_in[7525]),
   .I2(level4_in[7526]),
   .I3(level4_in[7527]),
   .I4(level4_in[7528]),
   .I5(level4_in[7529])
);

LUT6 #(
   .INIT(64'h5be581cd5be581cd)  
) LUT6_inst9031 (
   .O(to_level3[1255]),
   .I0(level4_in[7530]),
   .I1(level4_in[7531]),
   .I2(level4_in[7532]),
   .I3(level4_in[7533]),
   .I4(level4_in[7534]),
   .I5(level4_in[7535])
);

LUT6 #(
   .INIT(64'h7e714ad97e714ad9)  
) LUT6_inst9032 (
   .O(to_level3[1256]),
   .I0(level4_in[7536]),
   .I1(level4_in[7537]),
   .I2(level4_in[7538]),
   .I3(level4_in[7539]),
   .I4(level4_in[7540]),
   .I5(level4_in[7541])
);

LUT6 #(
   .INIT(64'h7b3e8b507b3e8b50)  
) LUT6_inst9033 (
   .O(to_level3[1257]),
   .I0(level4_in[7542]),
   .I1(level4_in[7543]),
   .I2(level4_in[7544]),
   .I3(level4_in[7545]),
   .I4(level4_in[7546]),
   .I5(level4_in[7547])
);

LUT6 #(
   .INIT(64'h29543c7029543c70)  
) LUT6_inst9034 (
   .O(to_level3[1258]),
   .I0(level4_in[7548]),
   .I1(level4_in[7549]),
   .I2(level4_in[7550]),
   .I3(level4_in[7551]),
   .I4(level4_in[7552]),
   .I5(level4_in[7553])
);

LUT6 #(
   .INIT(64'hf4cce45df4cce45d)  
) LUT6_inst9035 (
   .O(to_level3[1259]),
   .I0(level4_in[7554]),
   .I1(level4_in[7555]),
   .I2(level4_in[7556]),
   .I3(level4_in[7557]),
   .I4(level4_in[7558]),
   .I5(level4_in[7559])
);

LUT6 #(
   .INIT(64'h2e6e002b2e6e002b)  
) LUT6_inst9036 (
   .O(to_level3[1260]),
   .I0(level4_in[7560]),
   .I1(level4_in[7561]),
   .I2(level4_in[7562]),
   .I3(level4_in[7563]),
   .I4(level4_in[7564]),
   .I5(level4_in[7565])
);

LUT6 #(
   .INIT(64'h90ba586690ba5866)  
) LUT6_inst9037 (
   .O(to_level3[1261]),
   .I0(level4_in[7566]),
   .I1(level4_in[7567]),
   .I2(level4_in[7568]),
   .I3(level4_in[7569]),
   .I4(level4_in[7570]),
   .I5(level4_in[7571])
);

LUT6 #(
   .INIT(64'h327522b4327522b4)  
) LUT6_inst9038 (
   .O(to_level3[1262]),
   .I0(level4_in[7572]),
   .I1(level4_in[7573]),
   .I2(level4_in[7574]),
   .I3(level4_in[7575]),
   .I4(level4_in[7576]),
   .I5(level4_in[7577])
);

LUT6 #(
   .INIT(64'hc4662010c4662010)  
) LUT6_inst9039 (
   .O(to_level3[1263]),
   .I0(level4_in[7578]),
   .I1(level4_in[7579]),
   .I2(level4_in[7580]),
   .I3(level4_in[7581]),
   .I4(level4_in[7582]),
   .I5(level4_in[7583])
);

LUT6 #(
   .INIT(64'hf539b50ef539b50e)  
) LUT6_inst9040 (
   .O(to_level3[1264]),
   .I0(level4_in[7584]),
   .I1(level4_in[7585]),
   .I2(level4_in[7586]),
   .I3(level4_in[7587]),
   .I4(level4_in[7588]),
   .I5(level4_in[7589])
);

LUT6 #(
   .INIT(64'he19b36cbe19b36cb)  
) LUT6_inst9041 (
   .O(to_level3[1265]),
   .I0(level4_in[7590]),
   .I1(level4_in[7591]),
   .I2(level4_in[7592]),
   .I3(level4_in[7593]),
   .I4(level4_in[7594]),
   .I5(level4_in[7595])
);

LUT6 #(
   .INIT(64'hed6a79e8ed6a79e8)  
) LUT6_inst9042 (
   .O(to_level3[1266]),
   .I0(level4_in[7596]),
   .I1(level4_in[7597]),
   .I2(level4_in[7598]),
   .I3(level4_in[7599]),
   .I4(level4_in[7600]),
   .I5(level4_in[7601])
);

LUT6 #(
   .INIT(64'h18ab220b18ab220b)  
) LUT6_inst9043 (
   .O(to_level3[1267]),
   .I0(level4_in[7602]),
   .I1(level4_in[7603]),
   .I2(level4_in[7604]),
   .I3(level4_in[7605]),
   .I4(level4_in[7606]),
   .I5(level4_in[7607])
);

LUT6 #(
   .INIT(64'h7ea5cb5d7ea5cb5d)  
) LUT6_inst9044 (
   .O(to_level3[1268]),
   .I0(level4_in[7608]),
   .I1(level4_in[7609]),
   .I2(level4_in[7610]),
   .I3(level4_in[7611]),
   .I4(level4_in[7612]),
   .I5(level4_in[7613])
);

LUT6 #(
   .INIT(64'ha8985364a8985364)  
) LUT6_inst9045 (
   .O(to_level3[1269]),
   .I0(level4_in[7614]),
   .I1(level4_in[7615]),
   .I2(level4_in[7616]),
   .I3(level4_in[7617]),
   .I4(level4_in[7618]),
   .I5(level4_in[7619])
);

LUT6 #(
   .INIT(64'h57fc4a7e57fc4a7e)  
) LUT6_inst9046 (
   .O(to_level3[1270]),
   .I0(level4_in[7620]),
   .I1(level4_in[7621]),
   .I2(level4_in[7622]),
   .I3(level4_in[7623]),
   .I4(level4_in[7624]),
   .I5(level4_in[7625])
);

LUT6 #(
   .INIT(64'h25f0571425f05714)  
) LUT6_inst9047 (
   .O(to_level3[1271]),
   .I0(level4_in[7626]),
   .I1(level4_in[7627]),
   .I2(level4_in[7628]),
   .I3(level4_in[7629]),
   .I4(level4_in[7630]),
   .I5(level4_in[7631])
);

LUT6 #(
   .INIT(64'h59a345d959a345d9)  
) LUT6_inst9048 (
   .O(to_level3[1272]),
   .I0(level4_in[7632]),
   .I1(level4_in[7633]),
   .I2(level4_in[7634]),
   .I3(level4_in[7635]),
   .I4(level4_in[7636]),
   .I5(level4_in[7637])
);

LUT6 #(
   .INIT(64'h46939a4c46939a4c)  
) LUT6_inst9049 (
   .O(to_level3[1273]),
   .I0(level4_in[7638]),
   .I1(level4_in[7639]),
   .I2(level4_in[7640]),
   .I3(level4_in[7641]),
   .I4(level4_in[7642]),
   .I5(level4_in[7643])
);

LUT6 #(
   .INIT(64'hd4757082d4757082)  
) LUT6_inst9050 (
   .O(to_level3[1274]),
   .I0(level4_in[7644]),
   .I1(level4_in[7645]),
   .I2(level4_in[7646]),
   .I3(level4_in[7647]),
   .I4(level4_in[7648]),
   .I5(level4_in[7649])
);

LUT6 #(
   .INIT(64'h6904ec196904ec19)  
) LUT6_inst9051 (
   .O(to_level3[1275]),
   .I0(level4_in[7650]),
   .I1(level4_in[7651]),
   .I2(level4_in[7652]),
   .I3(level4_in[7653]),
   .I4(level4_in[7654]),
   .I5(level4_in[7655])
);

LUT6 #(
   .INIT(64'h8ec2c5338ec2c533)  
) LUT6_inst9052 (
   .O(to_level3[1276]),
   .I0(level4_in[7656]),
   .I1(level4_in[7657]),
   .I2(level4_in[7658]),
   .I3(level4_in[7659]),
   .I4(level4_in[7660]),
   .I5(level4_in[7661])
);

LUT6 #(
   .INIT(64'h432b6a02432b6a02)  
) LUT6_inst9053 (
   .O(to_level3[1277]),
   .I0(level4_in[7662]),
   .I1(level4_in[7663]),
   .I2(level4_in[7664]),
   .I3(level4_in[7665]),
   .I4(level4_in[7666]),
   .I5(level4_in[7667])
);

LUT6 #(
   .INIT(64'he2989741e2989741)  
) LUT6_inst9054 (
   .O(to_level3[1278]),
   .I0(level4_in[7668]),
   .I1(level4_in[7669]),
   .I2(level4_in[7670]),
   .I3(level4_in[7671]),
   .I4(level4_in[7672]),
   .I5(level4_in[7673])
);

LUT6 #(
   .INIT(64'h78f5adbb78f5adbb)  
) LUT6_inst9055 (
   .O(to_level3[1279]),
   .I0(level4_in[7674]),
   .I1(level4_in[7675]),
   .I2(level4_in[7676]),
   .I3(level4_in[7677]),
   .I4(level4_in[7678]),
   .I5(level4_in[7679])
);

LUT6 #(
   .INIT(64'h02dcb00602dcb006)  
) LUT6_inst9056 (
   .O(to_level3[1280]),
   .I0(level4_in[7680]),
   .I1(level4_in[7681]),
   .I2(level4_in[7682]),
   .I3(level4_in[7683]),
   .I4(level4_in[7684]),
   .I5(level4_in[7685])
);

LUT6 #(
   .INIT(64'h530bd058530bd058)  
) LUT6_inst9057 (
   .O(to_level3[1281]),
   .I0(level4_in[7686]),
   .I1(level4_in[7687]),
   .I2(level4_in[7688]),
   .I3(level4_in[7689]),
   .I4(level4_in[7690]),
   .I5(level4_in[7691])
);

LUT6 #(
   .INIT(64'h1865cabd1865cabd)  
) LUT6_inst9058 (
   .O(to_level3[1282]),
   .I0(level4_in[7692]),
   .I1(level4_in[7693]),
   .I2(level4_in[7694]),
   .I3(level4_in[7695]),
   .I4(level4_in[7696]),
   .I5(level4_in[7697])
);

LUT6 #(
   .INIT(64'h226c0aaf226c0aaf)  
) LUT6_inst9059 (
   .O(to_level3[1283]),
   .I0(level4_in[7698]),
   .I1(level4_in[7699]),
   .I2(level4_in[7700]),
   .I3(level4_in[7701]),
   .I4(level4_in[7702]),
   .I5(level4_in[7703])
);

LUT6 #(
   .INIT(64'h1d2609cd1d2609cd)  
) LUT6_inst9060 (
   .O(to_level3[1284]),
   .I0(level4_in[7704]),
   .I1(level4_in[7705]),
   .I2(level4_in[7706]),
   .I3(level4_in[7707]),
   .I4(level4_in[7708]),
   .I5(level4_in[7709])
);

LUT6 #(
   .INIT(64'h509ad9e7509ad9e7)  
) LUT6_inst9061 (
   .O(to_level3[1285]),
   .I0(level4_in[7710]),
   .I1(level4_in[7711]),
   .I2(level4_in[7712]),
   .I3(level4_in[7713]),
   .I4(level4_in[7714]),
   .I5(level4_in[7715])
);

LUT6 #(
   .INIT(64'h4459d6ce4459d6ce)  
) LUT6_inst9062 (
   .O(to_level3[1286]),
   .I0(level4_in[7716]),
   .I1(level4_in[7717]),
   .I2(level4_in[7718]),
   .I3(level4_in[7719]),
   .I4(level4_in[7720]),
   .I5(level4_in[7721])
);

LUT6 #(
   .INIT(64'h7e201f607e201f60)  
) LUT6_inst9063 (
   .O(to_level3[1287]),
   .I0(level4_in[7722]),
   .I1(level4_in[7723]),
   .I2(level4_in[7724]),
   .I3(level4_in[7725]),
   .I4(level4_in[7726]),
   .I5(level4_in[7727])
);

LUT6 #(
   .INIT(64'h046576da046576da)  
) LUT6_inst9064 (
   .O(to_level3[1288]),
   .I0(level4_in[7728]),
   .I1(level4_in[7729]),
   .I2(level4_in[7730]),
   .I3(level4_in[7731]),
   .I4(level4_in[7732]),
   .I5(level4_in[7733])
);

LUT6 #(
   .INIT(64'h5d6eb62c5d6eb62c)  
) LUT6_inst9065 (
   .O(to_level3[1289]),
   .I0(level4_in[7734]),
   .I1(level4_in[7735]),
   .I2(level4_in[7736]),
   .I3(level4_in[7737]),
   .I4(level4_in[7738]),
   .I5(level4_in[7739])
);

LUT6 #(
   .INIT(64'h4f4e576f4f4e576f)  
) LUT6_inst9066 (
   .O(to_level3[1290]),
   .I0(level4_in[7740]),
   .I1(level4_in[7741]),
   .I2(level4_in[7742]),
   .I3(level4_in[7743]),
   .I4(level4_in[7744]),
   .I5(level4_in[7745])
);

LUT6 #(
   .INIT(64'h5ab3bd6c5ab3bd6c)  
) LUT6_inst9067 (
   .O(to_level3[1291]),
   .I0(level4_in[7746]),
   .I1(level4_in[7747]),
   .I2(level4_in[7748]),
   .I3(level4_in[7749]),
   .I4(level4_in[7750]),
   .I5(level4_in[7751])
);

LUT6 #(
   .INIT(64'h51a83a8251a83a82)  
) LUT6_inst9068 (
   .O(to_level3[1292]),
   .I0(level4_in[7752]),
   .I1(level4_in[7753]),
   .I2(level4_in[7754]),
   .I3(level4_in[7755]),
   .I4(level4_in[7756]),
   .I5(level4_in[7757])
);

LUT6 #(
   .INIT(64'h7697947776979477)  
) LUT6_inst9069 (
   .O(to_level3[1293]),
   .I0(level4_in[7758]),
   .I1(level4_in[7759]),
   .I2(level4_in[7760]),
   .I3(level4_in[7761]),
   .I4(level4_in[7762]),
   .I5(level4_in[7763])
);

LUT6 #(
   .INIT(64'h46a94b2046a94b20)  
) LUT6_inst9070 (
   .O(to_level3[1294]),
   .I0(level4_in[7764]),
   .I1(level4_in[7765]),
   .I2(level4_in[7766]),
   .I3(level4_in[7767]),
   .I4(level4_in[7768]),
   .I5(level4_in[7769])
);

LUT6 #(
   .INIT(64'h3fd443053fd44305)  
) LUT6_inst9071 (
   .O(to_level3[1295]),
   .I0(level4_in[7770]),
   .I1(level4_in[7771]),
   .I2(level4_in[7772]),
   .I3(level4_in[7773]),
   .I4(level4_in[7774]),
   .I5(level4_in[7775])
);
////////////// level 3 starts below:/n
LUT6 #(
   .INIT(64'hb86c5c00b86c5c00)  
) LUT6_inst9072 (
   .O(to_level2[0]),
   .I0(level3_in[0]),
   .I1(level3_in[1]),
   .I2(level3_in[2]),
   .I3(level3_in[3]),
   .I4(level3_in[4]),
   .I5(level3_in[5])
);

LUT6 #(
   .INIT(64'h0e91443d0e91443d)  
) LUT6_inst9073 (
   .O(to_level2[1]),
   .I0(level3_in[6]),
   .I1(level3_in[7]),
   .I2(level3_in[8]),
   .I3(level3_in[9]),
   .I4(level3_in[10]),
   .I5(level3_in[11])
);

LUT6 #(
   .INIT(64'h74fd90d574fd90d5)  
) LUT6_inst9074 (
   .O(to_level2[2]),
   .I0(level3_in[12]),
   .I1(level3_in[13]),
   .I2(level3_in[14]),
   .I3(level3_in[15]),
   .I4(level3_in[16]),
   .I5(level3_in[17])
);

LUT6 #(
   .INIT(64'h5d9ed0955d9ed095)  
) LUT6_inst9075 (
   .O(to_level2[3]),
   .I0(level3_in[18]),
   .I1(level3_in[19]),
   .I2(level3_in[20]),
   .I3(level3_in[21]),
   .I4(level3_in[22]),
   .I5(level3_in[23])
);

LUT6 #(
   .INIT(64'h0798627207986272)  
) LUT6_inst9076 (
   .O(to_level2[4]),
   .I0(level3_in[24]),
   .I1(level3_in[25]),
   .I2(level3_in[26]),
   .I3(level3_in[27]),
   .I4(level3_in[28]),
   .I5(level3_in[29])
);

LUT6 #(
   .INIT(64'h9348168893481688)  
) LUT6_inst9077 (
   .O(to_level2[5]),
   .I0(level3_in[30]),
   .I1(level3_in[31]),
   .I2(level3_in[32]),
   .I3(level3_in[33]),
   .I4(level3_in[34]),
   .I5(level3_in[35])
);

LUT6 #(
   .INIT(64'h387ab408387ab408)  
) LUT6_inst9078 (
   .O(to_level2[6]),
   .I0(level3_in[36]),
   .I1(level3_in[37]),
   .I2(level3_in[38]),
   .I3(level3_in[39]),
   .I4(level3_in[40]),
   .I5(level3_in[41])
);

LUT6 #(
   .INIT(64'h6eba36276eba3627)  
) LUT6_inst9079 (
   .O(to_level2[7]),
   .I0(level3_in[42]),
   .I1(level3_in[43]),
   .I2(level3_in[44]),
   .I3(level3_in[45]),
   .I4(level3_in[46]),
   .I5(level3_in[47])
);

LUT6 #(
   .INIT(64'h2172a3ec2172a3ec)  
) LUT6_inst9080 (
   .O(to_level2[8]),
   .I0(level3_in[48]),
   .I1(level3_in[49]),
   .I2(level3_in[50]),
   .I3(level3_in[51]),
   .I4(level3_in[52]),
   .I5(level3_in[53])
);

LUT6 #(
   .INIT(64'hbaf13b87baf13b87)  
) LUT6_inst9081 (
   .O(to_level2[9]),
   .I0(level3_in[54]),
   .I1(level3_in[55]),
   .I2(level3_in[56]),
   .I3(level3_in[57]),
   .I4(level3_in[58]),
   .I5(level3_in[59])
);

LUT6 #(
   .INIT(64'h2ba9a6162ba9a616)  
) LUT6_inst9082 (
   .O(to_level2[10]),
   .I0(level3_in[60]),
   .I1(level3_in[61]),
   .I2(level3_in[62]),
   .I3(level3_in[63]),
   .I4(level3_in[64]),
   .I5(level3_in[65])
);

LUT6 #(
   .INIT(64'h011cb5db011cb5db)  
) LUT6_inst9083 (
   .O(to_level2[11]),
   .I0(level3_in[66]),
   .I1(level3_in[67]),
   .I2(level3_in[68]),
   .I3(level3_in[69]),
   .I4(level3_in[70]),
   .I5(level3_in[71])
);

LUT6 #(
   .INIT(64'h45cc252545cc2525)  
) LUT6_inst9084 (
   .O(to_level2[12]),
   .I0(level3_in[72]),
   .I1(level3_in[73]),
   .I2(level3_in[74]),
   .I3(level3_in[75]),
   .I4(level3_in[76]),
   .I5(level3_in[77])
);

LUT6 #(
   .INIT(64'h405f535c405f535c)  
) LUT6_inst9085 (
   .O(to_level2[13]),
   .I0(level3_in[78]),
   .I1(level3_in[79]),
   .I2(level3_in[80]),
   .I3(level3_in[81]),
   .I4(level3_in[82]),
   .I5(level3_in[83])
);

LUT6 #(
   .INIT(64'hf1543571f1543571)  
) LUT6_inst9086 (
   .O(to_level2[14]),
   .I0(level3_in[84]),
   .I1(level3_in[85]),
   .I2(level3_in[86]),
   .I3(level3_in[87]),
   .I4(level3_in[88]),
   .I5(level3_in[89])
);

LUT6 #(
   .INIT(64'h22256ea722256ea7)  
) LUT6_inst9087 (
   .O(to_level2[15]),
   .I0(level3_in[90]),
   .I1(level3_in[91]),
   .I2(level3_in[92]),
   .I3(level3_in[93]),
   .I4(level3_in[94]),
   .I5(level3_in[95])
);

LUT6 #(
   .INIT(64'ha9a4601aa9a4601a)  
) LUT6_inst9088 (
   .O(to_level2[16]),
   .I0(level3_in[96]),
   .I1(level3_in[97]),
   .I2(level3_in[98]),
   .I3(level3_in[99]),
   .I4(level3_in[100]),
   .I5(level3_in[101])
);

LUT6 #(
   .INIT(64'h2c72c1c02c72c1c0)  
) LUT6_inst9089 (
   .O(to_level2[17]),
   .I0(level3_in[102]),
   .I1(level3_in[103]),
   .I2(level3_in[104]),
   .I3(level3_in[105]),
   .I4(level3_in[106]),
   .I5(level3_in[107])
);

LUT6 #(
   .INIT(64'h82ffe06f82ffe06f)  
) LUT6_inst9090 (
   .O(to_level2[18]),
   .I0(level3_in[108]),
   .I1(level3_in[109]),
   .I2(level3_in[110]),
   .I3(level3_in[111]),
   .I4(level3_in[112]),
   .I5(level3_in[113])
);

LUT6 #(
   .INIT(64'hc3a30464c3a30464)  
) LUT6_inst9091 (
   .O(to_level2[19]),
   .I0(level3_in[114]),
   .I1(level3_in[115]),
   .I2(level3_in[116]),
   .I3(level3_in[117]),
   .I4(level3_in[118]),
   .I5(level3_in[119])
);

LUT6 #(
   .INIT(64'hcba4ac8bcba4ac8b)  
) LUT6_inst9092 (
   .O(to_level2[20]),
   .I0(level3_in[120]),
   .I1(level3_in[121]),
   .I2(level3_in[122]),
   .I3(level3_in[123]),
   .I4(level3_in[124]),
   .I5(level3_in[125])
);

LUT6 #(
   .INIT(64'h8bd5a6bd8bd5a6bd)  
) LUT6_inst9093 (
   .O(to_level2[21]),
   .I0(level3_in[126]),
   .I1(level3_in[127]),
   .I2(level3_in[128]),
   .I3(level3_in[129]),
   .I4(level3_in[130]),
   .I5(level3_in[131])
);

LUT6 #(
   .INIT(64'hd13aaa1cd13aaa1c)  
) LUT6_inst9094 (
   .O(to_level2[22]),
   .I0(level3_in[132]),
   .I1(level3_in[133]),
   .I2(level3_in[134]),
   .I3(level3_in[135]),
   .I4(level3_in[136]),
   .I5(level3_in[137])
);

LUT6 #(
   .INIT(64'h2ee0f9e02ee0f9e0)  
) LUT6_inst9095 (
   .O(to_level2[23]),
   .I0(level3_in[138]),
   .I1(level3_in[139]),
   .I2(level3_in[140]),
   .I3(level3_in[141]),
   .I4(level3_in[142]),
   .I5(level3_in[143])
);

LUT6 #(
   .INIT(64'h4294d1fe4294d1fe)  
) LUT6_inst9096 (
   .O(to_level2[24]),
   .I0(level3_in[144]),
   .I1(level3_in[145]),
   .I2(level3_in[146]),
   .I3(level3_in[147]),
   .I4(level3_in[148]),
   .I5(level3_in[149])
);

LUT6 #(
   .INIT(64'ha67096f4a67096f4)  
) LUT6_inst9097 (
   .O(to_level2[25]),
   .I0(level3_in[150]),
   .I1(level3_in[151]),
   .I2(level3_in[152]),
   .I3(level3_in[153]),
   .I4(level3_in[154]),
   .I5(level3_in[155])
);

LUT6 #(
   .INIT(64'h2b3351a62b3351a6)  
) LUT6_inst9098 (
   .O(to_level2[26]),
   .I0(level3_in[156]),
   .I1(level3_in[157]),
   .I2(level3_in[158]),
   .I3(level3_in[159]),
   .I4(level3_in[160]),
   .I5(level3_in[161])
);

LUT6 #(
   .INIT(64'h886230ef886230ef)  
) LUT6_inst9099 (
   .O(to_level2[27]),
   .I0(level3_in[162]),
   .I1(level3_in[163]),
   .I2(level3_in[164]),
   .I3(level3_in[165]),
   .I4(level3_in[166]),
   .I5(level3_in[167])
);

LUT6 #(
   .INIT(64'heef88a1ceef88a1c)  
) LUT6_inst9100 (
   .O(to_level2[28]),
   .I0(level3_in[168]),
   .I1(level3_in[169]),
   .I2(level3_in[170]),
   .I3(level3_in[171]),
   .I4(level3_in[172]),
   .I5(level3_in[173])
);

LUT6 #(
   .INIT(64'hec99f40bec99f40b)  
) LUT6_inst9101 (
   .O(to_level2[29]),
   .I0(level3_in[174]),
   .I1(level3_in[175]),
   .I2(level3_in[176]),
   .I3(level3_in[177]),
   .I4(level3_in[178]),
   .I5(level3_in[179])
);

LUT6 #(
   .INIT(64'hb2843813b2843813)  
) LUT6_inst9102 (
   .O(to_level2[30]),
   .I0(level3_in[180]),
   .I1(level3_in[181]),
   .I2(level3_in[182]),
   .I3(level3_in[183]),
   .I4(level3_in[184]),
   .I5(level3_in[185])
);

LUT6 #(
   .INIT(64'h7b3c7cf67b3c7cf6)  
) LUT6_inst9103 (
   .O(to_level2[31]),
   .I0(level3_in[186]),
   .I1(level3_in[187]),
   .I2(level3_in[188]),
   .I3(level3_in[189]),
   .I4(level3_in[190]),
   .I5(level3_in[191])
);

LUT6 #(
   .INIT(64'h776fef34776fef34)  
) LUT6_inst9104 (
   .O(to_level2[32]),
   .I0(level3_in[192]),
   .I1(level3_in[193]),
   .I2(level3_in[194]),
   .I3(level3_in[195]),
   .I4(level3_in[196]),
   .I5(level3_in[197])
);

LUT6 #(
   .INIT(64'hd5e0d399d5e0d399)  
) LUT6_inst9105 (
   .O(to_level2[33]),
   .I0(level3_in[198]),
   .I1(level3_in[199]),
   .I2(level3_in[200]),
   .I3(level3_in[201]),
   .I4(level3_in[202]),
   .I5(level3_in[203])
);

LUT6 #(
   .INIT(64'h0314704903147049)  
) LUT6_inst9106 (
   .O(to_level2[34]),
   .I0(level3_in[204]),
   .I1(level3_in[205]),
   .I2(level3_in[206]),
   .I3(level3_in[207]),
   .I4(level3_in[208]),
   .I5(level3_in[209])
);

LUT6 #(
   .INIT(64'h9dcf02929dcf0292)  
) LUT6_inst9107 (
   .O(to_level2[35]),
   .I0(level3_in[210]),
   .I1(level3_in[211]),
   .I2(level3_in[212]),
   .I3(level3_in[213]),
   .I4(level3_in[214]),
   .I5(level3_in[215])
);

LUT6 #(
   .INIT(64'h2d17dad82d17dad8)  
) LUT6_inst9108 (
   .O(to_level2[36]),
   .I0(level3_in[216]),
   .I1(level3_in[217]),
   .I2(level3_in[218]),
   .I3(level3_in[219]),
   .I4(level3_in[220]),
   .I5(level3_in[221])
);

LUT6 #(
   .INIT(64'h51a4c81e51a4c81e)  
) LUT6_inst9109 (
   .O(to_level2[37]),
   .I0(level3_in[222]),
   .I1(level3_in[223]),
   .I2(level3_in[224]),
   .I3(level3_in[225]),
   .I4(level3_in[226]),
   .I5(level3_in[227])
);

LUT6 #(
   .INIT(64'hc345bc07c345bc07)  
) LUT6_inst9110 (
   .O(to_level2[38]),
   .I0(level3_in[228]),
   .I1(level3_in[229]),
   .I2(level3_in[230]),
   .I3(level3_in[231]),
   .I4(level3_in[232]),
   .I5(level3_in[233])
);

LUT6 #(
   .INIT(64'hc9f5e533c9f5e533)  
) LUT6_inst9111 (
   .O(to_level2[39]),
   .I0(level3_in[234]),
   .I1(level3_in[235]),
   .I2(level3_in[236]),
   .I3(level3_in[237]),
   .I4(level3_in[238]),
   .I5(level3_in[239])
);

LUT6 #(
   .INIT(64'h29a8d62f29a8d62f)  
) LUT6_inst9112 (
   .O(to_level2[40]),
   .I0(level3_in[240]),
   .I1(level3_in[241]),
   .I2(level3_in[242]),
   .I3(level3_in[243]),
   .I4(level3_in[244]),
   .I5(level3_in[245])
);

LUT6 #(
   .INIT(64'h2b3e26db2b3e26db)  
) LUT6_inst9113 (
   .O(to_level2[41]),
   .I0(level3_in[246]),
   .I1(level3_in[247]),
   .I2(level3_in[248]),
   .I3(level3_in[249]),
   .I4(level3_in[250]),
   .I5(level3_in[251])
);

LUT6 #(
   .INIT(64'hced64f1fced64f1f)  
) LUT6_inst9114 (
   .O(to_level2[42]),
   .I0(level3_in[252]),
   .I1(level3_in[253]),
   .I2(level3_in[254]),
   .I3(level3_in[255]),
   .I4(level3_in[256]),
   .I5(level3_in[257])
);

LUT6 #(
   .INIT(64'hf7e8bb1ef7e8bb1e)  
) LUT6_inst9115 (
   .O(to_level2[43]),
   .I0(level3_in[258]),
   .I1(level3_in[259]),
   .I2(level3_in[260]),
   .I3(level3_in[261]),
   .I4(level3_in[262]),
   .I5(level3_in[263])
);

LUT6 #(
   .INIT(64'hdcf82f56dcf82f56)  
) LUT6_inst9116 (
   .O(to_level2[44]),
   .I0(level3_in[264]),
   .I1(level3_in[265]),
   .I2(level3_in[266]),
   .I3(level3_in[267]),
   .I4(level3_in[268]),
   .I5(level3_in[269])
);

LUT6 #(
   .INIT(64'h62a6f42862a6f428)  
) LUT6_inst9117 (
   .O(to_level2[45]),
   .I0(level3_in[270]),
   .I1(level3_in[271]),
   .I2(level3_in[272]),
   .I3(level3_in[273]),
   .I4(level3_in[274]),
   .I5(level3_in[275])
);

LUT6 #(
   .INIT(64'h0ce43b140ce43b14)  
) LUT6_inst9118 (
   .O(to_level2[46]),
   .I0(level3_in[276]),
   .I1(level3_in[277]),
   .I2(level3_in[278]),
   .I3(level3_in[279]),
   .I4(level3_in[280]),
   .I5(level3_in[281])
);

LUT6 #(
   .INIT(64'h425dda9b425dda9b)  
) LUT6_inst9119 (
   .O(to_level2[47]),
   .I0(level3_in[282]),
   .I1(level3_in[283]),
   .I2(level3_in[284]),
   .I3(level3_in[285]),
   .I4(level3_in[286]),
   .I5(level3_in[287])
);

LUT6 #(
   .INIT(64'hc26aaf7dc26aaf7d)  
) LUT6_inst9120 (
   .O(to_level2[48]),
   .I0(level3_in[288]),
   .I1(level3_in[289]),
   .I2(level3_in[290]),
   .I3(level3_in[291]),
   .I4(level3_in[292]),
   .I5(level3_in[293])
);

LUT6 #(
   .INIT(64'h434fc830434fc830)  
) LUT6_inst9121 (
   .O(to_level2[49]),
   .I0(level3_in[294]),
   .I1(level3_in[295]),
   .I2(level3_in[296]),
   .I3(level3_in[297]),
   .I4(level3_in[298]),
   .I5(level3_in[299])
);

LUT6 #(
   .INIT(64'h8918458489184584)  
) LUT6_inst9122 (
   .O(to_level2[50]),
   .I0(level3_in[300]),
   .I1(level3_in[301]),
   .I2(level3_in[302]),
   .I3(level3_in[303]),
   .I4(level3_in[304]),
   .I5(level3_in[305])
);

LUT6 #(
   .INIT(64'hf34527b8f34527b8)  
) LUT6_inst9123 (
   .O(to_level2[51]),
   .I0(level3_in[306]),
   .I1(level3_in[307]),
   .I2(level3_in[308]),
   .I3(level3_in[309]),
   .I4(level3_in[310]),
   .I5(level3_in[311])
);

LUT6 #(
   .INIT(64'haccbb387accbb387)  
) LUT6_inst9124 (
   .O(to_level2[52]),
   .I0(level3_in[312]),
   .I1(level3_in[313]),
   .I2(level3_in[314]),
   .I3(level3_in[315]),
   .I4(level3_in[316]),
   .I5(level3_in[317])
);

LUT6 #(
   .INIT(64'h1ed8f7121ed8f712)  
) LUT6_inst9125 (
   .O(to_level2[53]),
   .I0(level3_in[318]),
   .I1(level3_in[319]),
   .I2(level3_in[320]),
   .I3(level3_in[321]),
   .I4(level3_in[322]),
   .I5(level3_in[323])
);

LUT6 #(
   .INIT(64'hbd65a1dbbd65a1db)  
) LUT6_inst9126 (
   .O(to_level2[54]),
   .I0(level3_in[324]),
   .I1(level3_in[325]),
   .I2(level3_in[326]),
   .I3(level3_in[327]),
   .I4(level3_in[328]),
   .I5(level3_in[329])
);

LUT6 #(
   .INIT(64'h872e4887872e4887)  
) LUT6_inst9127 (
   .O(to_level2[55]),
   .I0(level3_in[330]),
   .I1(level3_in[331]),
   .I2(level3_in[332]),
   .I3(level3_in[333]),
   .I4(level3_in[334]),
   .I5(level3_in[335])
);

LUT6 #(
   .INIT(64'h5548976055489760)  
) LUT6_inst9128 (
   .O(to_level2[56]),
   .I0(level3_in[336]),
   .I1(level3_in[337]),
   .I2(level3_in[338]),
   .I3(level3_in[339]),
   .I4(level3_in[340]),
   .I5(level3_in[341])
);

LUT6 #(
   .INIT(64'h707e57c4707e57c4)  
) LUT6_inst9129 (
   .O(to_level2[57]),
   .I0(level3_in[342]),
   .I1(level3_in[343]),
   .I2(level3_in[344]),
   .I3(level3_in[345]),
   .I4(level3_in[346]),
   .I5(level3_in[347])
);

LUT6 #(
   .INIT(64'hd73e546fd73e546f)  
) LUT6_inst9130 (
   .O(to_level2[58]),
   .I0(level3_in[348]),
   .I1(level3_in[349]),
   .I2(level3_in[350]),
   .I3(level3_in[351]),
   .I4(level3_in[352]),
   .I5(level3_in[353])
);

LUT6 #(
   .INIT(64'h87e295f087e295f0)  
) LUT6_inst9131 (
   .O(to_level2[59]),
   .I0(level3_in[354]),
   .I1(level3_in[355]),
   .I2(level3_in[356]),
   .I3(level3_in[357]),
   .I4(level3_in[358]),
   .I5(level3_in[359])
);

LUT6 #(
   .INIT(64'hd18708e3d18708e3)  
) LUT6_inst9132 (
   .O(to_level2[60]),
   .I0(level3_in[360]),
   .I1(level3_in[361]),
   .I2(level3_in[362]),
   .I3(level3_in[363]),
   .I4(level3_in[364]),
   .I5(level3_in[365])
);

LUT6 #(
   .INIT(64'hfdcaa13dfdcaa13d)  
) LUT6_inst9133 (
   .O(to_level2[61]),
   .I0(level3_in[366]),
   .I1(level3_in[367]),
   .I2(level3_in[368]),
   .I3(level3_in[369]),
   .I4(level3_in[370]),
   .I5(level3_in[371])
);

LUT6 #(
   .INIT(64'haf401376af401376)  
) LUT6_inst9134 (
   .O(to_level2[62]),
   .I0(level3_in[372]),
   .I1(level3_in[373]),
   .I2(level3_in[374]),
   .I3(level3_in[375]),
   .I4(level3_in[376]),
   .I5(level3_in[377])
);

LUT6 #(
   .INIT(64'hb2bad5fcb2bad5fc)  
) LUT6_inst9135 (
   .O(to_level2[63]),
   .I0(level3_in[378]),
   .I1(level3_in[379]),
   .I2(level3_in[380]),
   .I3(level3_in[381]),
   .I4(level3_in[382]),
   .I5(level3_in[383])
);

LUT6 #(
   .INIT(64'h4c6e95b44c6e95b4)  
) LUT6_inst9136 (
   .O(to_level2[64]),
   .I0(level3_in[384]),
   .I1(level3_in[385]),
   .I2(level3_in[386]),
   .I3(level3_in[387]),
   .I4(level3_in[388]),
   .I5(level3_in[389])
);

LUT6 #(
   .INIT(64'h7fc10d2b7fc10d2b)  
) LUT6_inst9137 (
   .O(to_level2[65]),
   .I0(level3_in[390]),
   .I1(level3_in[391]),
   .I2(level3_in[392]),
   .I3(level3_in[393]),
   .I4(level3_in[394]),
   .I5(level3_in[395])
);

LUT6 #(
   .INIT(64'hc5d6242dc5d6242d)  
) LUT6_inst9138 (
   .O(to_level2[66]),
   .I0(level3_in[396]),
   .I1(level3_in[397]),
   .I2(level3_in[398]),
   .I3(level3_in[399]),
   .I4(level3_in[400]),
   .I5(level3_in[401])
);

LUT6 #(
   .INIT(64'hf058c03cf058c03c)  
) LUT6_inst9139 (
   .O(to_level2[67]),
   .I0(level3_in[402]),
   .I1(level3_in[403]),
   .I2(level3_in[404]),
   .I3(level3_in[405]),
   .I4(level3_in[406]),
   .I5(level3_in[407])
);

LUT6 #(
   .INIT(64'h0a6c4b790a6c4b79)  
) LUT6_inst9140 (
   .O(to_level2[68]),
   .I0(level3_in[408]),
   .I1(level3_in[409]),
   .I2(level3_in[410]),
   .I3(level3_in[411]),
   .I4(level3_in[412]),
   .I5(level3_in[413])
);

LUT6 #(
   .INIT(64'hfcb58141fcb58141)  
) LUT6_inst9141 (
   .O(to_level2[69]),
   .I0(level3_in[414]),
   .I1(level3_in[415]),
   .I2(level3_in[416]),
   .I3(level3_in[417]),
   .I4(level3_in[418]),
   .I5(level3_in[419])
);

LUT6 #(
   .INIT(64'h22776d9622776d96)  
) LUT6_inst9142 (
   .O(to_level2[70]),
   .I0(level3_in[420]),
   .I1(level3_in[421]),
   .I2(level3_in[422]),
   .I3(level3_in[423]),
   .I4(level3_in[424]),
   .I5(level3_in[425])
);

LUT6 #(
   .INIT(64'h72dc9f5472dc9f54)  
) LUT6_inst9143 (
   .O(to_level2[71]),
   .I0(level3_in[426]),
   .I1(level3_in[427]),
   .I2(level3_in[428]),
   .I3(level3_in[429]),
   .I4(level3_in[430]),
   .I5(level3_in[431])
);

LUT6 #(
   .INIT(64'h885ff8be885ff8be)  
) LUT6_inst9144 (
   .O(to_level2[72]),
   .I0(level3_in[432]),
   .I1(level3_in[433]),
   .I2(level3_in[434]),
   .I3(level3_in[435]),
   .I4(level3_in[436]),
   .I5(level3_in[437])
);

LUT6 #(
   .INIT(64'ha1848744a1848744)  
) LUT6_inst9145 (
   .O(to_level2[73]),
   .I0(level3_in[438]),
   .I1(level3_in[439]),
   .I2(level3_in[440]),
   .I3(level3_in[441]),
   .I4(level3_in[442]),
   .I5(level3_in[443])
);

LUT6 #(
   .INIT(64'he72685a5e72685a5)  
) LUT6_inst9146 (
   .O(to_level2[74]),
   .I0(level3_in[444]),
   .I1(level3_in[445]),
   .I2(level3_in[446]),
   .I3(level3_in[447]),
   .I4(level3_in[448]),
   .I5(level3_in[449])
);

LUT6 #(
   .INIT(64'h42a32a0c42a32a0c)  
) LUT6_inst9147 (
   .O(to_level2[75]),
   .I0(level3_in[450]),
   .I1(level3_in[451]),
   .I2(level3_in[452]),
   .I3(level3_in[453]),
   .I4(level3_in[454]),
   .I5(level3_in[455])
);

LUT6 #(
   .INIT(64'h7d610dd27d610dd2)  
) LUT6_inst9148 (
   .O(to_level2[76]),
   .I0(level3_in[456]),
   .I1(level3_in[457]),
   .I2(level3_in[458]),
   .I3(level3_in[459]),
   .I4(level3_in[460]),
   .I5(level3_in[461])
);

LUT6 #(
   .INIT(64'hb44968afb44968af)  
) LUT6_inst9149 (
   .O(to_level2[77]),
   .I0(level3_in[462]),
   .I1(level3_in[463]),
   .I2(level3_in[464]),
   .I3(level3_in[465]),
   .I4(level3_in[466]),
   .I5(level3_in[467])
);

LUT6 #(
   .INIT(64'h2d63b4462d63b446)  
) LUT6_inst9150 (
   .O(to_level2[78]),
   .I0(level3_in[468]),
   .I1(level3_in[469]),
   .I2(level3_in[470]),
   .I3(level3_in[471]),
   .I4(level3_in[472]),
   .I5(level3_in[473])
);

LUT6 #(
   .INIT(64'he2b70ba1e2b70ba1)  
) LUT6_inst9151 (
   .O(to_level2[79]),
   .I0(level3_in[474]),
   .I1(level3_in[475]),
   .I2(level3_in[476]),
   .I3(level3_in[477]),
   .I4(level3_in[478]),
   .I5(level3_in[479])
);

LUT6 #(
   .INIT(64'h9537871995378719)  
) LUT6_inst9152 (
   .O(to_level2[80]),
   .I0(level3_in[480]),
   .I1(level3_in[481]),
   .I2(level3_in[482]),
   .I3(level3_in[483]),
   .I4(level3_in[484]),
   .I5(level3_in[485])
);

LUT6 #(
   .INIT(64'hb2ab0fd2b2ab0fd2)  
) LUT6_inst9153 (
   .O(to_level2[81]),
   .I0(level3_in[486]),
   .I1(level3_in[487]),
   .I2(level3_in[488]),
   .I3(level3_in[489]),
   .I4(level3_in[490]),
   .I5(level3_in[491])
);

LUT6 #(
   .INIT(64'h48faf14548faf145)  
) LUT6_inst9154 (
   .O(to_level2[82]),
   .I0(level3_in[492]),
   .I1(level3_in[493]),
   .I2(level3_in[494]),
   .I3(level3_in[495]),
   .I4(level3_in[496]),
   .I5(level3_in[497])
);

LUT6 #(
   .INIT(64'hdc4b6ca6dc4b6ca6)  
) LUT6_inst9155 (
   .O(to_level2[83]),
   .I0(level3_in[498]),
   .I1(level3_in[499]),
   .I2(level3_in[500]),
   .I3(level3_in[501]),
   .I4(level3_in[502]),
   .I5(level3_in[503])
);

LUT6 #(
   .INIT(64'hd8c558ddd8c558dd)  
) LUT6_inst9156 (
   .O(to_level2[84]),
   .I0(level3_in[504]),
   .I1(level3_in[505]),
   .I2(level3_in[506]),
   .I3(level3_in[507]),
   .I4(level3_in[508]),
   .I5(level3_in[509])
);

LUT6 #(
   .INIT(64'h239ed421239ed421)  
) LUT6_inst9157 (
   .O(to_level2[85]),
   .I0(level3_in[510]),
   .I1(level3_in[511]),
   .I2(level3_in[512]),
   .I3(level3_in[513]),
   .I4(level3_in[514]),
   .I5(level3_in[515])
);

LUT6 #(
   .INIT(64'he215d537e215d537)  
) LUT6_inst9158 (
   .O(to_level2[86]),
   .I0(level3_in[516]),
   .I1(level3_in[517]),
   .I2(level3_in[518]),
   .I3(level3_in[519]),
   .I4(level3_in[520]),
   .I5(level3_in[521])
);

LUT6 #(
   .INIT(64'hb3242740b3242740)  
) LUT6_inst9159 (
   .O(to_level2[87]),
   .I0(level3_in[522]),
   .I1(level3_in[523]),
   .I2(level3_in[524]),
   .I3(level3_in[525]),
   .I4(level3_in[526]),
   .I5(level3_in[527])
);

LUT6 #(
   .INIT(64'h5599c02a5599c02a)  
) LUT6_inst9160 (
   .O(to_level2[88]),
   .I0(level3_in[528]),
   .I1(level3_in[529]),
   .I2(level3_in[530]),
   .I3(level3_in[531]),
   .I4(level3_in[532]),
   .I5(level3_in[533])
);

LUT6 #(
   .INIT(64'he69323d3e69323d3)  
) LUT6_inst9161 (
   .O(to_level2[89]),
   .I0(level3_in[534]),
   .I1(level3_in[535]),
   .I2(level3_in[536]),
   .I3(level3_in[537]),
   .I4(level3_in[538]),
   .I5(level3_in[539])
);

LUT6 #(
   .INIT(64'h9e6999d29e6999d2)  
) LUT6_inst9162 (
   .O(to_level2[90]),
   .I0(level3_in[540]),
   .I1(level3_in[541]),
   .I2(level3_in[542]),
   .I3(level3_in[543]),
   .I4(level3_in[544]),
   .I5(level3_in[545])
);

LUT6 #(
   .INIT(64'h726fd8c9726fd8c9)  
) LUT6_inst9163 (
   .O(to_level2[91]),
   .I0(level3_in[546]),
   .I1(level3_in[547]),
   .I2(level3_in[548]),
   .I3(level3_in[549]),
   .I4(level3_in[550]),
   .I5(level3_in[551])
);

LUT6 #(
   .INIT(64'h5260e0125260e012)  
) LUT6_inst9164 (
   .O(to_level2[92]),
   .I0(level3_in[552]),
   .I1(level3_in[553]),
   .I2(level3_in[554]),
   .I3(level3_in[555]),
   .I4(level3_in[556]),
   .I5(level3_in[557])
);

LUT6 #(
   .INIT(64'hd155b617d155b617)  
) LUT6_inst9165 (
   .O(to_level2[93]),
   .I0(level3_in[558]),
   .I1(level3_in[559]),
   .I2(level3_in[560]),
   .I3(level3_in[561]),
   .I4(level3_in[562]),
   .I5(level3_in[563])
);

LUT6 #(
   .INIT(64'h3807058438070584)  
) LUT6_inst9166 (
   .O(to_level2[94]),
   .I0(level3_in[564]),
   .I1(level3_in[565]),
   .I2(level3_in[566]),
   .I3(level3_in[567]),
   .I4(level3_in[568]),
   .I5(level3_in[569])
);

LUT6 #(
   .INIT(64'h0d7699220d769922)  
) LUT6_inst9167 (
   .O(to_level2[95]),
   .I0(level3_in[570]),
   .I1(level3_in[571]),
   .I2(level3_in[572]),
   .I3(level3_in[573]),
   .I4(level3_in[574]),
   .I5(level3_in[575])
);

LUT6 #(
   .INIT(64'h40817a9b40817a9b)  
) LUT6_inst9168 (
   .O(to_level2[96]),
   .I0(level3_in[576]),
   .I1(level3_in[577]),
   .I2(level3_in[578]),
   .I3(level3_in[579]),
   .I4(level3_in[580]),
   .I5(level3_in[581])
);

LUT6 #(
   .INIT(64'h063f0bec063f0bec)  
) LUT6_inst9169 (
   .O(to_level2[97]),
   .I0(level3_in[582]),
   .I1(level3_in[583]),
   .I2(level3_in[584]),
   .I3(level3_in[585]),
   .I4(level3_in[586]),
   .I5(level3_in[587])
);

LUT6 #(
   .INIT(64'hc44fb4cbc44fb4cb)  
) LUT6_inst9170 (
   .O(to_level2[98]),
   .I0(level3_in[588]),
   .I1(level3_in[589]),
   .I2(level3_in[590]),
   .I3(level3_in[591]),
   .I4(level3_in[592]),
   .I5(level3_in[593])
);

LUT6 #(
   .INIT(64'h9163478d9163478d)  
) LUT6_inst9171 (
   .O(to_level2[99]),
   .I0(level3_in[594]),
   .I1(level3_in[595]),
   .I2(level3_in[596]),
   .I3(level3_in[597]),
   .I4(level3_in[598]),
   .I5(level3_in[599])
);

LUT6 #(
   .INIT(64'hb891d091b891d091)  
) LUT6_inst9172 (
   .O(to_level2[100]),
   .I0(level3_in[600]),
   .I1(level3_in[601]),
   .I2(level3_in[602]),
   .I3(level3_in[603]),
   .I4(level3_in[604]),
   .I5(level3_in[605])
);

LUT6 #(
   .INIT(64'hbdb66c3abdb66c3a)  
) LUT6_inst9173 (
   .O(to_level2[101]),
   .I0(level3_in[606]),
   .I1(level3_in[607]),
   .I2(level3_in[608]),
   .I3(level3_in[609]),
   .I4(level3_in[610]),
   .I5(level3_in[611])
);

LUT6 #(
   .INIT(64'h7f1be0de7f1be0de)  
) LUT6_inst9174 (
   .O(to_level2[102]),
   .I0(level3_in[612]),
   .I1(level3_in[613]),
   .I2(level3_in[614]),
   .I3(level3_in[615]),
   .I4(level3_in[616]),
   .I5(level3_in[617])
);

LUT6 #(
   .INIT(64'h82786ec282786ec2)  
) LUT6_inst9175 (
   .O(to_level2[103]),
   .I0(level3_in[618]),
   .I1(level3_in[619]),
   .I2(level3_in[620]),
   .I3(level3_in[621]),
   .I4(level3_in[622]),
   .I5(level3_in[623])
);

LUT6 #(
   .INIT(64'h6bb104b26bb104b2)  
) LUT6_inst9176 (
   .O(to_level2[104]),
   .I0(level3_in[624]),
   .I1(level3_in[625]),
   .I2(level3_in[626]),
   .I3(level3_in[627]),
   .I4(level3_in[628]),
   .I5(level3_in[629])
);

LUT6 #(
   .INIT(64'h57ed77fa57ed77fa)  
) LUT6_inst9177 (
   .O(to_level2[105]),
   .I0(level3_in[630]),
   .I1(level3_in[631]),
   .I2(level3_in[632]),
   .I3(level3_in[633]),
   .I4(level3_in[634]),
   .I5(level3_in[635])
);

LUT6 #(
   .INIT(64'h8ec274f58ec274f5)  
) LUT6_inst9178 (
   .O(to_level2[106]),
   .I0(level3_in[636]),
   .I1(level3_in[637]),
   .I2(level3_in[638]),
   .I3(level3_in[639]),
   .I4(level3_in[640]),
   .I5(level3_in[641])
);

LUT6 #(
   .INIT(64'h2e670bbf2e670bbf)  
) LUT6_inst9179 (
   .O(to_level2[107]),
   .I0(level3_in[642]),
   .I1(level3_in[643]),
   .I2(level3_in[644]),
   .I3(level3_in[645]),
   .I4(level3_in[646]),
   .I5(level3_in[647])
);

LUT6 #(
   .INIT(64'h3140b9c23140b9c2)  
) LUT6_inst9180 (
   .O(to_level2[108]),
   .I0(level3_in[648]),
   .I1(level3_in[649]),
   .I2(level3_in[650]),
   .I3(level3_in[651]),
   .I4(level3_in[652]),
   .I5(level3_in[653])
);

LUT6 #(
   .INIT(64'h6e42d9fb6e42d9fb)  
) LUT6_inst9181 (
   .O(to_level2[109]),
   .I0(level3_in[654]),
   .I1(level3_in[655]),
   .I2(level3_in[656]),
   .I3(level3_in[657]),
   .I4(level3_in[658]),
   .I5(level3_in[659])
);

LUT6 #(
   .INIT(64'h7fe9da3f7fe9da3f)  
) LUT6_inst9182 (
   .O(to_level2[110]),
   .I0(level3_in[660]),
   .I1(level3_in[661]),
   .I2(level3_in[662]),
   .I3(level3_in[663]),
   .I4(level3_in[664]),
   .I5(level3_in[665])
);

LUT6 #(
   .INIT(64'h3b5c1b053b5c1b05)  
) LUT6_inst9183 (
   .O(to_level2[111]),
   .I0(level3_in[666]),
   .I1(level3_in[667]),
   .I2(level3_in[668]),
   .I3(level3_in[669]),
   .I4(level3_in[670]),
   .I5(level3_in[671])
);

LUT6 #(
   .INIT(64'h1e2643491e264349)  
) LUT6_inst9184 (
   .O(to_level2[112]),
   .I0(level3_in[672]),
   .I1(level3_in[673]),
   .I2(level3_in[674]),
   .I3(level3_in[675]),
   .I4(level3_in[676]),
   .I5(level3_in[677])
);

LUT6 #(
   .INIT(64'ha4a19fc1a4a19fc1)  
) LUT6_inst9185 (
   .O(to_level2[113]),
   .I0(level3_in[678]),
   .I1(level3_in[679]),
   .I2(level3_in[680]),
   .I3(level3_in[681]),
   .I4(level3_in[682]),
   .I5(level3_in[683])
);

LUT6 #(
   .INIT(64'hd99030bed99030be)  
) LUT6_inst9186 (
   .O(to_level2[114]),
   .I0(level3_in[684]),
   .I1(level3_in[685]),
   .I2(level3_in[686]),
   .I3(level3_in[687]),
   .I4(level3_in[688]),
   .I5(level3_in[689])
);

LUT6 #(
   .INIT(64'h88e1ee6888e1ee68)  
) LUT6_inst9187 (
   .O(to_level2[115]),
   .I0(level3_in[690]),
   .I1(level3_in[691]),
   .I2(level3_in[692]),
   .I3(level3_in[693]),
   .I4(level3_in[694]),
   .I5(level3_in[695])
);

LUT6 #(
   .INIT(64'h6bbca7a56bbca7a5)  
) LUT6_inst9188 (
   .O(to_level2[116]),
   .I0(level3_in[696]),
   .I1(level3_in[697]),
   .I2(level3_in[698]),
   .I3(level3_in[699]),
   .I4(level3_in[700]),
   .I5(level3_in[701])
);

LUT6 #(
   .INIT(64'hd3517803d3517803)  
) LUT6_inst9189 (
   .O(to_level2[117]),
   .I0(level3_in[702]),
   .I1(level3_in[703]),
   .I2(level3_in[704]),
   .I3(level3_in[705]),
   .I4(level3_in[706]),
   .I5(level3_in[707])
);

LUT6 #(
   .INIT(64'h8a4471598a447159)  
) LUT6_inst9190 (
   .O(to_level2[118]),
   .I0(level3_in[708]),
   .I1(level3_in[709]),
   .I2(level3_in[710]),
   .I3(level3_in[711]),
   .I4(level3_in[712]),
   .I5(level3_in[713])
);

LUT6 #(
   .INIT(64'heafdb063eafdb063)  
) LUT6_inst9191 (
   .O(to_level2[119]),
   .I0(level3_in[714]),
   .I1(level3_in[715]),
   .I2(level3_in[716]),
   .I3(level3_in[717]),
   .I4(level3_in[718]),
   .I5(level3_in[719])
);

LUT6 #(
   .INIT(64'h6c8398656c839865)  
) LUT6_inst9192 (
   .O(to_level2[120]),
   .I0(level3_in[720]),
   .I1(level3_in[721]),
   .I2(level3_in[722]),
   .I3(level3_in[723]),
   .I4(level3_in[724]),
   .I5(level3_in[725])
);

LUT6 #(
   .INIT(64'h2fd7023e2fd7023e)  
) LUT6_inst9193 (
   .O(to_level2[121]),
   .I0(level3_in[726]),
   .I1(level3_in[727]),
   .I2(level3_in[728]),
   .I3(level3_in[729]),
   .I4(level3_in[730]),
   .I5(level3_in[731])
);

LUT6 #(
   .INIT(64'h69fe0b0c69fe0b0c)  
) LUT6_inst9194 (
   .O(to_level2[122]),
   .I0(level3_in[732]),
   .I1(level3_in[733]),
   .I2(level3_in[734]),
   .I3(level3_in[735]),
   .I4(level3_in[736]),
   .I5(level3_in[737])
);

LUT6 #(
   .INIT(64'h82f0215582f02155)  
) LUT6_inst9195 (
   .O(to_level2[123]),
   .I0(level3_in[738]),
   .I1(level3_in[739]),
   .I2(level3_in[740]),
   .I3(level3_in[741]),
   .I4(level3_in[742]),
   .I5(level3_in[743])
);

LUT6 #(
   .INIT(64'h9ccc4cd19ccc4cd1)  
) LUT6_inst9196 (
   .O(to_level2[124]),
   .I0(level3_in[744]),
   .I1(level3_in[745]),
   .I2(level3_in[746]),
   .I3(level3_in[747]),
   .I4(level3_in[748]),
   .I5(level3_in[749])
);

LUT6 #(
   .INIT(64'h94633dc394633dc3)  
) LUT6_inst9197 (
   .O(to_level2[125]),
   .I0(level3_in[750]),
   .I1(level3_in[751]),
   .I2(level3_in[752]),
   .I3(level3_in[753]),
   .I4(level3_in[754]),
   .I5(level3_in[755])
);

LUT6 #(
   .INIT(64'h86d4196686d41966)  
) LUT6_inst9198 (
   .O(to_level2[126]),
   .I0(level3_in[756]),
   .I1(level3_in[757]),
   .I2(level3_in[758]),
   .I3(level3_in[759]),
   .I4(level3_in[760]),
   .I5(level3_in[761])
);

LUT6 #(
   .INIT(64'ha79cc0b1a79cc0b1)  
) LUT6_inst9199 (
   .O(to_level2[127]),
   .I0(level3_in[762]),
   .I1(level3_in[763]),
   .I2(level3_in[764]),
   .I3(level3_in[765]),
   .I4(level3_in[766]),
   .I5(level3_in[767])
);

LUT6 #(
   .INIT(64'hafe3c802afe3c802)  
) LUT6_inst9200 (
   .O(to_level2[128]),
   .I0(level3_in[768]),
   .I1(level3_in[769]),
   .I2(level3_in[770]),
   .I3(level3_in[771]),
   .I4(level3_in[772]),
   .I5(level3_in[773])
);

LUT6 #(
   .INIT(64'ha553f8f7a553f8f7)  
) LUT6_inst9201 (
   .O(to_level2[129]),
   .I0(level3_in[774]),
   .I1(level3_in[775]),
   .I2(level3_in[776]),
   .I3(level3_in[777]),
   .I4(level3_in[778]),
   .I5(level3_in[779])
);

LUT6 #(
   .INIT(64'h39986b2d39986b2d)  
) LUT6_inst9202 (
   .O(to_level2[130]),
   .I0(level3_in[780]),
   .I1(level3_in[781]),
   .I2(level3_in[782]),
   .I3(level3_in[783]),
   .I4(level3_in[784]),
   .I5(level3_in[785])
);

LUT6 #(
   .INIT(64'h9a1aaece9a1aaece)  
) LUT6_inst9203 (
   .O(to_level2[131]),
   .I0(level3_in[786]),
   .I1(level3_in[787]),
   .I2(level3_in[788]),
   .I3(level3_in[789]),
   .I4(level3_in[790]),
   .I5(level3_in[791])
);

LUT6 #(
   .INIT(64'h72c0b23872c0b238)  
) LUT6_inst9204 (
   .O(to_level2[132]),
   .I0(level3_in[792]),
   .I1(level3_in[793]),
   .I2(level3_in[794]),
   .I3(level3_in[795]),
   .I4(level3_in[796]),
   .I5(level3_in[797])
);

LUT6 #(
   .INIT(64'hafb18403afb18403)  
) LUT6_inst9205 (
   .O(to_level2[133]),
   .I0(level3_in[798]),
   .I1(level3_in[799]),
   .I2(level3_in[800]),
   .I3(level3_in[801]),
   .I4(level3_in[802]),
   .I5(level3_in[803])
);

LUT6 #(
   .INIT(64'hc46b6fe8c46b6fe8)  
) LUT6_inst9206 (
   .O(to_level2[134]),
   .I0(level3_in[804]),
   .I1(level3_in[805]),
   .I2(level3_in[806]),
   .I3(level3_in[807]),
   .I4(level3_in[808]),
   .I5(level3_in[809])
);

LUT6 #(
   .INIT(64'h13f46b9913f46b99)  
) LUT6_inst9207 (
   .O(to_level2[135]),
   .I0(level3_in[810]),
   .I1(level3_in[811]),
   .I2(level3_in[812]),
   .I3(level3_in[813]),
   .I4(level3_in[814]),
   .I5(level3_in[815])
);

LUT6 #(
   .INIT(64'head94244ead94244)  
) LUT6_inst9208 (
   .O(to_level2[136]),
   .I0(level3_in[816]),
   .I1(level3_in[817]),
   .I2(level3_in[818]),
   .I3(level3_in[819]),
   .I4(level3_in[820]),
   .I5(level3_in[821])
);

LUT6 #(
   .INIT(64'h67a3111767a31117)  
) LUT6_inst9209 (
   .O(to_level2[137]),
   .I0(level3_in[822]),
   .I1(level3_in[823]),
   .I2(level3_in[824]),
   .I3(level3_in[825]),
   .I4(level3_in[826]),
   .I5(level3_in[827])
);

LUT6 #(
   .INIT(64'hdfc63307dfc63307)  
) LUT6_inst9210 (
   .O(to_level2[138]),
   .I0(level3_in[828]),
   .I1(level3_in[829]),
   .I2(level3_in[830]),
   .I3(level3_in[831]),
   .I4(level3_in[832]),
   .I5(level3_in[833])
);

LUT6 #(
   .INIT(64'hb54e9742b54e9742)  
) LUT6_inst9211 (
   .O(to_level2[139]),
   .I0(level3_in[834]),
   .I1(level3_in[835]),
   .I2(level3_in[836]),
   .I3(level3_in[837]),
   .I4(level3_in[838]),
   .I5(level3_in[839])
);

LUT6 #(
   .INIT(64'h24af7e4f24af7e4f)  
) LUT6_inst9212 (
   .O(to_level2[140]),
   .I0(level3_in[840]),
   .I1(level3_in[841]),
   .I2(level3_in[842]),
   .I3(level3_in[843]),
   .I4(level3_in[844]),
   .I5(level3_in[845])
);

LUT6 #(
   .INIT(64'h9cdc50169cdc5016)  
) LUT6_inst9213 (
   .O(to_level2[141]),
   .I0(level3_in[846]),
   .I1(level3_in[847]),
   .I2(level3_in[848]),
   .I3(level3_in[849]),
   .I4(level3_in[850]),
   .I5(level3_in[851])
);

LUT6 #(
   .INIT(64'h1c92a70a1c92a70a)  
) LUT6_inst9214 (
   .O(to_level2[142]),
   .I0(level3_in[852]),
   .I1(level3_in[853]),
   .I2(level3_in[854]),
   .I3(level3_in[855]),
   .I4(level3_in[856]),
   .I5(level3_in[857])
);

LUT6 #(
   .INIT(64'h597825de597825de)  
) LUT6_inst9215 (
   .O(to_level2[143]),
   .I0(level3_in[858]),
   .I1(level3_in[859]),
   .I2(level3_in[860]),
   .I3(level3_in[861]),
   .I4(level3_in[862]),
   .I5(level3_in[863])
);

LUT6 #(
   .INIT(64'h8661edf68661edf6)  
) LUT6_inst9216 (
   .O(to_level2[144]),
   .I0(level3_in[864]),
   .I1(level3_in[865]),
   .I2(level3_in[866]),
   .I3(level3_in[867]),
   .I4(level3_in[868]),
   .I5(level3_in[869])
);

LUT6 #(
   .INIT(64'h228a9315228a9315)  
) LUT6_inst9217 (
   .O(to_level2[145]),
   .I0(level3_in[870]),
   .I1(level3_in[871]),
   .I2(level3_in[872]),
   .I3(level3_in[873]),
   .I4(level3_in[874]),
   .I5(level3_in[875])
);

LUT6 #(
   .INIT(64'h66231b0766231b07)  
) LUT6_inst9218 (
   .O(to_level2[146]),
   .I0(level3_in[876]),
   .I1(level3_in[877]),
   .I2(level3_in[878]),
   .I3(level3_in[879]),
   .I4(level3_in[880]),
   .I5(level3_in[881])
);

LUT6 #(
   .INIT(64'h1121d6181121d618)  
) LUT6_inst9219 (
   .O(to_level2[147]),
   .I0(level3_in[882]),
   .I1(level3_in[883]),
   .I2(level3_in[884]),
   .I3(level3_in[885]),
   .I4(level3_in[886]),
   .I5(level3_in[887])
);

LUT6 #(
   .INIT(64'h7fa9c8197fa9c819)  
) LUT6_inst9220 (
   .O(to_level2[148]),
   .I0(level3_in[888]),
   .I1(level3_in[889]),
   .I2(level3_in[890]),
   .I3(level3_in[891]),
   .I4(level3_in[892]),
   .I5(level3_in[893])
);

LUT6 #(
   .INIT(64'h591afdc2591afdc2)  
) LUT6_inst9221 (
   .O(to_level2[149]),
   .I0(level3_in[894]),
   .I1(level3_in[895]),
   .I2(level3_in[896]),
   .I3(level3_in[897]),
   .I4(level3_in[898]),
   .I5(level3_in[899])
);

LUT6 #(
   .INIT(64'hde3b9f5bde3b9f5b)  
) LUT6_inst9222 (
   .O(to_level2[150]),
   .I0(level3_in[900]),
   .I1(level3_in[901]),
   .I2(level3_in[902]),
   .I3(level3_in[903]),
   .I4(level3_in[904]),
   .I5(level3_in[905])
);

LUT6 #(
   .INIT(64'h28b20cec28b20cec)  
) LUT6_inst9223 (
   .O(to_level2[151]),
   .I0(level3_in[906]),
   .I1(level3_in[907]),
   .I2(level3_in[908]),
   .I3(level3_in[909]),
   .I4(level3_in[910]),
   .I5(level3_in[911])
);

LUT6 #(
   .INIT(64'h955f075d955f075d)  
) LUT6_inst9224 (
   .O(to_level2[152]),
   .I0(level3_in[912]),
   .I1(level3_in[913]),
   .I2(level3_in[914]),
   .I3(level3_in[915]),
   .I4(level3_in[916]),
   .I5(level3_in[917])
);

LUT6 #(
   .INIT(64'h4875200d4875200d)  
) LUT6_inst9225 (
   .O(to_level2[153]),
   .I0(level3_in[918]),
   .I1(level3_in[919]),
   .I2(level3_in[920]),
   .I3(level3_in[921]),
   .I4(level3_in[922]),
   .I5(level3_in[923])
);

LUT6 #(
   .INIT(64'h72f6e30572f6e305)  
) LUT6_inst9226 (
   .O(to_level2[154]),
   .I0(level3_in[924]),
   .I1(level3_in[925]),
   .I2(level3_in[926]),
   .I3(level3_in[927]),
   .I4(level3_in[928]),
   .I5(level3_in[929])
);

LUT6 #(
   .INIT(64'hc2b2bbedc2b2bbed)  
) LUT6_inst9227 (
   .O(to_level2[155]),
   .I0(level3_in[930]),
   .I1(level3_in[931]),
   .I2(level3_in[932]),
   .I3(level3_in[933]),
   .I4(level3_in[934]),
   .I5(level3_in[935])
);

LUT6 #(
   .INIT(64'h99b5343c99b5343c)  
) LUT6_inst9228 (
   .O(to_level2[156]),
   .I0(level3_in[936]),
   .I1(level3_in[937]),
   .I2(level3_in[938]),
   .I3(level3_in[939]),
   .I4(level3_in[940]),
   .I5(level3_in[941])
);

LUT6 #(
   .INIT(64'h7f0e6f7b7f0e6f7b)  
) LUT6_inst9229 (
   .O(to_level2[157]),
   .I0(level3_in[942]),
   .I1(level3_in[943]),
   .I2(level3_in[944]),
   .I3(level3_in[945]),
   .I4(level3_in[946]),
   .I5(level3_in[947])
);

LUT6 #(
   .INIT(64'hc3ef7a18c3ef7a18)  
) LUT6_inst9230 (
   .O(to_level2[158]),
   .I0(level3_in[948]),
   .I1(level3_in[949]),
   .I2(level3_in[950]),
   .I3(level3_in[951]),
   .I4(level3_in[952]),
   .I5(level3_in[953])
);

LUT6 #(
   .INIT(64'h9a2486c49a2486c4)  
) LUT6_inst9231 (
   .O(to_level2[159]),
   .I0(level3_in[954]),
   .I1(level3_in[955]),
   .I2(level3_in[956]),
   .I3(level3_in[957]),
   .I4(level3_in[958]),
   .I5(level3_in[959])
);

LUT6 #(
   .INIT(64'h729d9814729d9814)  
) LUT6_inst9232 (
   .O(to_level2[160]),
   .I0(level3_in[960]),
   .I1(level3_in[961]),
   .I2(level3_in[962]),
   .I3(level3_in[963]),
   .I4(level3_in[964]),
   .I5(level3_in[965])
);

LUT6 #(
   .INIT(64'h6568ee846568ee84)  
) LUT6_inst9233 (
   .O(to_level2[161]),
   .I0(level3_in[966]),
   .I1(level3_in[967]),
   .I2(level3_in[968]),
   .I3(level3_in[969]),
   .I4(level3_in[970]),
   .I5(level3_in[971])
);

LUT6 #(
   .INIT(64'h2ffc347d2ffc347d)  
) LUT6_inst9234 (
   .O(to_level2[162]),
   .I0(level3_in[972]),
   .I1(level3_in[973]),
   .I2(level3_in[974]),
   .I3(level3_in[975]),
   .I4(level3_in[976]),
   .I5(level3_in[977])
);

LUT6 #(
   .INIT(64'h2578f1fb2578f1fb)  
) LUT6_inst9235 (
   .O(to_level2[163]),
   .I0(level3_in[978]),
   .I1(level3_in[979]),
   .I2(level3_in[980]),
   .I3(level3_in[981]),
   .I4(level3_in[982]),
   .I5(level3_in[983])
);

LUT6 #(
   .INIT(64'h3213ed783213ed78)  
) LUT6_inst9236 (
   .O(to_level2[164]),
   .I0(level3_in[984]),
   .I1(level3_in[985]),
   .I2(level3_in[986]),
   .I3(level3_in[987]),
   .I4(level3_in[988]),
   .I5(level3_in[989])
);

LUT6 #(
   .INIT(64'hfbc021d7fbc021d7)  
) LUT6_inst9237 (
   .O(to_level2[165]),
   .I0(level3_in[990]),
   .I1(level3_in[991]),
   .I2(level3_in[992]),
   .I3(level3_in[993]),
   .I4(level3_in[994]),
   .I5(level3_in[995])
);

LUT6 #(
   .INIT(64'h4b70f5d14b70f5d1)  
) LUT6_inst9238 (
   .O(to_level2[166]),
   .I0(level3_in[996]),
   .I1(level3_in[997]),
   .I2(level3_in[998]),
   .I3(level3_in[999]),
   .I4(level3_in[1000]),
   .I5(level3_in[1001])
);

LUT6 #(
   .INIT(64'h4089d1d24089d1d2)  
) LUT6_inst9239 (
   .O(to_level2[167]),
   .I0(level3_in[1002]),
   .I1(level3_in[1003]),
   .I2(level3_in[1004]),
   .I3(level3_in[1005]),
   .I4(level3_in[1006]),
   .I5(level3_in[1007])
);

LUT6 #(
   .INIT(64'h10d0cd9f10d0cd9f)  
) LUT6_inst9240 (
   .O(to_level2[168]),
   .I0(level3_in[1008]),
   .I1(level3_in[1009]),
   .I2(level3_in[1010]),
   .I3(level3_in[1011]),
   .I4(level3_in[1012]),
   .I5(level3_in[1013])
);

LUT6 #(
   .INIT(64'hebb08da7ebb08da7)  
) LUT6_inst9241 (
   .O(to_level2[169]),
   .I0(level3_in[1014]),
   .I1(level3_in[1015]),
   .I2(level3_in[1016]),
   .I3(level3_in[1017]),
   .I4(level3_in[1018]),
   .I5(level3_in[1019])
);

LUT6 #(
   .INIT(64'hf34aff15f34aff15)  
) LUT6_inst9242 (
   .O(to_level2[170]),
   .I0(level3_in[1020]),
   .I1(level3_in[1021]),
   .I2(level3_in[1022]),
   .I3(level3_in[1023]),
   .I4(level3_in[1024]),
   .I5(level3_in[1025])
);

LUT6 #(
   .INIT(64'hf071eadef071eade)  
) LUT6_inst9243 (
   .O(to_level2[171]),
   .I0(level3_in[1026]),
   .I1(level3_in[1027]),
   .I2(level3_in[1028]),
   .I3(level3_in[1029]),
   .I4(level3_in[1030]),
   .I5(level3_in[1031])
);

LUT6 #(
   .INIT(64'h8eb964858eb96485)  
) LUT6_inst9244 (
   .O(to_level2[172]),
   .I0(level3_in[1032]),
   .I1(level3_in[1033]),
   .I2(level3_in[1034]),
   .I3(level3_in[1035]),
   .I4(level3_in[1036]),
   .I5(level3_in[1037])
);

LUT6 #(
   .INIT(64'h561ff849561ff849)  
) LUT6_inst9245 (
   .O(to_level2[173]),
   .I0(level3_in[1038]),
   .I1(level3_in[1039]),
   .I2(level3_in[1040]),
   .I3(level3_in[1041]),
   .I4(level3_in[1042]),
   .I5(level3_in[1043])
);

LUT6 #(
   .INIT(64'h2d8755b02d8755b0)  
) LUT6_inst9246 (
   .O(to_level2[174]),
   .I0(level3_in[1044]),
   .I1(level3_in[1045]),
   .I2(level3_in[1046]),
   .I3(level3_in[1047]),
   .I4(level3_in[1048]),
   .I5(level3_in[1049])
);

LUT6 #(
   .INIT(64'h6403622964036229)  
) LUT6_inst9247 (
   .O(to_level2[175]),
   .I0(level3_in[1050]),
   .I1(level3_in[1051]),
   .I2(level3_in[1052]),
   .I3(level3_in[1053]),
   .I4(level3_in[1054]),
   .I5(level3_in[1055])
);

LUT6 #(
   .INIT(64'h07129e7b07129e7b)  
) LUT6_inst9248 (
   .O(to_level2[176]),
   .I0(level3_in[1056]),
   .I1(level3_in[1057]),
   .I2(level3_in[1058]),
   .I3(level3_in[1059]),
   .I4(level3_in[1060]),
   .I5(level3_in[1061])
);

LUT6 #(
   .INIT(64'h774136ea774136ea)  
) LUT6_inst9249 (
   .O(to_level2[177]),
   .I0(level3_in[1062]),
   .I1(level3_in[1063]),
   .I2(level3_in[1064]),
   .I3(level3_in[1065]),
   .I4(level3_in[1066]),
   .I5(level3_in[1067])
);

LUT6 #(
   .INIT(64'h08cebc5c08cebc5c)  
) LUT6_inst9250 (
   .O(to_level2[178]),
   .I0(level3_in[1068]),
   .I1(level3_in[1069]),
   .I2(level3_in[1070]),
   .I3(level3_in[1071]),
   .I4(level3_in[1072]),
   .I5(level3_in[1073])
);

LUT6 #(
   .INIT(64'hc1435edfc1435edf)  
) LUT6_inst9251 (
   .O(to_level2[179]),
   .I0(level3_in[1074]),
   .I1(level3_in[1075]),
   .I2(level3_in[1076]),
   .I3(level3_in[1077]),
   .I4(level3_in[1078]),
   .I5(level3_in[1079])
);

LUT6 #(
   .INIT(64'h4cd8e6444cd8e644)  
) LUT6_inst9252 (
   .O(to_level2[180]),
   .I0(level3_in[1080]),
   .I1(level3_in[1081]),
   .I2(level3_in[1082]),
   .I3(level3_in[1083]),
   .I4(level3_in[1084]),
   .I5(level3_in[1085])
);

LUT6 #(
   .INIT(64'haf156da9af156da9)  
) LUT6_inst9253 (
   .O(to_level2[181]),
   .I0(level3_in[1086]),
   .I1(level3_in[1087]),
   .I2(level3_in[1088]),
   .I3(level3_in[1089]),
   .I4(level3_in[1090]),
   .I5(level3_in[1091])
);

LUT6 #(
   .INIT(64'hdaf55758daf55758)  
) LUT6_inst9254 (
   .O(to_level2[182]),
   .I0(level3_in[1092]),
   .I1(level3_in[1093]),
   .I2(level3_in[1094]),
   .I3(level3_in[1095]),
   .I4(level3_in[1096]),
   .I5(level3_in[1097])
);

LUT6 #(
   .INIT(64'h969d46f3969d46f3)  
) LUT6_inst9255 (
   .O(to_level2[183]),
   .I0(level3_in[1098]),
   .I1(level3_in[1099]),
   .I2(level3_in[1100]),
   .I3(level3_in[1101]),
   .I4(level3_in[1102]),
   .I5(level3_in[1103])
);

LUT6 #(
   .INIT(64'h1a1769fa1a1769fa)  
) LUT6_inst9256 (
   .O(to_level2[184]),
   .I0(level3_in[1104]),
   .I1(level3_in[1105]),
   .I2(level3_in[1106]),
   .I3(level3_in[1107]),
   .I4(level3_in[1108]),
   .I5(level3_in[1109])
);

LUT6 #(
   .INIT(64'h6a97a66b6a97a66b)  
) LUT6_inst9257 (
   .O(to_level2[185]),
   .I0(level3_in[1110]),
   .I1(level3_in[1111]),
   .I2(level3_in[1112]),
   .I3(level3_in[1113]),
   .I4(level3_in[1114]),
   .I5(level3_in[1115])
);

LUT6 #(
   .INIT(64'hf38d5c27f38d5c27)  
) LUT6_inst9258 (
   .O(to_level2[186]),
   .I0(level3_in[1116]),
   .I1(level3_in[1117]),
   .I2(level3_in[1118]),
   .I3(level3_in[1119]),
   .I4(level3_in[1120]),
   .I5(level3_in[1121])
);

LUT6 #(
   .INIT(64'h6bdd809c6bdd809c)  
) LUT6_inst9259 (
   .O(to_level2[187]),
   .I0(level3_in[1122]),
   .I1(level3_in[1123]),
   .I2(level3_in[1124]),
   .I3(level3_in[1125]),
   .I4(level3_in[1126]),
   .I5(level3_in[1127])
);

LUT6 #(
   .INIT(64'h9366e45c9366e45c)  
) LUT6_inst9260 (
   .O(to_level2[188]),
   .I0(level3_in[1128]),
   .I1(level3_in[1129]),
   .I2(level3_in[1130]),
   .I3(level3_in[1131]),
   .I4(level3_in[1132]),
   .I5(level3_in[1133])
);

LUT6 #(
   .INIT(64'h6c6167386c616738)  
) LUT6_inst9261 (
   .O(to_level2[189]),
   .I0(level3_in[1134]),
   .I1(level3_in[1135]),
   .I2(level3_in[1136]),
   .I3(level3_in[1137]),
   .I4(level3_in[1138]),
   .I5(level3_in[1139])
);

LUT6 #(
   .INIT(64'hfa4430e2fa4430e2)  
) LUT6_inst9262 (
   .O(to_level2[190]),
   .I0(level3_in[1140]),
   .I1(level3_in[1141]),
   .I2(level3_in[1142]),
   .I3(level3_in[1143]),
   .I4(level3_in[1144]),
   .I5(level3_in[1145])
);

LUT6 #(
   .INIT(64'hff590464ff590464)  
) LUT6_inst9263 (
   .O(to_level2[191]),
   .I0(level3_in[1146]),
   .I1(level3_in[1147]),
   .I2(level3_in[1148]),
   .I3(level3_in[1149]),
   .I4(level3_in[1150]),
   .I5(level3_in[1151])
);

LUT6 #(
   .INIT(64'hd4cbf4fad4cbf4fa)  
) LUT6_inst9264 (
   .O(to_level2[192]),
   .I0(level3_in[1152]),
   .I1(level3_in[1153]),
   .I2(level3_in[1154]),
   .I3(level3_in[1155]),
   .I4(level3_in[1156]),
   .I5(level3_in[1157])
);

LUT6 #(
   .INIT(64'h8078f7bf8078f7bf)  
) LUT6_inst9265 (
   .O(to_level2[193]),
   .I0(level3_in[1158]),
   .I1(level3_in[1159]),
   .I2(level3_in[1160]),
   .I3(level3_in[1161]),
   .I4(level3_in[1162]),
   .I5(level3_in[1163])
);

LUT6 #(
   .INIT(64'hb06468c5b06468c5)  
) LUT6_inst9266 (
   .O(to_level2[194]),
   .I0(level3_in[1164]),
   .I1(level3_in[1165]),
   .I2(level3_in[1166]),
   .I3(level3_in[1167]),
   .I4(level3_in[1168]),
   .I5(level3_in[1169])
);

LUT6 #(
   .INIT(64'h4cc55a4c4cc55a4c)  
) LUT6_inst9267 (
   .O(to_level2[195]),
   .I0(level3_in[1170]),
   .I1(level3_in[1171]),
   .I2(level3_in[1172]),
   .I3(level3_in[1173]),
   .I4(level3_in[1174]),
   .I5(level3_in[1175])
);

LUT6 #(
   .INIT(64'h30a4a99c30a4a99c)  
) LUT6_inst9268 (
   .O(to_level2[196]),
   .I0(level3_in[1176]),
   .I1(level3_in[1177]),
   .I2(level3_in[1178]),
   .I3(level3_in[1179]),
   .I4(level3_in[1180]),
   .I5(level3_in[1181])
);

LUT6 #(
   .INIT(64'had2c4fb0ad2c4fb0)  
) LUT6_inst9269 (
   .O(to_level2[197]),
   .I0(level3_in[1182]),
   .I1(level3_in[1183]),
   .I2(level3_in[1184]),
   .I3(level3_in[1185]),
   .I4(level3_in[1186]),
   .I5(level3_in[1187])
);

LUT6 #(
   .INIT(64'h1e75bbe01e75bbe0)  
) LUT6_inst9270 (
   .O(to_level2[198]),
   .I0(level3_in[1188]),
   .I1(level3_in[1189]),
   .I2(level3_in[1190]),
   .I3(level3_in[1191]),
   .I4(level3_in[1192]),
   .I5(level3_in[1193])
);

LUT6 #(
   .INIT(64'h3232b9c73232b9c7)  
) LUT6_inst9271 (
   .O(to_level2[199]),
   .I0(level3_in[1194]),
   .I1(level3_in[1195]),
   .I2(level3_in[1196]),
   .I3(level3_in[1197]),
   .I4(level3_in[1198]),
   .I5(level3_in[1199])
);

LUT6 #(
   .INIT(64'h36d0bfad36d0bfad)  
) LUT6_inst9272 (
   .O(to_level2[200]),
   .I0(level3_in[1200]),
   .I1(level3_in[1201]),
   .I2(level3_in[1202]),
   .I3(level3_in[1203]),
   .I4(level3_in[1204]),
   .I5(level3_in[1205])
);

LUT6 #(
   .INIT(64'hfd5ed7d2fd5ed7d2)  
) LUT6_inst9273 (
   .O(to_level2[201]),
   .I0(level3_in[1206]),
   .I1(level3_in[1207]),
   .I2(level3_in[1208]),
   .I3(level3_in[1209]),
   .I4(level3_in[1210]),
   .I5(level3_in[1211])
);

LUT6 #(
   .INIT(64'h0479d03a0479d03a)  
) LUT6_inst9274 (
   .O(to_level2[202]),
   .I0(level3_in[1212]),
   .I1(level3_in[1213]),
   .I2(level3_in[1214]),
   .I3(level3_in[1215]),
   .I4(level3_in[1216]),
   .I5(level3_in[1217])
);

LUT6 #(
   .INIT(64'h3a1a0c9e3a1a0c9e)  
) LUT6_inst9275 (
   .O(to_level2[203]),
   .I0(level3_in[1218]),
   .I1(level3_in[1219]),
   .I2(level3_in[1220]),
   .I3(level3_in[1221]),
   .I4(level3_in[1222]),
   .I5(level3_in[1223])
);

LUT6 #(
   .INIT(64'h6a88a89e6a88a89e)  
) LUT6_inst9276 (
   .O(to_level2[204]),
   .I0(level3_in[1224]),
   .I1(level3_in[1225]),
   .I2(level3_in[1226]),
   .I3(level3_in[1227]),
   .I4(level3_in[1228]),
   .I5(level3_in[1229])
);

LUT6 #(
   .INIT(64'hd817faa0d817faa0)  
) LUT6_inst9277 (
   .O(to_level2[205]),
   .I0(level3_in[1230]),
   .I1(level3_in[1231]),
   .I2(level3_in[1232]),
   .I3(level3_in[1233]),
   .I4(level3_in[1234]),
   .I5(level3_in[1235])
);

LUT6 #(
   .INIT(64'hdce10e9cdce10e9c)  
) LUT6_inst9278 (
   .O(to_level2[206]),
   .I0(level3_in[1236]),
   .I1(level3_in[1237]),
   .I2(level3_in[1238]),
   .I3(level3_in[1239]),
   .I4(level3_in[1240]),
   .I5(level3_in[1241])
);

LUT6 #(
   .INIT(64'h7659eb1e7659eb1e)  
) LUT6_inst9279 (
   .O(to_level2[207]),
   .I0(level3_in[1242]),
   .I1(level3_in[1243]),
   .I2(level3_in[1244]),
   .I3(level3_in[1245]),
   .I4(level3_in[1246]),
   .I5(level3_in[1247])
);

LUT6 #(
   .INIT(64'h9b5271b19b5271b1)  
) LUT6_inst9280 (
   .O(to_level2[208]),
   .I0(level3_in[1248]),
   .I1(level3_in[1249]),
   .I2(level3_in[1250]),
   .I3(level3_in[1251]),
   .I4(level3_in[1252]),
   .I5(level3_in[1253])
);

LUT6 #(
   .INIT(64'hac2f8f79ac2f8f79)  
) LUT6_inst9281 (
   .O(to_level2[209]),
   .I0(level3_in[1254]),
   .I1(level3_in[1255]),
   .I2(level3_in[1256]),
   .I3(level3_in[1257]),
   .I4(level3_in[1258]),
   .I5(level3_in[1259])
);

LUT6 #(
   .INIT(64'hea9a2dc6ea9a2dc6)  
) LUT6_inst9282 (
   .O(to_level2[210]),
   .I0(level3_in[1260]),
   .I1(level3_in[1261]),
   .I2(level3_in[1262]),
   .I3(level3_in[1263]),
   .I4(level3_in[1264]),
   .I5(level3_in[1265])
);

LUT6 #(
   .INIT(64'ha14271b8a14271b8)  
) LUT6_inst9283 (
   .O(to_level2[211]),
   .I0(level3_in[1266]),
   .I1(level3_in[1267]),
   .I2(level3_in[1268]),
   .I3(level3_in[1269]),
   .I4(level3_in[1270]),
   .I5(level3_in[1271])
);

LUT6 #(
   .INIT(64'hce520b50ce520b50)  
) LUT6_inst9284 (
   .O(to_level2[212]),
   .I0(level3_in[1272]),
   .I1(level3_in[1273]),
   .I2(level3_in[1274]),
   .I3(level3_in[1275]),
   .I4(level3_in[1276]),
   .I5(level3_in[1277])
);

LUT6 #(
   .INIT(64'h0e5a03a20e5a03a2)  
) LUT6_inst9285 (
   .O(to_level2[213]),
   .I0(level3_in[1278]),
   .I1(level3_in[1279]),
   .I2(level3_in[1280]),
   .I3(level3_in[1281]),
   .I4(level3_in[1282]),
   .I5(level3_in[1283])
);

LUT6 #(
   .INIT(64'ha7abe579a7abe579)  
) LUT6_inst9286 (
   .O(to_level2[214]),
   .I0(level3_in[1284]),
   .I1(level3_in[1285]),
   .I2(level3_in[1286]),
   .I3(level3_in[1287]),
   .I4(level3_in[1288]),
   .I5(level3_in[1289])
);

LUT6 #(
   .INIT(64'h5e9998c45e9998c4)  
) LUT6_inst9287 (
   .O(to_level2[215]),
   .I0(level3_in[1290]),
   .I1(level3_in[1291]),
   .I2(level3_in[1292]),
   .I3(level3_in[1293]),
   .I4(level3_in[1294]),
   .I5(level3_in[1295])
);
////////////// level 2 starts below:/n
LUT6 #(
   .INIT(64'h04e5a68804e5a688)  
) LUT6_inst9288 (
   .O(to_level1[0]),
   .I0(level2_in[0]),
   .I1(level2_in[1]),
   .I2(level2_in[2]),
   .I3(level2_in[3]),
   .I4(level2_in[4]),
   .I5(level2_in[5])
);

LUT6 #(
   .INIT(64'hbf389f82bf389f82)  
) LUT6_inst9289 (
   .O(to_level1[1]),
   .I0(level2_in[6]),
   .I1(level2_in[7]),
   .I2(level2_in[8]),
   .I3(level2_in[9]),
   .I4(level2_in[10]),
   .I5(level2_in[11])
);

LUT6 #(
   .INIT(64'he6db605de6db605d)  
) LUT6_inst9290 (
   .O(to_level1[2]),
   .I0(level2_in[12]),
   .I1(level2_in[13]),
   .I2(level2_in[14]),
   .I3(level2_in[15]),
   .I4(level2_in[16]),
   .I5(level2_in[17])
);

LUT6 #(
   .INIT(64'h787cda6b787cda6b)  
) LUT6_inst9291 (
   .O(to_level1[3]),
   .I0(level2_in[18]),
   .I1(level2_in[19]),
   .I2(level2_in[20]),
   .I3(level2_in[21]),
   .I4(level2_in[22]),
   .I5(level2_in[23])
);

LUT6 #(
   .INIT(64'ha4e9755ba4e9755b)  
) LUT6_inst9292 (
   .O(to_level1[4]),
   .I0(level2_in[24]),
   .I1(level2_in[25]),
   .I2(level2_in[26]),
   .I3(level2_in[27]),
   .I4(level2_in[28]),
   .I5(level2_in[29])
);

LUT6 #(
   .INIT(64'hb5953e26b5953e26)  
) LUT6_inst9293 (
   .O(to_level1[5]),
   .I0(level2_in[30]),
   .I1(level2_in[31]),
   .I2(level2_in[32]),
   .I3(level2_in[33]),
   .I4(level2_in[34]),
   .I5(level2_in[35])
);

LUT6 #(
   .INIT(64'h552b95cf552b95cf)  
) LUT6_inst9294 (
   .O(to_level1[6]),
   .I0(level2_in[36]),
   .I1(level2_in[37]),
   .I2(level2_in[38]),
   .I3(level2_in[39]),
   .I4(level2_in[40]),
   .I5(level2_in[41])
);

LUT6 #(
   .INIT(64'h024554bc024554bc)  
) LUT6_inst9295 (
   .O(to_level1[7]),
   .I0(level2_in[42]),
   .I1(level2_in[43]),
   .I2(level2_in[44]),
   .I3(level2_in[45]),
   .I4(level2_in[46]),
   .I5(level2_in[47])
);

LUT6 #(
   .INIT(64'hfd9518cefd9518ce)  
) LUT6_inst9296 (
   .O(to_level1[8]),
   .I0(level2_in[48]),
   .I1(level2_in[49]),
   .I2(level2_in[50]),
   .I3(level2_in[51]),
   .I4(level2_in[52]),
   .I5(level2_in[53])
);

LUT6 #(
   .INIT(64'h019b4c90019b4c90)  
) LUT6_inst9297 (
   .O(to_level1[9]),
   .I0(level2_in[54]),
   .I1(level2_in[55]),
   .I2(level2_in[56]),
   .I3(level2_in[57]),
   .I4(level2_in[58]),
   .I5(level2_in[59])
);

LUT6 #(
   .INIT(64'h161af14e161af14e)  
) LUT6_inst9298 (
   .O(to_level1[10]),
   .I0(level2_in[60]),
   .I1(level2_in[61]),
   .I2(level2_in[62]),
   .I3(level2_in[63]),
   .I4(level2_in[64]),
   .I5(level2_in[65])
);

LUT6 #(
   .INIT(64'h291df2cc291df2cc)  
) LUT6_inst9299 (
   .O(to_level1[11]),
   .I0(level2_in[66]),
   .I1(level2_in[67]),
   .I2(level2_in[68]),
   .I3(level2_in[69]),
   .I4(level2_in[70]),
   .I5(level2_in[71])
);

LUT6 #(
   .INIT(64'h989df19e989df19e)  
) LUT6_inst9300 (
   .O(to_level1[12]),
   .I0(level2_in[72]),
   .I1(level2_in[73]),
   .I2(level2_in[74]),
   .I3(level2_in[75]),
   .I4(level2_in[76]),
   .I5(level2_in[77])
);

LUT6 #(
   .INIT(64'hece107e6ece107e6)  
) LUT6_inst9301 (
   .O(to_level1[13]),
   .I0(level2_in[78]),
   .I1(level2_in[79]),
   .I2(level2_in[80]),
   .I3(level2_in[81]),
   .I4(level2_in[82]),
   .I5(level2_in[83])
);

LUT6 #(
   .INIT(64'h4663cb214663cb21)  
) LUT6_inst9302 (
   .O(to_level1[14]),
   .I0(level2_in[84]),
   .I1(level2_in[85]),
   .I2(level2_in[86]),
   .I3(level2_in[87]),
   .I4(level2_in[88]),
   .I5(level2_in[89])
);

LUT6 #(
   .INIT(64'h13273f7213273f72)  
) LUT6_inst9303 (
   .O(to_level1[15]),
   .I0(level2_in[90]),
   .I1(level2_in[91]),
   .I2(level2_in[92]),
   .I3(level2_in[93]),
   .I4(level2_in[94]),
   .I5(level2_in[95])
);

LUT6 #(
   .INIT(64'h470323a9470323a9)  
) LUT6_inst9304 (
   .O(to_level1[16]),
   .I0(level2_in[96]),
   .I1(level2_in[97]),
   .I2(level2_in[98]),
   .I3(level2_in[99]),
   .I4(level2_in[100]),
   .I5(level2_in[101])
);

LUT6 #(
   .INIT(64'hc79749d2c79749d2)  
) LUT6_inst9305 (
   .O(to_level1[17]),
   .I0(level2_in[102]),
   .I1(level2_in[103]),
   .I2(level2_in[104]),
   .I3(level2_in[105]),
   .I4(level2_in[106]),
   .I5(level2_in[107])
);

LUT6 #(
   .INIT(64'h2c6de18f2c6de18f)  
) LUT6_inst9306 (
   .O(to_level1[18]),
   .I0(level2_in[108]),
   .I1(level2_in[109]),
   .I2(level2_in[110]),
   .I3(level2_in[111]),
   .I4(level2_in[112]),
   .I5(level2_in[113])
);

LUT6 #(
   .INIT(64'h7c35388a7c35388a)  
) LUT6_inst9307 (
   .O(to_level1[19]),
   .I0(level2_in[114]),
   .I1(level2_in[115]),
   .I2(level2_in[116]),
   .I3(level2_in[117]),
   .I4(level2_in[118]),
   .I5(level2_in[119])
);

LUT6 #(
   .INIT(64'he2454192e2454192)  
) LUT6_inst9308 (
   .O(to_level1[20]),
   .I0(level2_in[120]),
   .I1(level2_in[121]),
   .I2(level2_in[122]),
   .I3(level2_in[123]),
   .I4(level2_in[124]),
   .I5(level2_in[125])
);

LUT6 #(
   .INIT(64'h2b0e70332b0e7033)  
) LUT6_inst9309 (
   .O(to_level1[21]),
   .I0(level2_in[126]),
   .I1(level2_in[127]),
   .I2(level2_in[128]),
   .I3(level2_in[129]),
   .I4(level2_in[130]),
   .I5(level2_in[131])
);

LUT6 #(
   .INIT(64'h34dccc9834dccc98)  
) LUT6_inst9310 (
   .O(to_level1[22]),
   .I0(level2_in[132]),
   .I1(level2_in[133]),
   .I2(level2_in[134]),
   .I3(level2_in[135]),
   .I4(level2_in[136]),
   .I5(level2_in[137])
);

LUT6 #(
   .INIT(64'hcb62ccd7cb62ccd7)  
) LUT6_inst9311 (
   .O(to_level1[23]),
   .I0(level2_in[138]),
   .I1(level2_in[139]),
   .I2(level2_in[140]),
   .I3(level2_in[141]),
   .I4(level2_in[142]),
   .I5(level2_in[143])
);

LUT6 #(
   .INIT(64'h7c4caf027c4caf02)  
) LUT6_inst9312 (
   .O(to_level1[24]),
   .I0(level2_in[144]),
   .I1(level2_in[145]),
   .I2(level2_in[146]),
   .I3(level2_in[147]),
   .I4(level2_in[148]),
   .I5(level2_in[149])
);

LUT6 #(
   .INIT(64'hcb2fabcccb2fabcc)  
) LUT6_inst9313 (
   .O(to_level1[25]),
   .I0(level2_in[150]),
   .I1(level2_in[151]),
   .I2(level2_in[152]),
   .I3(level2_in[153]),
   .I4(level2_in[154]),
   .I5(level2_in[155])
);

LUT6 #(
   .INIT(64'h15a1a86e15a1a86e)  
) LUT6_inst9314 (
   .O(to_level1[26]),
   .I0(level2_in[156]),
   .I1(level2_in[157]),
   .I2(level2_in[158]),
   .I3(level2_in[159]),
   .I4(level2_in[160]),
   .I5(level2_in[161])
);

LUT6 #(
   .INIT(64'hdd6959eddd6959ed)  
) LUT6_inst9315 (
   .O(to_level1[27]),
   .I0(level2_in[162]),
   .I1(level2_in[163]),
   .I2(level2_in[164]),
   .I3(level2_in[165]),
   .I4(level2_in[166]),
   .I5(level2_in[167])
);

LUT6 #(
   .INIT(64'h4f4050664f405066)  
) LUT6_inst9316 (
   .O(to_level1[28]),
   .I0(level2_in[168]),
   .I1(level2_in[169]),
   .I2(level2_in[170]),
   .I3(level2_in[171]),
   .I4(level2_in[172]),
   .I5(level2_in[173])
);

LUT6 #(
   .INIT(64'h7114c7f57114c7f5)  
) LUT6_inst9317 (
   .O(to_level1[29]),
   .I0(level2_in[174]),
   .I1(level2_in[175]),
   .I2(level2_in[176]),
   .I3(level2_in[177]),
   .I4(level2_in[178]),
   .I5(level2_in[179])
);

LUT6 #(
   .INIT(64'h8e6853d88e6853d8)  
) LUT6_inst9318 (
   .O(to_level1[30]),
   .I0(level2_in[180]),
   .I1(level2_in[181]),
   .I2(level2_in[182]),
   .I3(level2_in[183]),
   .I4(level2_in[184]),
   .I5(level2_in[185])
);

LUT6 #(
   .INIT(64'h9bff0b589bff0b58)  
) LUT6_inst9319 (
   .O(to_level1[31]),
   .I0(level2_in[186]),
   .I1(level2_in[187]),
   .I2(level2_in[188]),
   .I3(level2_in[189]),
   .I4(level2_in[190]),
   .I5(level2_in[191])
);

LUT6 #(
   .INIT(64'h8ee40a1f8ee40a1f)  
) LUT6_inst9320 (
   .O(to_level1[32]),
   .I0(level2_in[192]),
   .I1(level2_in[193]),
   .I2(level2_in[194]),
   .I3(level2_in[195]),
   .I4(level2_in[196]),
   .I5(level2_in[197])
);

LUT6 #(
   .INIT(64'h4090336b4090336b)  
) LUT6_inst9321 (
   .O(to_level1[33]),
   .I0(level2_in[198]),
   .I1(level2_in[199]),
   .I2(level2_in[200]),
   .I3(level2_in[201]),
   .I4(level2_in[202]),
   .I5(level2_in[203])
);

LUT6 #(
   .INIT(64'h76fb38c076fb38c0)  
) LUT6_inst9322 (
   .O(to_level1[34]),
   .I0(level2_in[204]),
   .I1(level2_in[205]),
   .I2(level2_in[206]),
   .I3(level2_in[207]),
   .I4(level2_in[208]),
   .I5(level2_in[209])
);

LUT6 #(
   .INIT(64'h2298a3942298a394)  
) LUT6_inst9323 (
   .O(to_level1[35]),
   .I0(level2_in[210]),
   .I1(level2_in[211]),
   .I2(level2_in[212]),
   .I3(level2_in[213]),
   .I4(level2_in[214]),
   .I5(level2_in[215])
);
////////////// level 1 starts below:/n
LUT6 #(
   .INIT(64'hd567f163d567f163)  
) LUT6_inst9324 (
   .O(to_level0[0]),
   .I0(level1_in[0]),
   .I1(level1_in[1]),
   .I2(level1_in[2]),
   .I3(level1_in[3]),
   .I4(level1_in[4]),
   .I5(level1_in[5])
);

LUT6 #(
   .INIT(64'h64c40f6e64c40f6e)  
) LUT6_inst9325 (
   .O(to_level0[1]),
   .I0(level1_in[6]),
   .I1(level1_in[7]),
   .I2(level1_in[8]),
   .I3(level1_in[9]),
   .I4(level1_in[10]),
   .I5(level1_in[11])
);

LUT6 #(
   .INIT(64'h0ca095f80ca095f8)  
) LUT6_inst9326 (
   .O(to_level0[2]),
   .I0(level1_in[12]),
   .I1(level1_in[13]),
   .I2(level1_in[14]),
   .I3(level1_in[15]),
   .I4(level1_in[16]),
   .I5(level1_in[17])
);

LUT6 #(
   .INIT(64'hcb1291e6cb1291e6)  
) LUT6_inst9327 (
   .O(to_level0[3]),
   .I0(level1_in[18]),
   .I1(level1_in[19]),
   .I2(level1_in[20]),
   .I3(level1_in[21]),
   .I4(level1_in[22]),
   .I5(level1_in[23])
);

LUT6 #(
   .INIT(64'he8251b8be8251b8b)  
) LUT6_inst9328 (
   .O(to_level0[4]),
   .I0(level1_in[24]),
   .I1(level1_in[25]),
   .I2(level1_in[26]),
   .I3(level1_in[27]),
   .I4(level1_in[28]),
   .I5(level1_in[29])
);

LUT6 #(
   .INIT(64'h12fe095412fe0954)  
) LUT6_inst9329 (
   .O(to_level0[5]),
   .I0(level1_in[30]),
   .I1(level1_in[31]),
   .I2(level1_in[32]),
   .I3(level1_in[33]),
   .I4(level1_in[34]),
   .I5(level1_in[35])
);
////////////// level 0 starts below:/n
LUT6 #(
   .INIT(64'h6a2919146a291914)  
) LUT6_inst9330 (
   .O(data_out_temp),
   .I0(level0_in[0]),
   .I1(level0_in[1]),
   .I2(level0_in[2]),
   .I3(level0_in[3]),
   .I4(level0_in[4]),
   .I5(level0_in[5])
);

endmodule