
module lut_4level_tree6(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [7775:0] data_in,
                       input       data_valid,
                       output  reg data_out     
                       );

wire    [7775:0] to_level4;
(*S="TRUE"*)reg     [7775:0] level4_in;
wire    [1295:0] to_level3;
(*S="TRUE"*)reg     [1295:0] level3_in;
wire    [215:0] to_level2;
(*S="TRUE"*)reg     [215:0] level2_in;
wire    [35:0] to_level1;
(*S="TRUE"*)reg     [35:0] level1_in;
wire    [5:0] to_level0;
(*S="TRUE"*)reg     [5:0] level0_in;
wire          data_out_temp;


assign  to_level4 = data_in;

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level4_in <= 7776'b0;
  else
    level4_in <= to_level4;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level3_in <= 1296'b0;
  else
    level3_in <= to_level3;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level2_in <= 216'b0;
  else
    level2_in <= to_level2;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level1_in <= 36'b0;
  else
    level1_in <= to_level1;
end


always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    level0_in <= 6'b0;
  else
    level0_in <= to_level0;
end

always @(posedge rx_fifo_clock)
begin
  if(!rx_fifo_resetn)
    data_out <= 1'b0;
  else
    if(data_valid == 1'b1)
      data_out <= data_out_temp;
    else;
end
////////////// level 4 starts below:/n
LUT6 #(
   .INIT(64'h7859d2527859d252)  
) LUT6_inst7776 (
   .O(to_level3[0]),
   .I0(level4_in[0]),
   .I1(level4_in[1]),
   .I2(level4_in[2]),
   .I3(level4_in[3]),
   .I4(level4_in[4]),
   .I5(level4_in[5])
);

LUT6 #(
   .INIT(64'h235ebcff235ebcff)  
) LUT6_inst7777 (
   .O(to_level3[1]),
   .I0(level4_in[6]),
   .I1(level4_in[7]),
   .I2(level4_in[8]),
   .I3(level4_in[9]),
   .I4(level4_in[10]),
   .I5(level4_in[11])
);

LUT6 #(
   .INIT(64'h938a7127938a7127)  
) LUT6_inst7778 (
   .O(to_level3[2]),
   .I0(level4_in[12]),
   .I1(level4_in[13]),
   .I2(level4_in[14]),
   .I3(level4_in[15]),
   .I4(level4_in[16]),
   .I5(level4_in[17])
);

LUT6 #(
   .INIT(64'h06dcb79206dcb792)  
) LUT6_inst7779 (
   .O(to_level3[3]),
   .I0(level4_in[18]),
   .I1(level4_in[19]),
   .I2(level4_in[20]),
   .I3(level4_in[21]),
   .I4(level4_in[22]),
   .I5(level4_in[23])
);

LUT6 #(
   .INIT(64'h4160ac4c4160ac4c)  
) LUT6_inst7780 (
   .O(to_level3[4]),
   .I0(level4_in[24]),
   .I1(level4_in[25]),
   .I2(level4_in[26]),
   .I3(level4_in[27]),
   .I4(level4_in[28]),
   .I5(level4_in[29])
);

LUT6 #(
   .INIT(64'hb982610fb982610f)  
) LUT6_inst7781 (
   .O(to_level3[5]),
   .I0(level4_in[30]),
   .I1(level4_in[31]),
   .I2(level4_in[32]),
   .I3(level4_in[33]),
   .I4(level4_in[34]),
   .I5(level4_in[35])
);

LUT6 #(
   .INIT(64'hdc57c3c7dc57c3c7)  
) LUT6_inst7782 (
   .O(to_level3[6]),
   .I0(level4_in[36]),
   .I1(level4_in[37]),
   .I2(level4_in[38]),
   .I3(level4_in[39]),
   .I4(level4_in[40]),
   .I5(level4_in[41])
);

LUT6 #(
   .INIT(64'h48b590d048b590d0)  
) LUT6_inst7783 (
   .O(to_level3[7]),
   .I0(level4_in[42]),
   .I1(level4_in[43]),
   .I2(level4_in[44]),
   .I3(level4_in[45]),
   .I4(level4_in[46]),
   .I5(level4_in[47])
);

LUT6 #(
   .INIT(64'h893bda1b893bda1b)  
) LUT6_inst7784 (
   .O(to_level3[8]),
   .I0(level4_in[48]),
   .I1(level4_in[49]),
   .I2(level4_in[50]),
   .I3(level4_in[51]),
   .I4(level4_in[52]),
   .I5(level4_in[53])
);

LUT6 #(
   .INIT(64'h867e8493867e8493)  
) LUT6_inst7785 (
   .O(to_level3[9]),
   .I0(level4_in[54]),
   .I1(level4_in[55]),
   .I2(level4_in[56]),
   .I3(level4_in[57]),
   .I4(level4_in[58]),
   .I5(level4_in[59])
);

LUT6 #(
   .INIT(64'h604b9232604b9232)  
) LUT6_inst7786 (
   .O(to_level3[10]),
   .I0(level4_in[60]),
   .I1(level4_in[61]),
   .I2(level4_in[62]),
   .I3(level4_in[63]),
   .I4(level4_in[64]),
   .I5(level4_in[65])
);

LUT6 #(
   .INIT(64'h56216c1d56216c1d)  
) LUT6_inst7787 (
   .O(to_level3[11]),
   .I0(level4_in[66]),
   .I1(level4_in[67]),
   .I2(level4_in[68]),
   .I3(level4_in[69]),
   .I4(level4_in[70]),
   .I5(level4_in[71])
);

LUT6 #(
   .INIT(64'ha599b3d1a599b3d1)  
) LUT6_inst7788 (
   .O(to_level3[12]),
   .I0(level4_in[72]),
   .I1(level4_in[73]),
   .I2(level4_in[74]),
   .I3(level4_in[75]),
   .I4(level4_in[76]),
   .I5(level4_in[77])
);

LUT6 #(
   .INIT(64'hb218483bb218483b)  
) LUT6_inst7789 (
   .O(to_level3[13]),
   .I0(level4_in[78]),
   .I1(level4_in[79]),
   .I2(level4_in[80]),
   .I3(level4_in[81]),
   .I4(level4_in[82]),
   .I5(level4_in[83])
);

LUT6 #(
   .INIT(64'ha0c3a56aa0c3a56a)  
) LUT6_inst7790 (
   .O(to_level3[14]),
   .I0(level4_in[84]),
   .I1(level4_in[85]),
   .I2(level4_in[86]),
   .I3(level4_in[87]),
   .I4(level4_in[88]),
   .I5(level4_in[89])
);

LUT6 #(
   .INIT(64'h0a4c58440a4c5844)  
) LUT6_inst7791 (
   .O(to_level3[15]),
   .I0(level4_in[90]),
   .I1(level4_in[91]),
   .I2(level4_in[92]),
   .I3(level4_in[93]),
   .I4(level4_in[94]),
   .I5(level4_in[95])
);

LUT6 #(
   .INIT(64'h1e992d711e992d71)  
) LUT6_inst7792 (
   .O(to_level3[16]),
   .I0(level4_in[96]),
   .I1(level4_in[97]),
   .I2(level4_in[98]),
   .I3(level4_in[99]),
   .I4(level4_in[100]),
   .I5(level4_in[101])
);

LUT6 #(
   .INIT(64'hdbd1c21adbd1c21a)  
) LUT6_inst7793 (
   .O(to_level3[17]),
   .I0(level4_in[102]),
   .I1(level4_in[103]),
   .I2(level4_in[104]),
   .I3(level4_in[105]),
   .I4(level4_in[106]),
   .I5(level4_in[107])
);

LUT6 #(
   .INIT(64'h23bb246723bb2467)  
) LUT6_inst7794 (
   .O(to_level3[18]),
   .I0(level4_in[108]),
   .I1(level4_in[109]),
   .I2(level4_in[110]),
   .I3(level4_in[111]),
   .I4(level4_in[112]),
   .I5(level4_in[113])
);

LUT6 #(
   .INIT(64'h59ad312159ad3121)  
) LUT6_inst7795 (
   .O(to_level3[19]),
   .I0(level4_in[114]),
   .I1(level4_in[115]),
   .I2(level4_in[116]),
   .I3(level4_in[117]),
   .I4(level4_in[118]),
   .I5(level4_in[119])
);

LUT6 #(
   .INIT(64'h89e1d0e589e1d0e5)  
) LUT6_inst7796 (
   .O(to_level3[20]),
   .I0(level4_in[120]),
   .I1(level4_in[121]),
   .I2(level4_in[122]),
   .I3(level4_in[123]),
   .I4(level4_in[124]),
   .I5(level4_in[125])
);

LUT6 #(
   .INIT(64'h6966a8986966a898)  
) LUT6_inst7797 (
   .O(to_level3[21]),
   .I0(level4_in[126]),
   .I1(level4_in[127]),
   .I2(level4_in[128]),
   .I3(level4_in[129]),
   .I4(level4_in[130]),
   .I5(level4_in[131])
);

LUT6 #(
   .INIT(64'hb85805f4b85805f4)  
) LUT6_inst7798 (
   .O(to_level3[22]),
   .I0(level4_in[132]),
   .I1(level4_in[133]),
   .I2(level4_in[134]),
   .I3(level4_in[135]),
   .I4(level4_in[136]),
   .I5(level4_in[137])
);

LUT6 #(
   .INIT(64'h8e6984778e698477)  
) LUT6_inst7799 (
   .O(to_level3[23]),
   .I0(level4_in[138]),
   .I1(level4_in[139]),
   .I2(level4_in[140]),
   .I3(level4_in[141]),
   .I4(level4_in[142]),
   .I5(level4_in[143])
);

LUT6 #(
   .INIT(64'hd178f4fad178f4fa)  
) LUT6_inst7800 (
   .O(to_level3[24]),
   .I0(level4_in[144]),
   .I1(level4_in[145]),
   .I2(level4_in[146]),
   .I3(level4_in[147]),
   .I4(level4_in[148]),
   .I5(level4_in[149])
);

LUT6 #(
   .INIT(64'h2e0310c32e0310c3)  
) LUT6_inst7801 (
   .O(to_level3[25]),
   .I0(level4_in[150]),
   .I1(level4_in[151]),
   .I2(level4_in[152]),
   .I3(level4_in[153]),
   .I4(level4_in[154]),
   .I5(level4_in[155])
);

LUT6 #(
   .INIT(64'h3850d0d03850d0d0)  
) LUT6_inst7802 (
   .O(to_level3[26]),
   .I0(level4_in[156]),
   .I1(level4_in[157]),
   .I2(level4_in[158]),
   .I3(level4_in[159]),
   .I4(level4_in[160]),
   .I5(level4_in[161])
);

LUT6 #(
   .INIT(64'hced050cdced050cd)  
) LUT6_inst7803 (
   .O(to_level3[27]),
   .I0(level4_in[162]),
   .I1(level4_in[163]),
   .I2(level4_in[164]),
   .I3(level4_in[165]),
   .I4(level4_in[166]),
   .I5(level4_in[167])
);

LUT6 #(
   .INIT(64'h0c9081510c908151)  
) LUT6_inst7804 (
   .O(to_level3[28]),
   .I0(level4_in[168]),
   .I1(level4_in[169]),
   .I2(level4_in[170]),
   .I3(level4_in[171]),
   .I4(level4_in[172]),
   .I5(level4_in[173])
);

LUT6 #(
   .INIT(64'h005f2fda005f2fda)  
) LUT6_inst7805 (
   .O(to_level3[29]),
   .I0(level4_in[174]),
   .I1(level4_in[175]),
   .I2(level4_in[176]),
   .I3(level4_in[177]),
   .I4(level4_in[178]),
   .I5(level4_in[179])
);

LUT6 #(
   .INIT(64'hb4c2efcfb4c2efcf)  
) LUT6_inst7806 (
   .O(to_level3[30]),
   .I0(level4_in[180]),
   .I1(level4_in[181]),
   .I2(level4_in[182]),
   .I3(level4_in[183]),
   .I4(level4_in[184]),
   .I5(level4_in[185])
);

LUT6 #(
   .INIT(64'hb6bf74aeb6bf74ae)  
) LUT6_inst7807 (
   .O(to_level3[31]),
   .I0(level4_in[186]),
   .I1(level4_in[187]),
   .I2(level4_in[188]),
   .I3(level4_in[189]),
   .I4(level4_in[190]),
   .I5(level4_in[191])
);

LUT6 #(
   .INIT(64'h2626ffa12626ffa1)  
) LUT6_inst7808 (
   .O(to_level3[32]),
   .I0(level4_in[192]),
   .I1(level4_in[193]),
   .I2(level4_in[194]),
   .I3(level4_in[195]),
   .I4(level4_in[196]),
   .I5(level4_in[197])
);

LUT6 #(
   .INIT(64'h026b6d93026b6d93)  
) LUT6_inst7809 (
   .O(to_level3[33]),
   .I0(level4_in[198]),
   .I1(level4_in[199]),
   .I2(level4_in[200]),
   .I3(level4_in[201]),
   .I4(level4_in[202]),
   .I5(level4_in[203])
);

LUT6 #(
   .INIT(64'h752a094a752a094a)  
) LUT6_inst7810 (
   .O(to_level3[34]),
   .I0(level4_in[204]),
   .I1(level4_in[205]),
   .I2(level4_in[206]),
   .I3(level4_in[207]),
   .I4(level4_in[208]),
   .I5(level4_in[209])
);

LUT6 #(
   .INIT(64'hdc605d89dc605d89)  
) LUT6_inst7811 (
   .O(to_level3[35]),
   .I0(level4_in[210]),
   .I1(level4_in[211]),
   .I2(level4_in[212]),
   .I3(level4_in[213]),
   .I4(level4_in[214]),
   .I5(level4_in[215])
);

LUT6 #(
   .INIT(64'h8645a7658645a765)  
) LUT6_inst7812 (
   .O(to_level3[36]),
   .I0(level4_in[216]),
   .I1(level4_in[217]),
   .I2(level4_in[218]),
   .I3(level4_in[219]),
   .I4(level4_in[220]),
   .I5(level4_in[221])
);

LUT6 #(
   .INIT(64'h7d7a11097d7a1109)  
) LUT6_inst7813 (
   .O(to_level3[37]),
   .I0(level4_in[222]),
   .I1(level4_in[223]),
   .I2(level4_in[224]),
   .I3(level4_in[225]),
   .I4(level4_in[226]),
   .I5(level4_in[227])
);

LUT6 #(
   .INIT(64'hdd62d9eddd62d9ed)  
) LUT6_inst7814 (
   .O(to_level3[38]),
   .I0(level4_in[228]),
   .I1(level4_in[229]),
   .I2(level4_in[230]),
   .I3(level4_in[231]),
   .I4(level4_in[232]),
   .I5(level4_in[233])
);

LUT6 #(
   .INIT(64'h0c5a0ca40c5a0ca4)  
) LUT6_inst7815 (
   .O(to_level3[39]),
   .I0(level4_in[234]),
   .I1(level4_in[235]),
   .I2(level4_in[236]),
   .I3(level4_in[237]),
   .I4(level4_in[238]),
   .I5(level4_in[239])
);

LUT6 #(
   .INIT(64'ha895541ca895541c)  
) LUT6_inst7816 (
   .O(to_level3[40]),
   .I0(level4_in[240]),
   .I1(level4_in[241]),
   .I2(level4_in[242]),
   .I3(level4_in[243]),
   .I4(level4_in[244]),
   .I5(level4_in[245])
);

LUT6 #(
   .INIT(64'h948633e9948633e9)  
) LUT6_inst7817 (
   .O(to_level3[41]),
   .I0(level4_in[246]),
   .I1(level4_in[247]),
   .I2(level4_in[248]),
   .I3(level4_in[249]),
   .I4(level4_in[250]),
   .I5(level4_in[251])
);

LUT6 #(
   .INIT(64'h57be88ec57be88ec)  
) LUT6_inst7818 (
   .O(to_level3[42]),
   .I0(level4_in[252]),
   .I1(level4_in[253]),
   .I2(level4_in[254]),
   .I3(level4_in[255]),
   .I4(level4_in[256]),
   .I5(level4_in[257])
);

LUT6 #(
   .INIT(64'h3fbf52563fbf5256)  
) LUT6_inst7819 (
   .O(to_level3[43]),
   .I0(level4_in[258]),
   .I1(level4_in[259]),
   .I2(level4_in[260]),
   .I3(level4_in[261]),
   .I4(level4_in[262]),
   .I5(level4_in[263])
);

LUT6 #(
   .INIT(64'h252a9f0a252a9f0a)  
) LUT6_inst7820 (
   .O(to_level3[44]),
   .I0(level4_in[264]),
   .I1(level4_in[265]),
   .I2(level4_in[266]),
   .I3(level4_in[267]),
   .I4(level4_in[268]),
   .I5(level4_in[269])
);

LUT6 #(
   .INIT(64'h01b93be801b93be8)  
) LUT6_inst7821 (
   .O(to_level3[45]),
   .I0(level4_in[270]),
   .I1(level4_in[271]),
   .I2(level4_in[272]),
   .I3(level4_in[273]),
   .I4(level4_in[274]),
   .I5(level4_in[275])
);

LUT6 #(
   .INIT(64'ha5f2e2bba5f2e2bb)  
) LUT6_inst7822 (
   .O(to_level3[46]),
   .I0(level4_in[276]),
   .I1(level4_in[277]),
   .I2(level4_in[278]),
   .I3(level4_in[279]),
   .I4(level4_in[280]),
   .I5(level4_in[281])
);

LUT6 #(
   .INIT(64'h83dd9ebd83dd9ebd)  
) LUT6_inst7823 (
   .O(to_level3[47]),
   .I0(level4_in[282]),
   .I1(level4_in[283]),
   .I2(level4_in[284]),
   .I3(level4_in[285]),
   .I4(level4_in[286]),
   .I5(level4_in[287])
);

LUT6 #(
   .INIT(64'hbb34b467bb34b467)  
) LUT6_inst7824 (
   .O(to_level3[48]),
   .I0(level4_in[288]),
   .I1(level4_in[289]),
   .I2(level4_in[290]),
   .I3(level4_in[291]),
   .I4(level4_in[292]),
   .I5(level4_in[293])
);

LUT6 #(
   .INIT(64'h68c9729b68c9729b)  
) LUT6_inst7825 (
   .O(to_level3[49]),
   .I0(level4_in[294]),
   .I1(level4_in[295]),
   .I2(level4_in[296]),
   .I3(level4_in[297]),
   .I4(level4_in[298]),
   .I5(level4_in[299])
);

LUT6 #(
   .INIT(64'ha31b8f65a31b8f65)  
) LUT6_inst7826 (
   .O(to_level3[50]),
   .I0(level4_in[300]),
   .I1(level4_in[301]),
   .I2(level4_in[302]),
   .I3(level4_in[303]),
   .I4(level4_in[304]),
   .I5(level4_in[305])
);

LUT6 #(
   .INIT(64'h2fa1f1ca2fa1f1ca)  
) LUT6_inst7827 (
   .O(to_level3[51]),
   .I0(level4_in[306]),
   .I1(level4_in[307]),
   .I2(level4_in[308]),
   .I3(level4_in[309]),
   .I4(level4_in[310]),
   .I5(level4_in[311])
);

LUT6 #(
   .INIT(64'h51cf6d6151cf6d61)  
) LUT6_inst7828 (
   .O(to_level3[52]),
   .I0(level4_in[312]),
   .I1(level4_in[313]),
   .I2(level4_in[314]),
   .I3(level4_in[315]),
   .I4(level4_in[316]),
   .I5(level4_in[317])
);

LUT6 #(
   .INIT(64'h9597b17f9597b17f)  
) LUT6_inst7829 (
   .O(to_level3[53]),
   .I0(level4_in[318]),
   .I1(level4_in[319]),
   .I2(level4_in[320]),
   .I3(level4_in[321]),
   .I4(level4_in[322]),
   .I5(level4_in[323])
);

LUT6 #(
   .INIT(64'h55b6ad2a55b6ad2a)  
) LUT6_inst7830 (
   .O(to_level3[54]),
   .I0(level4_in[324]),
   .I1(level4_in[325]),
   .I2(level4_in[326]),
   .I3(level4_in[327]),
   .I4(level4_in[328]),
   .I5(level4_in[329])
);

LUT6 #(
   .INIT(64'h84540e8584540e85)  
) LUT6_inst7831 (
   .O(to_level3[55]),
   .I0(level4_in[330]),
   .I1(level4_in[331]),
   .I2(level4_in[332]),
   .I3(level4_in[333]),
   .I4(level4_in[334]),
   .I5(level4_in[335])
);

LUT6 #(
   .INIT(64'h18e5461918e54619)  
) LUT6_inst7832 (
   .O(to_level3[56]),
   .I0(level4_in[336]),
   .I1(level4_in[337]),
   .I2(level4_in[338]),
   .I3(level4_in[339]),
   .I4(level4_in[340]),
   .I5(level4_in[341])
);

LUT6 #(
   .INIT(64'h8bb2a2f68bb2a2f6)  
) LUT6_inst7833 (
   .O(to_level3[57]),
   .I0(level4_in[342]),
   .I1(level4_in[343]),
   .I2(level4_in[344]),
   .I3(level4_in[345]),
   .I4(level4_in[346]),
   .I5(level4_in[347])
);

LUT6 #(
   .INIT(64'he7c8f8fde7c8f8fd)  
) LUT6_inst7834 (
   .O(to_level3[58]),
   .I0(level4_in[348]),
   .I1(level4_in[349]),
   .I2(level4_in[350]),
   .I3(level4_in[351]),
   .I4(level4_in[352]),
   .I5(level4_in[353])
);

LUT6 #(
   .INIT(64'h4a9845c74a9845c7)  
) LUT6_inst7835 (
   .O(to_level3[59]),
   .I0(level4_in[354]),
   .I1(level4_in[355]),
   .I2(level4_in[356]),
   .I3(level4_in[357]),
   .I4(level4_in[358]),
   .I5(level4_in[359])
);

LUT6 #(
   .INIT(64'h296c6b64296c6b64)  
) LUT6_inst7836 (
   .O(to_level3[60]),
   .I0(level4_in[360]),
   .I1(level4_in[361]),
   .I2(level4_in[362]),
   .I3(level4_in[363]),
   .I4(level4_in[364]),
   .I5(level4_in[365])
);

LUT6 #(
   .INIT(64'h6804606368046063)  
) LUT6_inst7837 (
   .O(to_level3[61]),
   .I0(level4_in[366]),
   .I1(level4_in[367]),
   .I2(level4_in[368]),
   .I3(level4_in[369]),
   .I4(level4_in[370]),
   .I5(level4_in[371])
);

LUT6 #(
   .INIT(64'h9e971bb69e971bb6)  
) LUT6_inst7838 (
   .O(to_level3[62]),
   .I0(level4_in[372]),
   .I1(level4_in[373]),
   .I2(level4_in[374]),
   .I3(level4_in[375]),
   .I4(level4_in[376]),
   .I5(level4_in[377])
);

LUT6 #(
   .INIT(64'h0161ab600161ab60)  
) LUT6_inst7839 (
   .O(to_level3[63]),
   .I0(level4_in[378]),
   .I1(level4_in[379]),
   .I2(level4_in[380]),
   .I3(level4_in[381]),
   .I4(level4_in[382]),
   .I5(level4_in[383])
);

LUT6 #(
   .INIT(64'h0415aa3d0415aa3d)  
) LUT6_inst7840 (
   .O(to_level3[64]),
   .I0(level4_in[384]),
   .I1(level4_in[385]),
   .I2(level4_in[386]),
   .I3(level4_in[387]),
   .I4(level4_in[388]),
   .I5(level4_in[389])
);

LUT6 #(
   .INIT(64'h80b5c6f080b5c6f0)  
) LUT6_inst7841 (
   .O(to_level3[65]),
   .I0(level4_in[390]),
   .I1(level4_in[391]),
   .I2(level4_in[392]),
   .I3(level4_in[393]),
   .I4(level4_in[394]),
   .I5(level4_in[395])
);

LUT6 #(
   .INIT(64'he7d21331e7d21331)  
) LUT6_inst7842 (
   .O(to_level3[66]),
   .I0(level4_in[396]),
   .I1(level4_in[397]),
   .I2(level4_in[398]),
   .I3(level4_in[399]),
   .I4(level4_in[400]),
   .I5(level4_in[401])
);

LUT6 #(
   .INIT(64'hd55be2e4d55be2e4)  
) LUT6_inst7843 (
   .O(to_level3[67]),
   .I0(level4_in[402]),
   .I1(level4_in[403]),
   .I2(level4_in[404]),
   .I3(level4_in[405]),
   .I4(level4_in[406]),
   .I5(level4_in[407])
);

LUT6 #(
   .INIT(64'h24918f4224918f42)  
) LUT6_inst7844 (
   .O(to_level3[68]),
   .I0(level4_in[408]),
   .I1(level4_in[409]),
   .I2(level4_in[410]),
   .I3(level4_in[411]),
   .I4(level4_in[412]),
   .I5(level4_in[413])
);

LUT6 #(
   .INIT(64'h627a6ecb627a6ecb)  
) LUT6_inst7845 (
   .O(to_level3[69]),
   .I0(level4_in[414]),
   .I1(level4_in[415]),
   .I2(level4_in[416]),
   .I3(level4_in[417]),
   .I4(level4_in[418]),
   .I5(level4_in[419])
);

LUT6 #(
   .INIT(64'h78b8cf4178b8cf41)  
) LUT6_inst7846 (
   .O(to_level3[70]),
   .I0(level4_in[420]),
   .I1(level4_in[421]),
   .I2(level4_in[422]),
   .I3(level4_in[423]),
   .I4(level4_in[424]),
   .I5(level4_in[425])
);

LUT6 #(
   .INIT(64'h96215d0a96215d0a)  
) LUT6_inst7847 (
   .O(to_level3[71]),
   .I0(level4_in[426]),
   .I1(level4_in[427]),
   .I2(level4_in[428]),
   .I3(level4_in[429]),
   .I4(level4_in[430]),
   .I5(level4_in[431])
);

LUT6 #(
   .INIT(64'h4aba28584aba2858)  
) LUT6_inst7848 (
   .O(to_level3[72]),
   .I0(level4_in[432]),
   .I1(level4_in[433]),
   .I2(level4_in[434]),
   .I3(level4_in[435]),
   .I4(level4_in[436]),
   .I5(level4_in[437])
);

LUT6 #(
   .INIT(64'h846264f7846264f7)  
) LUT6_inst7849 (
   .O(to_level3[73]),
   .I0(level4_in[438]),
   .I1(level4_in[439]),
   .I2(level4_in[440]),
   .I3(level4_in[441]),
   .I4(level4_in[442]),
   .I5(level4_in[443])
);

LUT6 #(
   .INIT(64'h01b1ab7a01b1ab7a)  
) LUT6_inst7850 (
   .O(to_level3[74]),
   .I0(level4_in[444]),
   .I1(level4_in[445]),
   .I2(level4_in[446]),
   .I3(level4_in[447]),
   .I4(level4_in[448]),
   .I5(level4_in[449])
);

LUT6 #(
   .INIT(64'h8f39f1218f39f121)  
) LUT6_inst7851 (
   .O(to_level3[75]),
   .I0(level4_in[450]),
   .I1(level4_in[451]),
   .I2(level4_in[452]),
   .I3(level4_in[453]),
   .I4(level4_in[454]),
   .I5(level4_in[455])
);

LUT6 #(
   .INIT(64'h419743f6419743f6)  
) LUT6_inst7852 (
   .O(to_level3[76]),
   .I0(level4_in[456]),
   .I1(level4_in[457]),
   .I2(level4_in[458]),
   .I3(level4_in[459]),
   .I4(level4_in[460]),
   .I5(level4_in[461])
);

LUT6 #(
   .INIT(64'hd4fa855bd4fa855b)  
) LUT6_inst7853 (
   .O(to_level3[77]),
   .I0(level4_in[462]),
   .I1(level4_in[463]),
   .I2(level4_in[464]),
   .I3(level4_in[465]),
   .I4(level4_in[466]),
   .I5(level4_in[467])
);

LUT6 #(
   .INIT(64'h96e3d84696e3d846)  
) LUT6_inst7854 (
   .O(to_level3[78]),
   .I0(level4_in[468]),
   .I1(level4_in[469]),
   .I2(level4_in[470]),
   .I3(level4_in[471]),
   .I4(level4_in[472]),
   .I5(level4_in[473])
);

LUT6 #(
   .INIT(64'h032671a8032671a8)  
) LUT6_inst7855 (
   .O(to_level3[79]),
   .I0(level4_in[474]),
   .I1(level4_in[475]),
   .I2(level4_in[476]),
   .I3(level4_in[477]),
   .I4(level4_in[478]),
   .I5(level4_in[479])
);

LUT6 #(
   .INIT(64'h2c1e5f982c1e5f98)  
) LUT6_inst7856 (
   .O(to_level3[80]),
   .I0(level4_in[480]),
   .I1(level4_in[481]),
   .I2(level4_in[482]),
   .I3(level4_in[483]),
   .I4(level4_in[484]),
   .I5(level4_in[485])
);

LUT6 #(
   .INIT(64'h1a0c6ec11a0c6ec1)  
) LUT6_inst7857 (
   .O(to_level3[81]),
   .I0(level4_in[486]),
   .I1(level4_in[487]),
   .I2(level4_in[488]),
   .I3(level4_in[489]),
   .I4(level4_in[490]),
   .I5(level4_in[491])
);

LUT6 #(
   .INIT(64'h4992024549920245)  
) LUT6_inst7858 (
   .O(to_level3[82]),
   .I0(level4_in[492]),
   .I1(level4_in[493]),
   .I2(level4_in[494]),
   .I3(level4_in[495]),
   .I4(level4_in[496]),
   .I5(level4_in[497])
);

LUT6 #(
   .INIT(64'h9e1915f59e1915f5)  
) LUT6_inst7859 (
   .O(to_level3[83]),
   .I0(level4_in[498]),
   .I1(level4_in[499]),
   .I2(level4_in[500]),
   .I3(level4_in[501]),
   .I4(level4_in[502]),
   .I5(level4_in[503])
);

LUT6 #(
   .INIT(64'h081f7bbf081f7bbf)  
) LUT6_inst7860 (
   .O(to_level3[84]),
   .I0(level4_in[504]),
   .I1(level4_in[505]),
   .I2(level4_in[506]),
   .I3(level4_in[507]),
   .I4(level4_in[508]),
   .I5(level4_in[509])
);

LUT6 #(
   .INIT(64'h86ed0c1b86ed0c1b)  
) LUT6_inst7861 (
   .O(to_level3[85]),
   .I0(level4_in[510]),
   .I1(level4_in[511]),
   .I2(level4_in[512]),
   .I3(level4_in[513]),
   .I4(level4_in[514]),
   .I5(level4_in[515])
);

LUT6 #(
   .INIT(64'h318bbab9318bbab9)  
) LUT6_inst7862 (
   .O(to_level3[86]),
   .I0(level4_in[516]),
   .I1(level4_in[517]),
   .I2(level4_in[518]),
   .I3(level4_in[519]),
   .I4(level4_in[520]),
   .I5(level4_in[521])
);

LUT6 #(
   .INIT(64'hd48de023d48de023)  
) LUT6_inst7863 (
   .O(to_level3[87]),
   .I0(level4_in[522]),
   .I1(level4_in[523]),
   .I2(level4_in[524]),
   .I3(level4_in[525]),
   .I4(level4_in[526]),
   .I5(level4_in[527])
);

LUT6 #(
   .INIT(64'h5728668157286681)  
) LUT6_inst7864 (
   .O(to_level3[88]),
   .I0(level4_in[528]),
   .I1(level4_in[529]),
   .I2(level4_in[530]),
   .I3(level4_in[531]),
   .I4(level4_in[532]),
   .I5(level4_in[533])
);

LUT6 #(
   .INIT(64'h4f414ced4f414ced)  
) LUT6_inst7865 (
   .O(to_level3[89]),
   .I0(level4_in[534]),
   .I1(level4_in[535]),
   .I2(level4_in[536]),
   .I3(level4_in[537]),
   .I4(level4_in[538]),
   .I5(level4_in[539])
);

LUT6 #(
   .INIT(64'heedcf1eaeedcf1ea)  
) LUT6_inst7866 (
   .O(to_level3[90]),
   .I0(level4_in[540]),
   .I1(level4_in[541]),
   .I2(level4_in[542]),
   .I3(level4_in[543]),
   .I4(level4_in[544]),
   .I5(level4_in[545])
);

LUT6 #(
   .INIT(64'ha05b6851a05b6851)  
) LUT6_inst7867 (
   .O(to_level3[91]),
   .I0(level4_in[546]),
   .I1(level4_in[547]),
   .I2(level4_in[548]),
   .I3(level4_in[549]),
   .I4(level4_in[550]),
   .I5(level4_in[551])
);

LUT6 #(
   .INIT(64'h8721924787219247)  
) LUT6_inst7868 (
   .O(to_level3[92]),
   .I0(level4_in[552]),
   .I1(level4_in[553]),
   .I2(level4_in[554]),
   .I3(level4_in[555]),
   .I4(level4_in[556]),
   .I5(level4_in[557])
);

LUT6 #(
   .INIT(64'hd8459ebfd8459ebf)  
) LUT6_inst7869 (
   .O(to_level3[93]),
   .I0(level4_in[558]),
   .I1(level4_in[559]),
   .I2(level4_in[560]),
   .I3(level4_in[561]),
   .I4(level4_in[562]),
   .I5(level4_in[563])
);

LUT6 #(
   .INIT(64'he93b85f4e93b85f4)  
) LUT6_inst7870 (
   .O(to_level3[94]),
   .I0(level4_in[564]),
   .I1(level4_in[565]),
   .I2(level4_in[566]),
   .I3(level4_in[567]),
   .I4(level4_in[568]),
   .I5(level4_in[569])
);

LUT6 #(
   .INIT(64'h09e8f6a209e8f6a2)  
) LUT6_inst7871 (
   .O(to_level3[95]),
   .I0(level4_in[570]),
   .I1(level4_in[571]),
   .I2(level4_in[572]),
   .I3(level4_in[573]),
   .I4(level4_in[574]),
   .I5(level4_in[575])
);

LUT6 #(
   .INIT(64'h3c520f203c520f20)  
) LUT6_inst7872 (
   .O(to_level3[96]),
   .I0(level4_in[576]),
   .I1(level4_in[577]),
   .I2(level4_in[578]),
   .I3(level4_in[579]),
   .I4(level4_in[580]),
   .I5(level4_in[581])
);

LUT6 #(
   .INIT(64'hb866001fb866001f)  
) LUT6_inst7873 (
   .O(to_level3[97]),
   .I0(level4_in[582]),
   .I1(level4_in[583]),
   .I2(level4_in[584]),
   .I3(level4_in[585]),
   .I4(level4_in[586]),
   .I5(level4_in[587])
);

LUT6 #(
   .INIT(64'hf3adc908f3adc908)  
) LUT6_inst7874 (
   .O(to_level3[98]),
   .I0(level4_in[588]),
   .I1(level4_in[589]),
   .I2(level4_in[590]),
   .I3(level4_in[591]),
   .I4(level4_in[592]),
   .I5(level4_in[593])
);

LUT6 #(
   .INIT(64'h0cc67fed0cc67fed)  
) LUT6_inst7875 (
   .O(to_level3[99]),
   .I0(level4_in[594]),
   .I1(level4_in[595]),
   .I2(level4_in[596]),
   .I3(level4_in[597]),
   .I4(level4_in[598]),
   .I5(level4_in[599])
);

LUT6 #(
   .INIT(64'h357d8d1f357d8d1f)  
) LUT6_inst7876 (
   .O(to_level3[100]),
   .I0(level4_in[600]),
   .I1(level4_in[601]),
   .I2(level4_in[602]),
   .I3(level4_in[603]),
   .I4(level4_in[604]),
   .I5(level4_in[605])
);

LUT6 #(
   .INIT(64'ha19c716fa19c716f)  
) LUT6_inst7877 (
   .O(to_level3[101]),
   .I0(level4_in[606]),
   .I1(level4_in[607]),
   .I2(level4_in[608]),
   .I3(level4_in[609]),
   .I4(level4_in[610]),
   .I5(level4_in[611])
);

LUT6 #(
   .INIT(64'hd864ce0bd864ce0b)  
) LUT6_inst7878 (
   .O(to_level3[102]),
   .I0(level4_in[612]),
   .I1(level4_in[613]),
   .I2(level4_in[614]),
   .I3(level4_in[615]),
   .I4(level4_in[616]),
   .I5(level4_in[617])
);

LUT6 #(
   .INIT(64'hfe439beffe439bef)  
) LUT6_inst7879 (
   .O(to_level3[103]),
   .I0(level4_in[618]),
   .I1(level4_in[619]),
   .I2(level4_in[620]),
   .I3(level4_in[621]),
   .I4(level4_in[622]),
   .I5(level4_in[623])
);

LUT6 #(
   .INIT(64'h78926f0b78926f0b)  
) LUT6_inst7880 (
   .O(to_level3[104]),
   .I0(level4_in[624]),
   .I1(level4_in[625]),
   .I2(level4_in[626]),
   .I3(level4_in[627]),
   .I4(level4_in[628]),
   .I5(level4_in[629])
);

LUT6 #(
   .INIT(64'h7f2a31d67f2a31d6)  
) LUT6_inst7881 (
   .O(to_level3[105]),
   .I0(level4_in[630]),
   .I1(level4_in[631]),
   .I2(level4_in[632]),
   .I3(level4_in[633]),
   .I4(level4_in[634]),
   .I5(level4_in[635])
);

LUT6 #(
   .INIT(64'hb76c35d5b76c35d5)  
) LUT6_inst7882 (
   .O(to_level3[106]),
   .I0(level4_in[636]),
   .I1(level4_in[637]),
   .I2(level4_in[638]),
   .I3(level4_in[639]),
   .I4(level4_in[640]),
   .I5(level4_in[641])
);

LUT6 #(
   .INIT(64'h5fca72885fca7288)  
) LUT6_inst7883 (
   .O(to_level3[107]),
   .I0(level4_in[642]),
   .I1(level4_in[643]),
   .I2(level4_in[644]),
   .I3(level4_in[645]),
   .I4(level4_in[646]),
   .I5(level4_in[647])
);

LUT6 #(
   .INIT(64'h232cc7ef232cc7ef)  
) LUT6_inst7884 (
   .O(to_level3[108]),
   .I0(level4_in[648]),
   .I1(level4_in[649]),
   .I2(level4_in[650]),
   .I3(level4_in[651]),
   .I4(level4_in[652]),
   .I5(level4_in[653])
);

LUT6 #(
   .INIT(64'h34d251ae34d251ae)  
) LUT6_inst7885 (
   .O(to_level3[109]),
   .I0(level4_in[654]),
   .I1(level4_in[655]),
   .I2(level4_in[656]),
   .I3(level4_in[657]),
   .I4(level4_in[658]),
   .I5(level4_in[659])
);

LUT6 #(
   .INIT(64'haed18157aed18157)  
) LUT6_inst7886 (
   .O(to_level3[110]),
   .I0(level4_in[660]),
   .I1(level4_in[661]),
   .I2(level4_in[662]),
   .I3(level4_in[663]),
   .I4(level4_in[664]),
   .I5(level4_in[665])
);

LUT6 #(
   .INIT(64'hb5420d4eb5420d4e)  
) LUT6_inst7887 (
   .O(to_level3[111]),
   .I0(level4_in[666]),
   .I1(level4_in[667]),
   .I2(level4_in[668]),
   .I3(level4_in[669]),
   .I4(level4_in[670]),
   .I5(level4_in[671])
);

LUT6 #(
   .INIT(64'h6d33384d6d33384d)  
) LUT6_inst7888 (
   .O(to_level3[112]),
   .I0(level4_in[672]),
   .I1(level4_in[673]),
   .I2(level4_in[674]),
   .I3(level4_in[675]),
   .I4(level4_in[676]),
   .I5(level4_in[677])
);

LUT6 #(
   .INIT(64'h0ab2b1e70ab2b1e7)  
) LUT6_inst7889 (
   .O(to_level3[113]),
   .I0(level4_in[678]),
   .I1(level4_in[679]),
   .I2(level4_in[680]),
   .I3(level4_in[681]),
   .I4(level4_in[682]),
   .I5(level4_in[683])
);

LUT6 #(
   .INIT(64'h1f48b6111f48b611)  
) LUT6_inst7890 (
   .O(to_level3[114]),
   .I0(level4_in[684]),
   .I1(level4_in[685]),
   .I2(level4_in[686]),
   .I3(level4_in[687]),
   .I4(level4_in[688]),
   .I5(level4_in[689])
);

LUT6 #(
   .INIT(64'hd02ee5bbd02ee5bb)  
) LUT6_inst7891 (
   .O(to_level3[115]),
   .I0(level4_in[690]),
   .I1(level4_in[691]),
   .I2(level4_in[692]),
   .I3(level4_in[693]),
   .I4(level4_in[694]),
   .I5(level4_in[695])
);

LUT6 #(
   .INIT(64'hc6fd24f9c6fd24f9)  
) LUT6_inst7892 (
   .O(to_level3[116]),
   .I0(level4_in[696]),
   .I1(level4_in[697]),
   .I2(level4_in[698]),
   .I3(level4_in[699]),
   .I4(level4_in[700]),
   .I5(level4_in[701])
);

LUT6 #(
   .INIT(64'h566292a6566292a6)  
) LUT6_inst7893 (
   .O(to_level3[117]),
   .I0(level4_in[702]),
   .I1(level4_in[703]),
   .I2(level4_in[704]),
   .I3(level4_in[705]),
   .I4(level4_in[706]),
   .I5(level4_in[707])
);

LUT6 #(
   .INIT(64'h76b456bc76b456bc)  
) LUT6_inst7894 (
   .O(to_level3[118]),
   .I0(level4_in[708]),
   .I1(level4_in[709]),
   .I2(level4_in[710]),
   .I3(level4_in[711]),
   .I4(level4_in[712]),
   .I5(level4_in[713])
);

LUT6 #(
   .INIT(64'ha71f446ca71f446c)  
) LUT6_inst7895 (
   .O(to_level3[119]),
   .I0(level4_in[714]),
   .I1(level4_in[715]),
   .I2(level4_in[716]),
   .I3(level4_in[717]),
   .I4(level4_in[718]),
   .I5(level4_in[719])
);

LUT6 #(
   .INIT(64'hc73b907dc73b907d)  
) LUT6_inst7896 (
   .O(to_level3[120]),
   .I0(level4_in[720]),
   .I1(level4_in[721]),
   .I2(level4_in[722]),
   .I3(level4_in[723]),
   .I4(level4_in[724]),
   .I5(level4_in[725])
);

LUT6 #(
   .INIT(64'h94da07c294da07c2)  
) LUT6_inst7897 (
   .O(to_level3[121]),
   .I0(level4_in[726]),
   .I1(level4_in[727]),
   .I2(level4_in[728]),
   .I3(level4_in[729]),
   .I4(level4_in[730]),
   .I5(level4_in[731])
);

LUT6 #(
   .INIT(64'h77a6e5d377a6e5d3)  
) LUT6_inst7898 (
   .O(to_level3[122]),
   .I0(level4_in[732]),
   .I1(level4_in[733]),
   .I2(level4_in[734]),
   .I3(level4_in[735]),
   .I4(level4_in[736]),
   .I5(level4_in[737])
);

LUT6 #(
   .INIT(64'h3c42f3953c42f395)  
) LUT6_inst7899 (
   .O(to_level3[123]),
   .I0(level4_in[738]),
   .I1(level4_in[739]),
   .I2(level4_in[740]),
   .I3(level4_in[741]),
   .I4(level4_in[742]),
   .I5(level4_in[743])
);

LUT6 #(
   .INIT(64'h3f0a2f353f0a2f35)  
) LUT6_inst7900 (
   .O(to_level3[124]),
   .I0(level4_in[744]),
   .I1(level4_in[745]),
   .I2(level4_in[746]),
   .I3(level4_in[747]),
   .I4(level4_in[748]),
   .I5(level4_in[749])
);

LUT6 #(
   .INIT(64'h795cd208795cd208)  
) LUT6_inst7901 (
   .O(to_level3[125]),
   .I0(level4_in[750]),
   .I1(level4_in[751]),
   .I2(level4_in[752]),
   .I3(level4_in[753]),
   .I4(level4_in[754]),
   .I5(level4_in[755])
);

LUT6 #(
   .INIT(64'hefe949c5efe949c5)  
) LUT6_inst7902 (
   .O(to_level3[126]),
   .I0(level4_in[756]),
   .I1(level4_in[757]),
   .I2(level4_in[758]),
   .I3(level4_in[759]),
   .I4(level4_in[760]),
   .I5(level4_in[761])
);

LUT6 #(
   .INIT(64'hb83f9d9cb83f9d9c)  
) LUT6_inst7903 (
   .O(to_level3[127]),
   .I0(level4_in[762]),
   .I1(level4_in[763]),
   .I2(level4_in[764]),
   .I3(level4_in[765]),
   .I4(level4_in[766]),
   .I5(level4_in[767])
);

LUT6 #(
   .INIT(64'he8f63796e8f63796)  
) LUT6_inst7904 (
   .O(to_level3[128]),
   .I0(level4_in[768]),
   .I1(level4_in[769]),
   .I2(level4_in[770]),
   .I3(level4_in[771]),
   .I4(level4_in[772]),
   .I5(level4_in[773])
);

LUT6 #(
   .INIT(64'hb2a8363ab2a8363a)  
) LUT6_inst7905 (
   .O(to_level3[129]),
   .I0(level4_in[774]),
   .I1(level4_in[775]),
   .I2(level4_in[776]),
   .I3(level4_in[777]),
   .I4(level4_in[778]),
   .I5(level4_in[779])
);

LUT6 #(
   .INIT(64'hc5b535d8c5b535d8)  
) LUT6_inst7906 (
   .O(to_level3[130]),
   .I0(level4_in[780]),
   .I1(level4_in[781]),
   .I2(level4_in[782]),
   .I3(level4_in[783]),
   .I4(level4_in[784]),
   .I5(level4_in[785])
);

LUT6 #(
   .INIT(64'habfc3e8eabfc3e8e)  
) LUT6_inst7907 (
   .O(to_level3[131]),
   .I0(level4_in[786]),
   .I1(level4_in[787]),
   .I2(level4_in[788]),
   .I3(level4_in[789]),
   .I4(level4_in[790]),
   .I5(level4_in[791])
);

LUT6 #(
   .INIT(64'he4f3bce5e4f3bce5)  
) LUT6_inst7908 (
   .O(to_level3[132]),
   .I0(level4_in[792]),
   .I1(level4_in[793]),
   .I2(level4_in[794]),
   .I3(level4_in[795]),
   .I4(level4_in[796]),
   .I5(level4_in[797])
);

LUT6 #(
   .INIT(64'h550a55ef550a55ef)  
) LUT6_inst7909 (
   .O(to_level3[133]),
   .I0(level4_in[798]),
   .I1(level4_in[799]),
   .I2(level4_in[800]),
   .I3(level4_in[801]),
   .I4(level4_in[802]),
   .I5(level4_in[803])
);

LUT6 #(
   .INIT(64'h34b0e05534b0e055)  
) LUT6_inst7910 (
   .O(to_level3[134]),
   .I0(level4_in[804]),
   .I1(level4_in[805]),
   .I2(level4_in[806]),
   .I3(level4_in[807]),
   .I4(level4_in[808]),
   .I5(level4_in[809])
);

LUT6 #(
   .INIT(64'h70ccd09a70ccd09a)  
) LUT6_inst7911 (
   .O(to_level3[135]),
   .I0(level4_in[810]),
   .I1(level4_in[811]),
   .I2(level4_in[812]),
   .I3(level4_in[813]),
   .I4(level4_in[814]),
   .I5(level4_in[815])
);

LUT6 #(
   .INIT(64'h7c57454e7c57454e)  
) LUT6_inst7912 (
   .O(to_level3[136]),
   .I0(level4_in[816]),
   .I1(level4_in[817]),
   .I2(level4_in[818]),
   .I3(level4_in[819]),
   .I4(level4_in[820]),
   .I5(level4_in[821])
);

LUT6 #(
   .INIT(64'h700ac4bf700ac4bf)  
) LUT6_inst7913 (
   .O(to_level3[137]),
   .I0(level4_in[822]),
   .I1(level4_in[823]),
   .I2(level4_in[824]),
   .I3(level4_in[825]),
   .I4(level4_in[826]),
   .I5(level4_in[827])
);

LUT6 #(
   .INIT(64'h65eb5f5965eb5f59)  
) LUT6_inst7914 (
   .O(to_level3[138]),
   .I0(level4_in[828]),
   .I1(level4_in[829]),
   .I2(level4_in[830]),
   .I3(level4_in[831]),
   .I4(level4_in[832]),
   .I5(level4_in[833])
);

LUT6 #(
   .INIT(64'hda8dd0a6da8dd0a6)  
) LUT6_inst7915 (
   .O(to_level3[139]),
   .I0(level4_in[834]),
   .I1(level4_in[835]),
   .I2(level4_in[836]),
   .I3(level4_in[837]),
   .I4(level4_in[838]),
   .I5(level4_in[839])
);

LUT6 #(
   .INIT(64'he4f137d0e4f137d0)  
) LUT6_inst7916 (
   .O(to_level3[140]),
   .I0(level4_in[840]),
   .I1(level4_in[841]),
   .I2(level4_in[842]),
   .I3(level4_in[843]),
   .I4(level4_in[844]),
   .I5(level4_in[845])
);

LUT6 #(
   .INIT(64'h4a8ed8fc4a8ed8fc)  
) LUT6_inst7917 (
   .O(to_level3[141]),
   .I0(level4_in[846]),
   .I1(level4_in[847]),
   .I2(level4_in[848]),
   .I3(level4_in[849]),
   .I4(level4_in[850]),
   .I5(level4_in[851])
);

LUT6 #(
   .INIT(64'he6d529e7e6d529e7)  
) LUT6_inst7918 (
   .O(to_level3[142]),
   .I0(level4_in[852]),
   .I1(level4_in[853]),
   .I2(level4_in[854]),
   .I3(level4_in[855]),
   .I4(level4_in[856]),
   .I5(level4_in[857])
);

LUT6 #(
   .INIT(64'hb36a7b9bb36a7b9b)  
) LUT6_inst7919 (
   .O(to_level3[143]),
   .I0(level4_in[858]),
   .I1(level4_in[859]),
   .I2(level4_in[860]),
   .I3(level4_in[861]),
   .I4(level4_in[862]),
   .I5(level4_in[863])
);

LUT6 #(
   .INIT(64'hc7dc7991c7dc7991)  
) LUT6_inst7920 (
   .O(to_level3[144]),
   .I0(level4_in[864]),
   .I1(level4_in[865]),
   .I2(level4_in[866]),
   .I3(level4_in[867]),
   .I4(level4_in[868]),
   .I5(level4_in[869])
);

LUT6 #(
   .INIT(64'h5206940752069407)  
) LUT6_inst7921 (
   .O(to_level3[145]),
   .I0(level4_in[870]),
   .I1(level4_in[871]),
   .I2(level4_in[872]),
   .I3(level4_in[873]),
   .I4(level4_in[874]),
   .I5(level4_in[875])
);

LUT6 #(
   .INIT(64'h3e48a4f43e48a4f4)  
) LUT6_inst7922 (
   .O(to_level3[146]),
   .I0(level4_in[876]),
   .I1(level4_in[877]),
   .I2(level4_in[878]),
   .I3(level4_in[879]),
   .I4(level4_in[880]),
   .I5(level4_in[881])
);

LUT6 #(
   .INIT(64'h0feb6d560feb6d56)  
) LUT6_inst7923 (
   .O(to_level3[147]),
   .I0(level4_in[882]),
   .I1(level4_in[883]),
   .I2(level4_in[884]),
   .I3(level4_in[885]),
   .I4(level4_in[886]),
   .I5(level4_in[887])
);

LUT6 #(
   .INIT(64'hb7a2a359b7a2a359)  
) LUT6_inst7924 (
   .O(to_level3[148]),
   .I0(level4_in[888]),
   .I1(level4_in[889]),
   .I2(level4_in[890]),
   .I3(level4_in[891]),
   .I4(level4_in[892]),
   .I5(level4_in[893])
);

LUT6 #(
   .INIT(64'h30409f3930409f39)  
) LUT6_inst7925 (
   .O(to_level3[149]),
   .I0(level4_in[894]),
   .I1(level4_in[895]),
   .I2(level4_in[896]),
   .I3(level4_in[897]),
   .I4(level4_in[898]),
   .I5(level4_in[899])
);

LUT6 #(
   .INIT(64'h2d9ab95d2d9ab95d)  
) LUT6_inst7926 (
   .O(to_level3[150]),
   .I0(level4_in[900]),
   .I1(level4_in[901]),
   .I2(level4_in[902]),
   .I3(level4_in[903]),
   .I4(level4_in[904]),
   .I5(level4_in[905])
);

LUT6 #(
   .INIT(64'h0924357909243579)  
) LUT6_inst7927 (
   .O(to_level3[151]),
   .I0(level4_in[906]),
   .I1(level4_in[907]),
   .I2(level4_in[908]),
   .I3(level4_in[909]),
   .I4(level4_in[910]),
   .I5(level4_in[911])
);

LUT6 #(
   .INIT(64'h9249fc059249fc05)  
) LUT6_inst7928 (
   .O(to_level3[152]),
   .I0(level4_in[912]),
   .I1(level4_in[913]),
   .I2(level4_in[914]),
   .I3(level4_in[915]),
   .I4(level4_in[916]),
   .I5(level4_in[917])
);

LUT6 #(
   .INIT(64'h94772daf94772daf)  
) LUT6_inst7929 (
   .O(to_level3[153]),
   .I0(level4_in[918]),
   .I1(level4_in[919]),
   .I2(level4_in[920]),
   .I3(level4_in[921]),
   .I4(level4_in[922]),
   .I5(level4_in[923])
);

LUT6 #(
   .INIT(64'hac60ffe0ac60ffe0)  
) LUT6_inst7930 (
   .O(to_level3[154]),
   .I0(level4_in[924]),
   .I1(level4_in[925]),
   .I2(level4_in[926]),
   .I3(level4_in[927]),
   .I4(level4_in[928]),
   .I5(level4_in[929])
);

LUT6 #(
   .INIT(64'hf86600acf86600ac)  
) LUT6_inst7931 (
   .O(to_level3[155]),
   .I0(level4_in[930]),
   .I1(level4_in[931]),
   .I2(level4_in[932]),
   .I3(level4_in[933]),
   .I4(level4_in[934]),
   .I5(level4_in[935])
);

LUT6 #(
   .INIT(64'h5c215c485c215c48)  
) LUT6_inst7932 (
   .O(to_level3[156]),
   .I0(level4_in[936]),
   .I1(level4_in[937]),
   .I2(level4_in[938]),
   .I3(level4_in[939]),
   .I4(level4_in[940]),
   .I5(level4_in[941])
);

LUT6 #(
   .INIT(64'h5733476957334769)  
) LUT6_inst7933 (
   .O(to_level3[157]),
   .I0(level4_in[942]),
   .I1(level4_in[943]),
   .I2(level4_in[944]),
   .I3(level4_in[945]),
   .I4(level4_in[946]),
   .I5(level4_in[947])
);

LUT6 #(
   .INIT(64'hbbca9f32bbca9f32)  
) LUT6_inst7934 (
   .O(to_level3[158]),
   .I0(level4_in[948]),
   .I1(level4_in[949]),
   .I2(level4_in[950]),
   .I3(level4_in[951]),
   .I4(level4_in[952]),
   .I5(level4_in[953])
);

LUT6 #(
   .INIT(64'h479e8c59479e8c59)  
) LUT6_inst7935 (
   .O(to_level3[159]),
   .I0(level4_in[954]),
   .I1(level4_in[955]),
   .I2(level4_in[956]),
   .I3(level4_in[957]),
   .I4(level4_in[958]),
   .I5(level4_in[959])
);

LUT6 #(
   .INIT(64'h221a5cb7221a5cb7)  
) LUT6_inst7936 (
   .O(to_level3[160]),
   .I0(level4_in[960]),
   .I1(level4_in[961]),
   .I2(level4_in[962]),
   .I3(level4_in[963]),
   .I4(level4_in[964]),
   .I5(level4_in[965])
);

LUT6 #(
   .INIT(64'haa95816caa95816c)  
) LUT6_inst7937 (
   .O(to_level3[161]),
   .I0(level4_in[966]),
   .I1(level4_in[967]),
   .I2(level4_in[968]),
   .I3(level4_in[969]),
   .I4(level4_in[970]),
   .I5(level4_in[971])
);

LUT6 #(
   .INIT(64'h843381dc843381dc)  
) LUT6_inst7938 (
   .O(to_level3[162]),
   .I0(level4_in[972]),
   .I1(level4_in[973]),
   .I2(level4_in[974]),
   .I3(level4_in[975]),
   .I4(level4_in[976]),
   .I5(level4_in[977])
);

LUT6 #(
   .INIT(64'hbcd64901bcd64901)  
) LUT6_inst7939 (
   .O(to_level3[163]),
   .I0(level4_in[978]),
   .I1(level4_in[979]),
   .I2(level4_in[980]),
   .I3(level4_in[981]),
   .I4(level4_in[982]),
   .I5(level4_in[983])
);

LUT6 #(
   .INIT(64'h5a4e36dd5a4e36dd)  
) LUT6_inst7940 (
   .O(to_level3[164]),
   .I0(level4_in[984]),
   .I1(level4_in[985]),
   .I2(level4_in[986]),
   .I3(level4_in[987]),
   .I4(level4_in[988]),
   .I5(level4_in[989])
);

LUT6 #(
   .INIT(64'h97ef349497ef3494)  
) LUT6_inst7941 (
   .O(to_level3[165]),
   .I0(level4_in[990]),
   .I1(level4_in[991]),
   .I2(level4_in[992]),
   .I3(level4_in[993]),
   .I4(level4_in[994]),
   .I5(level4_in[995])
);

LUT6 #(
   .INIT(64'h99a64f5a99a64f5a)  
) LUT6_inst7942 (
   .O(to_level3[166]),
   .I0(level4_in[996]),
   .I1(level4_in[997]),
   .I2(level4_in[998]),
   .I3(level4_in[999]),
   .I4(level4_in[1000]),
   .I5(level4_in[1001])
);

LUT6 #(
   .INIT(64'h05e4470705e44707)  
) LUT6_inst7943 (
   .O(to_level3[167]),
   .I0(level4_in[1002]),
   .I1(level4_in[1003]),
   .I2(level4_in[1004]),
   .I3(level4_in[1005]),
   .I4(level4_in[1006]),
   .I5(level4_in[1007])
);

LUT6 #(
   .INIT(64'h4134e22b4134e22b)  
) LUT6_inst7944 (
   .O(to_level3[168]),
   .I0(level4_in[1008]),
   .I1(level4_in[1009]),
   .I2(level4_in[1010]),
   .I3(level4_in[1011]),
   .I4(level4_in[1012]),
   .I5(level4_in[1013])
);

LUT6 #(
   .INIT(64'ha10c38aea10c38ae)  
) LUT6_inst7945 (
   .O(to_level3[169]),
   .I0(level4_in[1014]),
   .I1(level4_in[1015]),
   .I2(level4_in[1016]),
   .I3(level4_in[1017]),
   .I4(level4_in[1018]),
   .I5(level4_in[1019])
);

LUT6 #(
   .INIT(64'h545713fe545713fe)  
) LUT6_inst7946 (
   .O(to_level3[170]),
   .I0(level4_in[1020]),
   .I1(level4_in[1021]),
   .I2(level4_in[1022]),
   .I3(level4_in[1023]),
   .I4(level4_in[1024]),
   .I5(level4_in[1025])
);

LUT6 #(
   .INIT(64'h18aa559518aa5595)  
) LUT6_inst7947 (
   .O(to_level3[171]),
   .I0(level4_in[1026]),
   .I1(level4_in[1027]),
   .I2(level4_in[1028]),
   .I3(level4_in[1029]),
   .I4(level4_in[1030]),
   .I5(level4_in[1031])
);

LUT6 #(
   .INIT(64'haf00dcf3af00dcf3)  
) LUT6_inst7948 (
   .O(to_level3[172]),
   .I0(level4_in[1032]),
   .I1(level4_in[1033]),
   .I2(level4_in[1034]),
   .I3(level4_in[1035]),
   .I4(level4_in[1036]),
   .I5(level4_in[1037])
);

LUT6 #(
   .INIT(64'h4136146e4136146e)  
) LUT6_inst7949 (
   .O(to_level3[173]),
   .I0(level4_in[1038]),
   .I1(level4_in[1039]),
   .I2(level4_in[1040]),
   .I3(level4_in[1041]),
   .I4(level4_in[1042]),
   .I5(level4_in[1043])
);

LUT6 #(
   .INIT(64'h780ad82f780ad82f)  
) LUT6_inst7950 (
   .O(to_level3[174]),
   .I0(level4_in[1044]),
   .I1(level4_in[1045]),
   .I2(level4_in[1046]),
   .I3(level4_in[1047]),
   .I4(level4_in[1048]),
   .I5(level4_in[1049])
);

LUT6 #(
   .INIT(64'h2698c5d72698c5d7)  
) LUT6_inst7951 (
   .O(to_level3[175]),
   .I0(level4_in[1050]),
   .I1(level4_in[1051]),
   .I2(level4_in[1052]),
   .I3(level4_in[1053]),
   .I4(level4_in[1054]),
   .I5(level4_in[1055])
);

LUT6 #(
   .INIT(64'h33033d8e33033d8e)  
) LUT6_inst7952 (
   .O(to_level3[176]),
   .I0(level4_in[1056]),
   .I1(level4_in[1057]),
   .I2(level4_in[1058]),
   .I3(level4_in[1059]),
   .I4(level4_in[1060]),
   .I5(level4_in[1061])
);

LUT6 #(
   .INIT(64'h2c02124a2c02124a)  
) LUT6_inst7953 (
   .O(to_level3[177]),
   .I0(level4_in[1062]),
   .I1(level4_in[1063]),
   .I2(level4_in[1064]),
   .I3(level4_in[1065]),
   .I4(level4_in[1066]),
   .I5(level4_in[1067])
);

LUT6 #(
   .INIT(64'hd0cb1807d0cb1807)  
) LUT6_inst7954 (
   .O(to_level3[178]),
   .I0(level4_in[1068]),
   .I1(level4_in[1069]),
   .I2(level4_in[1070]),
   .I3(level4_in[1071]),
   .I4(level4_in[1072]),
   .I5(level4_in[1073])
);

LUT6 #(
   .INIT(64'h5489c7c05489c7c0)  
) LUT6_inst7955 (
   .O(to_level3[179]),
   .I0(level4_in[1074]),
   .I1(level4_in[1075]),
   .I2(level4_in[1076]),
   .I3(level4_in[1077]),
   .I4(level4_in[1078]),
   .I5(level4_in[1079])
);

LUT6 #(
   .INIT(64'he419f2e9e419f2e9)  
) LUT6_inst7956 (
   .O(to_level3[180]),
   .I0(level4_in[1080]),
   .I1(level4_in[1081]),
   .I2(level4_in[1082]),
   .I3(level4_in[1083]),
   .I4(level4_in[1084]),
   .I5(level4_in[1085])
);

LUT6 #(
   .INIT(64'h2da11bff2da11bff)  
) LUT6_inst7957 (
   .O(to_level3[181]),
   .I0(level4_in[1086]),
   .I1(level4_in[1087]),
   .I2(level4_in[1088]),
   .I3(level4_in[1089]),
   .I4(level4_in[1090]),
   .I5(level4_in[1091])
);

LUT6 #(
   .INIT(64'h8127eeb58127eeb5)  
) LUT6_inst7958 (
   .O(to_level3[182]),
   .I0(level4_in[1092]),
   .I1(level4_in[1093]),
   .I2(level4_in[1094]),
   .I3(level4_in[1095]),
   .I4(level4_in[1096]),
   .I5(level4_in[1097])
);

LUT6 #(
   .INIT(64'h14c6ec6514c6ec65)  
) LUT6_inst7959 (
   .O(to_level3[183]),
   .I0(level4_in[1098]),
   .I1(level4_in[1099]),
   .I2(level4_in[1100]),
   .I3(level4_in[1101]),
   .I4(level4_in[1102]),
   .I5(level4_in[1103])
);

LUT6 #(
   .INIT(64'hc37b8545c37b8545)  
) LUT6_inst7960 (
   .O(to_level3[184]),
   .I0(level4_in[1104]),
   .I1(level4_in[1105]),
   .I2(level4_in[1106]),
   .I3(level4_in[1107]),
   .I4(level4_in[1108]),
   .I5(level4_in[1109])
);

LUT6 #(
   .INIT(64'h4863b9be4863b9be)  
) LUT6_inst7961 (
   .O(to_level3[185]),
   .I0(level4_in[1110]),
   .I1(level4_in[1111]),
   .I2(level4_in[1112]),
   .I3(level4_in[1113]),
   .I4(level4_in[1114]),
   .I5(level4_in[1115])
);

LUT6 #(
   .INIT(64'h9714382c9714382c)  
) LUT6_inst7962 (
   .O(to_level3[186]),
   .I0(level4_in[1116]),
   .I1(level4_in[1117]),
   .I2(level4_in[1118]),
   .I3(level4_in[1119]),
   .I4(level4_in[1120]),
   .I5(level4_in[1121])
);

LUT6 #(
   .INIT(64'h0df3b8910df3b891)  
) LUT6_inst7963 (
   .O(to_level3[187]),
   .I0(level4_in[1122]),
   .I1(level4_in[1123]),
   .I2(level4_in[1124]),
   .I3(level4_in[1125]),
   .I4(level4_in[1126]),
   .I5(level4_in[1127])
);

LUT6 #(
   .INIT(64'h08b0238908b02389)  
) LUT6_inst7964 (
   .O(to_level3[188]),
   .I0(level4_in[1128]),
   .I1(level4_in[1129]),
   .I2(level4_in[1130]),
   .I3(level4_in[1131]),
   .I4(level4_in[1132]),
   .I5(level4_in[1133])
);

LUT6 #(
   .INIT(64'hab2315eaab2315ea)  
) LUT6_inst7965 (
   .O(to_level3[189]),
   .I0(level4_in[1134]),
   .I1(level4_in[1135]),
   .I2(level4_in[1136]),
   .I3(level4_in[1137]),
   .I4(level4_in[1138]),
   .I5(level4_in[1139])
);

LUT6 #(
   .INIT(64'h56d8715556d87155)  
) LUT6_inst7966 (
   .O(to_level3[190]),
   .I0(level4_in[1140]),
   .I1(level4_in[1141]),
   .I2(level4_in[1142]),
   .I3(level4_in[1143]),
   .I4(level4_in[1144]),
   .I5(level4_in[1145])
);

LUT6 #(
   .INIT(64'hd0111c04d0111c04)  
) LUT6_inst7967 (
   .O(to_level3[191]),
   .I0(level4_in[1146]),
   .I1(level4_in[1147]),
   .I2(level4_in[1148]),
   .I3(level4_in[1149]),
   .I4(level4_in[1150]),
   .I5(level4_in[1151])
);

LUT6 #(
   .INIT(64'h14ea898e14ea898e)  
) LUT6_inst7968 (
   .O(to_level3[192]),
   .I0(level4_in[1152]),
   .I1(level4_in[1153]),
   .I2(level4_in[1154]),
   .I3(level4_in[1155]),
   .I4(level4_in[1156]),
   .I5(level4_in[1157])
);

LUT6 #(
   .INIT(64'h99370ccf99370ccf)  
) LUT6_inst7969 (
   .O(to_level3[193]),
   .I0(level4_in[1158]),
   .I1(level4_in[1159]),
   .I2(level4_in[1160]),
   .I3(level4_in[1161]),
   .I4(level4_in[1162]),
   .I5(level4_in[1163])
);

LUT6 #(
   .INIT(64'h5c32c61d5c32c61d)  
) LUT6_inst7970 (
   .O(to_level3[194]),
   .I0(level4_in[1164]),
   .I1(level4_in[1165]),
   .I2(level4_in[1166]),
   .I3(level4_in[1167]),
   .I4(level4_in[1168]),
   .I5(level4_in[1169])
);

LUT6 #(
   .INIT(64'h78bfbb8178bfbb81)  
) LUT6_inst7971 (
   .O(to_level3[195]),
   .I0(level4_in[1170]),
   .I1(level4_in[1171]),
   .I2(level4_in[1172]),
   .I3(level4_in[1173]),
   .I4(level4_in[1174]),
   .I5(level4_in[1175])
);

LUT6 #(
   .INIT(64'h9077341390773413)  
) LUT6_inst7972 (
   .O(to_level3[196]),
   .I0(level4_in[1176]),
   .I1(level4_in[1177]),
   .I2(level4_in[1178]),
   .I3(level4_in[1179]),
   .I4(level4_in[1180]),
   .I5(level4_in[1181])
);

LUT6 #(
   .INIT(64'h9243286992432869)  
) LUT6_inst7973 (
   .O(to_level3[197]),
   .I0(level4_in[1182]),
   .I1(level4_in[1183]),
   .I2(level4_in[1184]),
   .I3(level4_in[1185]),
   .I4(level4_in[1186]),
   .I5(level4_in[1187])
);

LUT6 #(
   .INIT(64'h2f6005042f600504)  
) LUT6_inst7974 (
   .O(to_level3[198]),
   .I0(level4_in[1188]),
   .I1(level4_in[1189]),
   .I2(level4_in[1190]),
   .I3(level4_in[1191]),
   .I4(level4_in[1192]),
   .I5(level4_in[1193])
);

LUT6 #(
   .INIT(64'he7950980e7950980)  
) LUT6_inst7975 (
   .O(to_level3[199]),
   .I0(level4_in[1194]),
   .I1(level4_in[1195]),
   .I2(level4_in[1196]),
   .I3(level4_in[1197]),
   .I4(level4_in[1198]),
   .I5(level4_in[1199])
);

LUT6 #(
   .INIT(64'h104341dc104341dc)  
) LUT6_inst7976 (
   .O(to_level3[200]),
   .I0(level4_in[1200]),
   .I1(level4_in[1201]),
   .I2(level4_in[1202]),
   .I3(level4_in[1203]),
   .I4(level4_in[1204]),
   .I5(level4_in[1205])
);

LUT6 #(
   .INIT(64'h2b5995dc2b5995dc)  
) LUT6_inst7977 (
   .O(to_level3[201]),
   .I0(level4_in[1206]),
   .I1(level4_in[1207]),
   .I2(level4_in[1208]),
   .I3(level4_in[1209]),
   .I4(level4_in[1210]),
   .I5(level4_in[1211])
);

LUT6 #(
   .INIT(64'h8edbace08edbace0)  
) LUT6_inst7978 (
   .O(to_level3[202]),
   .I0(level4_in[1212]),
   .I1(level4_in[1213]),
   .I2(level4_in[1214]),
   .I3(level4_in[1215]),
   .I4(level4_in[1216]),
   .I5(level4_in[1217])
);

LUT6 #(
   .INIT(64'h462cfb9f462cfb9f)  
) LUT6_inst7979 (
   .O(to_level3[203]),
   .I0(level4_in[1218]),
   .I1(level4_in[1219]),
   .I2(level4_in[1220]),
   .I3(level4_in[1221]),
   .I4(level4_in[1222]),
   .I5(level4_in[1223])
);

LUT6 #(
   .INIT(64'h9e85af619e85af61)  
) LUT6_inst7980 (
   .O(to_level3[204]),
   .I0(level4_in[1224]),
   .I1(level4_in[1225]),
   .I2(level4_in[1226]),
   .I3(level4_in[1227]),
   .I4(level4_in[1228]),
   .I5(level4_in[1229])
);

LUT6 #(
   .INIT(64'h34e4200e34e4200e)  
) LUT6_inst7981 (
   .O(to_level3[205]),
   .I0(level4_in[1230]),
   .I1(level4_in[1231]),
   .I2(level4_in[1232]),
   .I3(level4_in[1233]),
   .I4(level4_in[1234]),
   .I5(level4_in[1235])
);

LUT6 #(
   .INIT(64'h7e88b84b7e88b84b)  
) LUT6_inst7982 (
   .O(to_level3[206]),
   .I0(level4_in[1236]),
   .I1(level4_in[1237]),
   .I2(level4_in[1238]),
   .I3(level4_in[1239]),
   .I4(level4_in[1240]),
   .I5(level4_in[1241])
);

LUT6 #(
   .INIT(64'h18f6350e18f6350e)  
) LUT6_inst7983 (
   .O(to_level3[207]),
   .I0(level4_in[1242]),
   .I1(level4_in[1243]),
   .I2(level4_in[1244]),
   .I3(level4_in[1245]),
   .I4(level4_in[1246]),
   .I5(level4_in[1247])
);

LUT6 #(
   .INIT(64'hfcf29d4dfcf29d4d)  
) LUT6_inst7984 (
   .O(to_level3[208]),
   .I0(level4_in[1248]),
   .I1(level4_in[1249]),
   .I2(level4_in[1250]),
   .I3(level4_in[1251]),
   .I4(level4_in[1252]),
   .I5(level4_in[1253])
);

LUT6 #(
   .INIT(64'h93ef55da93ef55da)  
) LUT6_inst7985 (
   .O(to_level3[209]),
   .I0(level4_in[1254]),
   .I1(level4_in[1255]),
   .I2(level4_in[1256]),
   .I3(level4_in[1257]),
   .I4(level4_in[1258]),
   .I5(level4_in[1259])
);

LUT6 #(
   .INIT(64'h11dc1a7411dc1a74)  
) LUT6_inst7986 (
   .O(to_level3[210]),
   .I0(level4_in[1260]),
   .I1(level4_in[1261]),
   .I2(level4_in[1262]),
   .I3(level4_in[1263]),
   .I4(level4_in[1264]),
   .I5(level4_in[1265])
);

LUT6 #(
   .INIT(64'hca121b43ca121b43)  
) LUT6_inst7987 (
   .O(to_level3[211]),
   .I0(level4_in[1266]),
   .I1(level4_in[1267]),
   .I2(level4_in[1268]),
   .I3(level4_in[1269]),
   .I4(level4_in[1270]),
   .I5(level4_in[1271])
);

LUT6 #(
   .INIT(64'h879b5ad3879b5ad3)  
) LUT6_inst7988 (
   .O(to_level3[212]),
   .I0(level4_in[1272]),
   .I1(level4_in[1273]),
   .I2(level4_in[1274]),
   .I3(level4_in[1275]),
   .I4(level4_in[1276]),
   .I5(level4_in[1277])
);

LUT6 #(
   .INIT(64'h689051f2689051f2)  
) LUT6_inst7989 (
   .O(to_level3[213]),
   .I0(level4_in[1278]),
   .I1(level4_in[1279]),
   .I2(level4_in[1280]),
   .I3(level4_in[1281]),
   .I4(level4_in[1282]),
   .I5(level4_in[1283])
);

LUT6 #(
   .INIT(64'h9c9410ee9c9410ee)  
) LUT6_inst7990 (
   .O(to_level3[214]),
   .I0(level4_in[1284]),
   .I1(level4_in[1285]),
   .I2(level4_in[1286]),
   .I3(level4_in[1287]),
   .I4(level4_in[1288]),
   .I5(level4_in[1289])
);

LUT6 #(
   .INIT(64'h002e8469002e8469)  
) LUT6_inst7991 (
   .O(to_level3[215]),
   .I0(level4_in[1290]),
   .I1(level4_in[1291]),
   .I2(level4_in[1292]),
   .I3(level4_in[1293]),
   .I4(level4_in[1294]),
   .I5(level4_in[1295])
);

LUT6 #(
   .INIT(64'h73dc956673dc9566)  
) LUT6_inst7992 (
   .O(to_level3[216]),
   .I0(level4_in[1296]),
   .I1(level4_in[1297]),
   .I2(level4_in[1298]),
   .I3(level4_in[1299]),
   .I4(level4_in[1300]),
   .I5(level4_in[1301])
);

LUT6 #(
   .INIT(64'heba7c318eba7c318)  
) LUT6_inst7993 (
   .O(to_level3[217]),
   .I0(level4_in[1302]),
   .I1(level4_in[1303]),
   .I2(level4_in[1304]),
   .I3(level4_in[1305]),
   .I4(level4_in[1306]),
   .I5(level4_in[1307])
);

LUT6 #(
   .INIT(64'h52eddbc152eddbc1)  
) LUT6_inst7994 (
   .O(to_level3[218]),
   .I0(level4_in[1308]),
   .I1(level4_in[1309]),
   .I2(level4_in[1310]),
   .I3(level4_in[1311]),
   .I4(level4_in[1312]),
   .I5(level4_in[1313])
);

LUT6 #(
   .INIT(64'h95f1269d95f1269d)  
) LUT6_inst7995 (
   .O(to_level3[219]),
   .I0(level4_in[1314]),
   .I1(level4_in[1315]),
   .I2(level4_in[1316]),
   .I3(level4_in[1317]),
   .I4(level4_in[1318]),
   .I5(level4_in[1319])
);

LUT6 #(
   .INIT(64'h6cb1be226cb1be22)  
) LUT6_inst7996 (
   .O(to_level3[220]),
   .I0(level4_in[1320]),
   .I1(level4_in[1321]),
   .I2(level4_in[1322]),
   .I3(level4_in[1323]),
   .I4(level4_in[1324]),
   .I5(level4_in[1325])
);

LUT6 #(
   .INIT(64'h8e3648c78e3648c7)  
) LUT6_inst7997 (
   .O(to_level3[221]),
   .I0(level4_in[1326]),
   .I1(level4_in[1327]),
   .I2(level4_in[1328]),
   .I3(level4_in[1329]),
   .I4(level4_in[1330]),
   .I5(level4_in[1331])
);

LUT6 #(
   .INIT(64'h0a5e1a680a5e1a68)  
) LUT6_inst7998 (
   .O(to_level3[222]),
   .I0(level4_in[1332]),
   .I1(level4_in[1333]),
   .I2(level4_in[1334]),
   .I3(level4_in[1335]),
   .I4(level4_in[1336]),
   .I5(level4_in[1337])
);

LUT6 #(
   .INIT(64'h8fd136d58fd136d5)  
) LUT6_inst7999 (
   .O(to_level3[223]),
   .I0(level4_in[1338]),
   .I1(level4_in[1339]),
   .I2(level4_in[1340]),
   .I3(level4_in[1341]),
   .I4(level4_in[1342]),
   .I5(level4_in[1343])
);

LUT6 #(
   .INIT(64'he77fd744e77fd744)  
) LUT6_inst8000 (
   .O(to_level3[224]),
   .I0(level4_in[1344]),
   .I1(level4_in[1345]),
   .I2(level4_in[1346]),
   .I3(level4_in[1347]),
   .I4(level4_in[1348]),
   .I5(level4_in[1349])
);

LUT6 #(
   .INIT(64'hcad7e17ccad7e17c)  
) LUT6_inst8001 (
   .O(to_level3[225]),
   .I0(level4_in[1350]),
   .I1(level4_in[1351]),
   .I2(level4_in[1352]),
   .I3(level4_in[1353]),
   .I4(level4_in[1354]),
   .I5(level4_in[1355])
);

LUT6 #(
   .INIT(64'h47ec30b547ec30b5)  
) LUT6_inst8002 (
   .O(to_level3[226]),
   .I0(level4_in[1356]),
   .I1(level4_in[1357]),
   .I2(level4_in[1358]),
   .I3(level4_in[1359]),
   .I4(level4_in[1360]),
   .I5(level4_in[1361])
);

LUT6 #(
   .INIT(64'hfb80bd06fb80bd06)  
) LUT6_inst8003 (
   .O(to_level3[227]),
   .I0(level4_in[1362]),
   .I1(level4_in[1363]),
   .I2(level4_in[1364]),
   .I3(level4_in[1365]),
   .I4(level4_in[1366]),
   .I5(level4_in[1367])
);

LUT6 #(
   .INIT(64'hd2b8b0b0d2b8b0b0)  
) LUT6_inst8004 (
   .O(to_level3[228]),
   .I0(level4_in[1368]),
   .I1(level4_in[1369]),
   .I2(level4_in[1370]),
   .I3(level4_in[1371]),
   .I4(level4_in[1372]),
   .I5(level4_in[1373])
);

LUT6 #(
   .INIT(64'h5f526b985f526b98)  
) LUT6_inst8005 (
   .O(to_level3[229]),
   .I0(level4_in[1374]),
   .I1(level4_in[1375]),
   .I2(level4_in[1376]),
   .I3(level4_in[1377]),
   .I4(level4_in[1378]),
   .I5(level4_in[1379])
);

LUT6 #(
   .INIT(64'hf1085dbcf1085dbc)  
) LUT6_inst8006 (
   .O(to_level3[230]),
   .I0(level4_in[1380]),
   .I1(level4_in[1381]),
   .I2(level4_in[1382]),
   .I3(level4_in[1383]),
   .I4(level4_in[1384]),
   .I5(level4_in[1385])
);

LUT6 #(
   .INIT(64'h202b311e202b311e)  
) LUT6_inst8007 (
   .O(to_level3[231]),
   .I0(level4_in[1386]),
   .I1(level4_in[1387]),
   .I2(level4_in[1388]),
   .I3(level4_in[1389]),
   .I4(level4_in[1390]),
   .I5(level4_in[1391])
);

LUT6 #(
   .INIT(64'h049dbc7c049dbc7c)  
) LUT6_inst8008 (
   .O(to_level3[232]),
   .I0(level4_in[1392]),
   .I1(level4_in[1393]),
   .I2(level4_in[1394]),
   .I3(level4_in[1395]),
   .I4(level4_in[1396]),
   .I5(level4_in[1397])
);

LUT6 #(
   .INIT(64'h3a1b27633a1b2763)  
) LUT6_inst8009 (
   .O(to_level3[233]),
   .I0(level4_in[1398]),
   .I1(level4_in[1399]),
   .I2(level4_in[1400]),
   .I3(level4_in[1401]),
   .I4(level4_in[1402]),
   .I5(level4_in[1403])
);

LUT6 #(
   .INIT(64'h3d7f13473d7f1347)  
) LUT6_inst8010 (
   .O(to_level3[234]),
   .I0(level4_in[1404]),
   .I1(level4_in[1405]),
   .I2(level4_in[1406]),
   .I3(level4_in[1407]),
   .I4(level4_in[1408]),
   .I5(level4_in[1409])
);

LUT6 #(
   .INIT(64'h8b3dfcad8b3dfcad)  
) LUT6_inst8011 (
   .O(to_level3[235]),
   .I0(level4_in[1410]),
   .I1(level4_in[1411]),
   .I2(level4_in[1412]),
   .I3(level4_in[1413]),
   .I4(level4_in[1414]),
   .I5(level4_in[1415])
);

LUT6 #(
   .INIT(64'hba98cc44ba98cc44)  
) LUT6_inst8012 (
   .O(to_level3[236]),
   .I0(level4_in[1416]),
   .I1(level4_in[1417]),
   .I2(level4_in[1418]),
   .I3(level4_in[1419]),
   .I4(level4_in[1420]),
   .I5(level4_in[1421])
);

LUT6 #(
   .INIT(64'h4bd355164bd35516)  
) LUT6_inst8013 (
   .O(to_level3[237]),
   .I0(level4_in[1422]),
   .I1(level4_in[1423]),
   .I2(level4_in[1424]),
   .I3(level4_in[1425]),
   .I4(level4_in[1426]),
   .I5(level4_in[1427])
);

LUT6 #(
   .INIT(64'h138ce544138ce544)  
) LUT6_inst8014 (
   .O(to_level3[238]),
   .I0(level4_in[1428]),
   .I1(level4_in[1429]),
   .I2(level4_in[1430]),
   .I3(level4_in[1431]),
   .I4(level4_in[1432]),
   .I5(level4_in[1433])
);

LUT6 #(
   .INIT(64'hc5aee568c5aee568)  
) LUT6_inst8015 (
   .O(to_level3[239]),
   .I0(level4_in[1434]),
   .I1(level4_in[1435]),
   .I2(level4_in[1436]),
   .I3(level4_in[1437]),
   .I4(level4_in[1438]),
   .I5(level4_in[1439])
);

LUT6 #(
   .INIT(64'h1da3b4091da3b409)  
) LUT6_inst8016 (
   .O(to_level3[240]),
   .I0(level4_in[1440]),
   .I1(level4_in[1441]),
   .I2(level4_in[1442]),
   .I3(level4_in[1443]),
   .I4(level4_in[1444]),
   .I5(level4_in[1445])
);

LUT6 #(
   .INIT(64'hcfb996b2cfb996b2)  
) LUT6_inst8017 (
   .O(to_level3[241]),
   .I0(level4_in[1446]),
   .I1(level4_in[1447]),
   .I2(level4_in[1448]),
   .I3(level4_in[1449]),
   .I4(level4_in[1450]),
   .I5(level4_in[1451])
);

LUT6 #(
   .INIT(64'h08a5b55608a5b556)  
) LUT6_inst8018 (
   .O(to_level3[242]),
   .I0(level4_in[1452]),
   .I1(level4_in[1453]),
   .I2(level4_in[1454]),
   .I3(level4_in[1455]),
   .I4(level4_in[1456]),
   .I5(level4_in[1457])
);

LUT6 #(
   .INIT(64'h9bc185e99bc185e9)  
) LUT6_inst8019 (
   .O(to_level3[243]),
   .I0(level4_in[1458]),
   .I1(level4_in[1459]),
   .I2(level4_in[1460]),
   .I3(level4_in[1461]),
   .I4(level4_in[1462]),
   .I5(level4_in[1463])
);

LUT6 #(
   .INIT(64'hab12d531ab12d531)  
) LUT6_inst8020 (
   .O(to_level3[244]),
   .I0(level4_in[1464]),
   .I1(level4_in[1465]),
   .I2(level4_in[1466]),
   .I3(level4_in[1467]),
   .I4(level4_in[1468]),
   .I5(level4_in[1469])
);

LUT6 #(
   .INIT(64'h0a455b5b0a455b5b)  
) LUT6_inst8021 (
   .O(to_level3[245]),
   .I0(level4_in[1470]),
   .I1(level4_in[1471]),
   .I2(level4_in[1472]),
   .I3(level4_in[1473]),
   .I4(level4_in[1474]),
   .I5(level4_in[1475])
);

LUT6 #(
   .INIT(64'h880d4803880d4803)  
) LUT6_inst8022 (
   .O(to_level3[246]),
   .I0(level4_in[1476]),
   .I1(level4_in[1477]),
   .I2(level4_in[1478]),
   .I3(level4_in[1479]),
   .I4(level4_in[1480]),
   .I5(level4_in[1481])
);

LUT6 #(
   .INIT(64'he867168fe867168f)  
) LUT6_inst8023 (
   .O(to_level3[247]),
   .I0(level4_in[1482]),
   .I1(level4_in[1483]),
   .I2(level4_in[1484]),
   .I3(level4_in[1485]),
   .I4(level4_in[1486]),
   .I5(level4_in[1487])
);

LUT6 #(
   .INIT(64'heda61573eda61573)  
) LUT6_inst8024 (
   .O(to_level3[248]),
   .I0(level4_in[1488]),
   .I1(level4_in[1489]),
   .I2(level4_in[1490]),
   .I3(level4_in[1491]),
   .I4(level4_in[1492]),
   .I5(level4_in[1493])
);

LUT6 #(
   .INIT(64'h976e96d9976e96d9)  
) LUT6_inst8025 (
   .O(to_level3[249]),
   .I0(level4_in[1494]),
   .I1(level4_in[1495]),
   .I2(level4_in[1496]),
   .I3(level4_in[1497]),
   .I4(level4_in[1498]),
   .I5(level4_in[1499])
);

LUT6 #(
   .INIT(64'h27f4e1e927f4e1e9)  
) LUT6_inst8026 (
   .O(to_level3[250]),
   .I0(level4_in[1500]),
   .I1(level4_in[1501]),
   .I2(level4_in[1502]),
   .I3(level4_in[1503]),
   .I4(level4_in[1504]),
   .I5(level4_in[1505])
);

LUT6 #(
   .INIT(64'hcaac73cbcaac73cb)  
) LUT6_inst8027 (
   .O(to_level3[251]),
   .I0(level4_in[1506]),
   .I1(level4_in[1507]),
   .I2(level4_in[1508]),
   .I3(level4_in[1509]),
   .I4(level4_in[1510]),
   .I5(level4_in[1511])
);

LUT6 #(
   .INIT(64'h936d374e936d374e)  
) LUT6_inst8028 (
   .O(to_level3[252]),
   .I0(level4_in[1512]),
   .I1(level4_in[1513]),
   .I2(level4_in[1514]),
   .I3(level4_in[1515]),
   .I4(level4_in[1516]),
   .I5(level4_in[1517])
);

LUT6 #(
   .INIT(64'h0c871a0a0c871a0a)  
) LUT6_inst8029 (
   .O(to_level3[253]),
   .I0(level4_in[1518]),
   .I1(level4_in[1519]),
   .I2(level4_in[1520]),
   .I3(level4_in[1521]),
   .I4(level4_in[1522]),
   .I5(level4_in[1523])
);

LUT6 #(
   .INIT(64'hd2559465d2559465)  
) LUT6_inst8030 (
   .O(to_level3[254]),
   .I0(level4_in[1524]),
   .I1(level4_in[1525]),
   .I2(level4_in[1526]),
   .I3(level4_in[1527]),
   .I4(level4_in[1528]),
   .I5(level4_in[1529])
);

LUT6 #(
   .INIT(64'h6b0826c66b0826c6)  
) LUT6_inst8031 (
   .O(to_level3[255]),
   .I0(level4_in[1530]),
   .I1(level4_in[1531]),
   .I2(level4_in[1532]),
   .I3(level4_in[1533]),
   .I4(level4_in[1534]),
   .I5(level4_in[1535])
);

LUT6 #(
   .INIT(64'hb7e28004b7e28004)  
) LUT6_inst8032 (
   .O(to_level3[256]),
   .I0(level4_in[1536]),
   .I1(level4_in[1537]),
   .I2(level4_in[1538]),
   .I3(level4_in[1539]),
   .I4(level4_in[1540]),
   .I5(level4_in[1541])
);

LUT6 #(
   .INIT(64'h356039ad356039ad)  
) LUT6_inst8033 (
   .O(to_level3[257]),
   .I0(level4_in[1542]),
   .I1(level4_in[1543]),
   .I2(level4_in[1544]),
   .I3(level4_in[1545]),
   .I4(level4_in[1546]),
   .I5(level4_in[1547])
);

LUT6 #(
   .INIT(64'h7e5ae7de7e5ae7de)  
) LUT6_inst8034 (
   .O(to_level3[258]),
   .I0(level4_in[1548]),
   .I1(level4_in[1549]),
   .I2(level4_in[1550]),
   .I3(level4_in[1551]),
   .I4(level4_in[1552]),
   .I5(level4_in[1553])
);

LUT6 #(
   .INIT(64'h4d9359cc4d9359cc)  
) LUT6_inst8035 (
   .O(to_level3[259]),
   .I0(level4_in[1554]),
   .I1(level4_in[1555]),
   .I2(level4_in[1556]),
   .I3(level4_in[1557]),
   .I4(level4_in[1558]),
   .I5(level4_in[1559])
);

LUT6 #(
   .INIT(64'h2a1bf6dd2a1bf6dd)  
) LUT6_inst8036 (
   .O(to_level3[260]),
   .I0(level4_in[1560]),
   .I1(level4_in[1561]),
   .I2(level4_in[1562]),
   .I3(level4_in[1563]),
   .I4(level4_in[1564]),
   .I5(level4_in[1565])
);

LUT6 #(
   .INIT(64'h1924f74b1924f74b)  
) LUT6_inst8037 (
   .O(to_level3[261]),
   .I0(level4_in[1566]),
   .I1(level4_in[1567]),
   .I2(level4_in[1568]),
   .I3(level4_in[1569]),
   .I4(level4_in[1570]),
   .I5(level4_in[1571])
);

LUT6 #(
   .INIT(64'h49b74f6c49b74f6c)  
) LUT6_inst8038 (
   .O(to_level3[262]),
   .I0(level4_in[1572]),
   .I1(level4_in[1573]),
   .I2(level4_in[1574]),
   .I3(level4_in[1575]),
   .I4(level4_in[1576]),
   .I5(level4_in[1577])
);

LUT6 #(
   .INIT(64'heaaef9dbeaaef9db)  
) LUT6_inst8039 (
   .O(to_level3[263]),
   .I0(level4_in[1578]),
   .I1(level4_in[1579]),
   .I2(level4_in[1580]),
   .I3(level4_in[1581]),
   .I4(level4_in[1582]),
   .I5(level4_in[1583])
);

LUT6 #(
   .INIT(64'h365c2d13365c2d13)  
) LUT6_inst8040 (
   .O(to_level3[264]),
   .I0(level4_in[1584]),
   .I1(level4_in[1585]),
   .I2(level4_in[1586]),
   .I3(level4_in[1587]),
   .I4(level4_in[1588]),
   .I5(level4_in[1589])
);

LUT6 #(
   .INIT(64'hc66cf77cc66cf77c)  
) LUT6_inst8041 (
   .O(to_level3[265]),
   .I0(level4_in[1590]),
   .I1(level4_in[1591]),
   .I2(level4_in[1592]),
   .I3(level4_in[1593]),
   .I4(level4_in[1594]),
   .I5(level4_in[1595])
);

LUT6 #(
   .INIT(64'h6a7e923e6a7e923e)  
) LUT6_inst8042 (
   .O(to_level3[266]),
   .I0(level4_in[1596]),
   .I1(level4_in[1597]),
   .I2(level4_in[1598]),
   .I3(level4_in[1599]),
   .I4(level4_in[1600]),
   .I5(level4_in[1601])
);

LUT6 #(
   .INIT(64'he3f861f9e3f861f9)  
) LUT6_inst8043 (
   .O(to_level3[267]),
   .I0(level4_in[1602]),
   .I1(level4_in[1603]),
   .I2(level4_in[1604]),
   .I3(level4_in[1605]),
   .I4(level4_in[1606]),
   .I5(level4_in[1607])
);

LUT6 #(
   .INIT(64'h4e646cb74e646cb7)  
) LUT6_inst8044 (
   .O(to_level3[268]),
   .I0(level4_in[1608]),
   .I1(level4_in[1609]),
   .I2(level4_in[1610]),
   .I3(level4_in[1611]),
   .I4(level4_in[1612]),
   .I5(level4_in[1613])
);

LUT6 #(
   .INIT(64'h821d9da1821d9da1)  
) LUT6_inst8045 (
   .O(to_level3[269]),
   .I0(level4_in[1614]),
   .I1(level4_in[1615]),
   .I2(level4_in[1616]),
   .I3(level4_in[1617]),
   .I4(level4_in[1618]),
   .I5(level4_in[1619])
);

LUT6 #(
   .INIT(64'h600e7754600e7754)  
) LUT6_inst8046 (
   .O(to_level3[270]),
   .I0(level4_in[1620]),
   .I1(level4_in[1621]),
   .I2(level4_in[1622]),
   .I3(level4_in[1623]),
   .I4(level4_in[1624]),
   .I5(level4_in[1625])
);

LUT6 #(
   .INIT(64'h34cbde0034cbde00)  
) LUT6_inst8047 (
   .O(to_level3[271]),
   .I0(level4_in[1626]),
   .I1(level4_in[1627]),
   .I2(level4_in[1628]),
   .I3(level4_in[1629]),
   .I4(level4_in[1630]),
   .I5(level4_in[1631])
);

LUT6 #(
   .INIT(64'hce60baccce60bacc)  
) LUT6_inst8048 (
   .O(to_level3[272]),
   .I0(level4_in[1632]),
   .I1(level4_in[1633]),
   .I2(level4_in[1634]),
   .I3(level4_in[1635]),
   .I4(level4_in[1636]),
   .I5(level4_in[1637])
);

LUT6 #(
   .INIT(64'hdca8c02cdca8c02c)  
) LUT6_inst8049 (
   .O(to_level3[273]),
   .I0(level4_in[1638]),
   .I1(level4_in[1639]),
   .I2(level4_in[1640]),
   .I3(level4_in[1641]),
   .I4(level4_in[1642]),
   .I5(level4_in[1643])
);

LUT6 #(
   .INIT(64'hd14f33c6d14f33c6)  
) LUT6_inst8050 (
   .O(to_level3[274]),
   .I0(level4_in[1644]),
   .I1(level4_in[1645]),
   .I2(level4_in[1646]),
   .I3(level4_in[1647]),
   .I4(level4_in[1648]),
   .I5(level4_in[1649])
);

LUT6 #(
   .INIT(64'hc1a02ecdc1a02ecd)  
) LUT6_inst8051 (
   .O(to_level3[275]),
   .I0(level4_in[1650]),
   .I1(level4_in[1651]),
   .I2(level4_in[1652]),
   .I3(level4_in[1653]),
   .I4(level4_in[1654]),
   .I5(level4_in[1655])
);

LUT6 #(
   .INIT(64'h78e89e2c78e89e2c)  
) LUT6_inst8052 (
   .O(to_level3[276]),
   .I0(level4_in[1656]),
   .I1(level4_in[1657]),
   .I2(level4_in[1658]),
   .I3(level4_in[1659]),
   .I4(level4_in[1660]),
   .I5(level4_in[1661])
);

LUT6 #(
   .INIT(64'h2ecb33462ecb3346)  
) LUT6_inst8053 (
   .O(to_level3[277]),
   .I0(level4_in[1662]),
   .I1(level4_in[1663]),
   .I2(level4_in[1664]),
   .I3(level4_in[1665]),
   .I4(level4_in[1666]),
   .I5(level4_in[1667])
);

LUT6 #(
   .INIT(64'h6f8ab04e6f8ab04e)  
) LUT6_inst8054 (
   .O(to_level3[278]),
   .I0(level4_in[1668]),
   .I1(level4_in[1669]),
   .I2(level4_in[1670]),
   .I3(level4_in[1671]),
   .I4(level4_in[1672]),
   .I5(level4_in[1673])
);

LUT6 #(
   .INIT(64'hd6abcdf1d6abcdf1)  
) LUT6_inst8055 (
   .O(to_level3[279]),
   .I0(level4_in[1674]),
   .I1(level4_in[1675]),
   .I2(level4_in[1676]),
   .I3(level4_in[1677]),
   .I4(level4_in[1678]),
   .I5(level4_in[1679])
);

LUT6 #(
   .INIT(64'h29e240b429e240b4)  
) LUT6_inst8056 (
   .O(to_level3[280]),
   .I0(level4_in[1680]),
   .I1(level4_in[1681]),
   .I2(level4_in[1682]),
   .I3(level4_in[1683]),
   .I4(level4_in[1684]),
   .I5(level4_in[1685])
);

LUT6 #(
   .INIT(64'h66c13d2a66c13d2a)  
) LUT6_inst8057 (
   .O(to_level3[281]),
   .I0(level4_in[1686]),
   .I1(level4_in[1687]),
   .I2(level4_in[1688]),
   .I3(level4_in[1689]),
   .I4(level4_in[1690]),
   .I5(level4_in[1691])
);

LUT6 #(
   .INIT(64'h105394ad105394ad)  
) LUT6_inst8058 (
   .O(to_level3[282]),
   .I0(level4_in[1692]),
   .I1(level4_in[1693]),
   .I2(level4_in[1694]),
   .I3(level4_in[1695]),
   .I4(level4_in[1696]),
   .I5(level4_in[1697])
);

LUT6 #(
   .INIT(64'ha70ccb35a70ccb35)  
) LUT6_inst8059 (
   .O(to_level3[283]),
   .I0(level4_in[1698]),
   .I1(level4_in[1699]),
   .I2(level4_in[1700]),
   .I3(level4_in[1701]),
   .I4(level4_in[1702]),
   .I5(level4_in[1703])
);

LUT6 #(
   .INIT(64'hc6d0c806c6d0c806)  
) LUT6_inst8060 (
   .O(to_level3[284]),
   .I0(level4_in[1704]),
   .I1(level4_in[1705]),
   .I2(level4_in[1706]),
   .I3(level4_in[1707]),
   .I4(level4_in[1708]),
   .I5(level4_in[1709])
);

LUT6 #(
   .INIT(64'h5d40a4db5d40a4db)  
) LUT6_inst8061 (
   .O(to_level3[285]),
   .I0(level4_in[1710]),
   .I1(level4_in[1711]),
   .I2(level4_in[1712]),
   .I3(level4_in[1713]),
   .I4(level4_in[1714]),
   .I5(level4_in[1715])
);

LUT6 #(
   .INIT(64'he7f80996e7f80996)  
) LUT6_inst8062 (
   .O(to_level3[286]),
   .I0(level4_in[1716]),
   .I1(level4_in[1717]),
   .I2(level4_in[1718]),
   .I3(level4_in[1719]),
   .I4(level4_in[1720]),
   .I5(level4_in[1721])
);

LUT6 #(
   .INIT(64'hb1b1f413b1b1f413)  
) LUT6_inst8063 (
   .O(to_level3[287]),
   .I0(level4_in[1722]),
   .I1(level4_in[1723]),
   .I2(level4_in[1724]),
   .I3(level4_in[1725]),
   .I4(level4_in[1726]),
   .I5(level4_in[1727])
);

LUT6 #(
   .INIT(64'h8c5f9fd88c5f9fd8)  
) LUT6_inst8064 (
   .O(to_level3[288]),
   .I0(level4_in[1728]),
   .I1(level4_in[1729]),
   .I2(level4_in[1730]),
   .I3(level4_in[1731]),
   .I4(level4_in[1732]),
   .I5(level4_in[1733])
);

LUT6 #(
   .INIT(64'h262c2f5d262c2f5d)  
) LUT6_inst8065 (
   .O(to_level3[289]),
   .I0(level4_in[1734]),
   .I1(level4_in[1735]),
   .I2(level4_in[1736]),
   .I3(level4_in[1737]),
   .I4(level4_in[1738]),
   .I5(level4_in[1739])
);

LUT6 #(
   .INIT(64'h1cb7f7931cb7f793)  
) LUT6_inst8066 (
   .O(to_level3[290]),
   .I0(level4_in[1740]),
   .I1(level4_in[1741]),
   .I2(level4_in[1742]),
   .I3(level4_in[1743]),
   .I4(level4_in[1744]),
   .I5(level4_in[1745])
);

LUT6 #(
   .INIT(64'ha9e3c9dba9e3c9db)  
) LUT6_inst8067 (
   .O(to_level3[291]),
   .I0(level4_in[1746]),
   .I1(level4_in[1747]),
   .I2(level4_in[1748]),
   .I3(level4_in[1749]),
   .I4(level4_in[1750]),
   .I5(level4_in[1751])
);

LUT6 #(
   .INIT(64'hb0cb0da5b0cb0da5)  
) LUT6_inst8068 (
   .O(to_level3[292]),
   .I0(level4_in[1752]),
   .I1(level4_in[1753]),
   .I2(level4_in[1754]),
   .I3(level4_in[1755]),
   .I4(level4_in[1756]),
   .I5(level4_in[1757])
);

LUT6 #(
   .INIT(64'he9e5057be9e5057b)  
) LUT6_inst8069 (
   .O(to_level3[293]),
   .I0(level4_in[1758]),
   .I1(level4_in[1759]),
   .I2(level4_in[1760]),
   .I3(level4_in[1761]),
   .I4(level4_in[1762]),
   .I5(level4_in[1763])
);

LUT6 #(
   .INIT(64'h1199f7301199f730)  
) LUT6_inst8070 (
   .O(to_level3[294]),
   .I0(level4_in[1764]),
   .I1(level4_in[1765]),
   .I2(level4_in[1766]),
   .I3(level4_in[1767]),
   .I4(level4_in[1768]),
   .I5(level4_in[1769])
);

LUT6 #(
   .INIT(64'h4f295af14f295af1)  
) LUT6_inst8071 (
   .O(to_level3[295]),
   .I0(level4_in[1770]),
   .I1(level4_in[1771]),
   .I2(level4_in[1772]),
   .I3(level4_in[1773]),
   .I4(level4_in[1774]),
   .I5(level4_in[1775])
);

LUT6 #(
   .INIT(64'hc0abddddc0abdddd)  
) LUT6_inst8072 (
   .O(to_level3[296]),
   .I0(level4_in[1776]),
   .I1(level4_in[1777]),
   .I2(level4_in[1778]),
   .I3(level4_in[1779]),
   .I4(level4_in[1780]),
   .I5(level4_in[1781])
);

LUT6 #(
   .INIT(64'h19672e1319672e13)  
) LUT6_inst8073 (
   .O(to_level3[297]),
   .I0(level4_in[1782]),
   .I1(level4_in[1783]),
   .I2(level4_in[1784]),
   .I3(level4_in[1785]),
   .I4(level4_in[1786]),
   .I5(level4_in[1787])
);

LUT6 #(
   .INIT(64'h51e334ce51e334ce)  
) LUT6_inst8074 (
   .O(to_level3[298]),
   .I0(level4_in[1788]),
   .I1(level4_in[1789]),
   .I2(level4_in[1790]),
   .I3(level4_in[1791]),
   .I4(level4_in[1792]),
   .I5(level4_in[1793])
);

LUT6 #(
   .INIT(64'h978565af978565af)  
) LUT6_inst8075 (
   .O(to_level3[299]),
   .I0(level4_in[1794]),
   .I1(level4_in[1795]),
   .I2(level4_in[1796]),
   .I3(level4_in[1797]),
   .I4(level4_in[1798]),
   .I5(level4_in[1799])
);

LUT6 #(
   .INIT(64'h44f3a9d344f3a9d3)  
) LUT6_inst8076 (
   .O(to_level3[300]),
   .I0(level4_in[1800]),
   .I1(level4_in[1801]),
   .I2(level4_in[1802]),
   .I3(level4_in[1803]),
   .I4(level4_in[1804]),
   .I5(level4_in[1805])
);

LUT6 #(
   .INIT(64'h21cc13c821cc13c8)  
) LUT6_inst8077 (
   .O(to_level3[301]),
   .I0(level4_in[1806]),
   .I1(level4_in[1807]),
   .I2(level4_in[1808]),
   .I3(level4_in[1809]),
   .I4(level4_in[1810]),
   .I5(level4_in[1811])
);

LUT6 #(
   .INIT(64'h8f4898958f489895)  
) LUT6_inst8078 (
   .O(to_level3[302]),
   .I0(level4_in[1812]),
   .I1(level4_in[1813]),
   .I2(level4_in[1814]),
   .I3(level4_in[1815]),
   .I4(level4_in[1816]),
   .I5(level4_in[1817])
);

LUT6 #(
   .INIT(64'h92865cf092865cf0)  
) LUT6_inst8079 (
   .O(to_level3[303]),
   .I0(level4_in[1818]),
   .I1(level4_in[1819]),
   .I2(level4_in[1820]),
   .I3(level4_in[1821]),
   .I4(level4_in[1822]),
   .I5(level4_in[1823])
);

LUT6 #(
   .INIT(64'h1a23abc01a23abc0)  
) LUT6_inst8080 (
   .O(to_level3[304]),
   .I0(level4_in[1824]),
   .I1(level4_in[1825]),
   .I2(level4_in[1826]),
   .I3(level4_in[1827]),
   .I4(level4_in[1828]),
   .I5(level4_in[1829])
);

LUT6 #(
   .INIT(64'hd3b72c31d3b72c31)  
) LUT6_inst8081 (
   .O(to_level3[305]),
   .I0(level4_in[1830]),
   .I1(level4_in[1831]),
   .I2(level4_in[1832]),
   .I3(level4_in[1833]),
   .I4(level4_in[1834]),
   .I5(level4_in[1835])
);

LUT6 #(
   .INIT(64'h96e5afee96e5afee)  
) LUT6_inst8082 (
   .O(to_level3[306]),
   .I0(level4_in[1836]),
   .I1(level4_in[1837]),
   .I2(level4_in[1838]),
   .I3(level4_in[1839]),
   .I4(level4_in[1840]),
   .I5(level4_in[1841])
);

LUT6 #(
   .INIT(64'h96e8201796e82017)  
) LUT6_inst8083 (
   .O(to_level3[307]),
   .I0(level4_in[1842]),
   .I1(level4_in[1843]),
   .I2(level4_in[1844]),
   .I3(level4_in[1845]),
   .I4(level4_in[1846]),
   .I5(level4_in[1847])
);

LUT6 #(
   .INIT(64'h1a08bfd01a08bfd0)  
) LUT6_inst8084 (
   .O(to_level3[308]),
   .I0(level4_in[1848]),
   .I1(level4_in[1849]),
   .I2(level4_in[1850]),
   .I3(level4_in[1851]),
   .I4(level4_in[1852]),
   .I5(level4_in[1853])
);

LUT6 #(
   .INIT(64'hfd4d32dbfd4d32db)  
) LUT6_inst8085 (
   .O(to_level3[309]),
   .I0(level4_in[1854]),
   .I1(level4_in[1855]),
   .I2(level4_in[1856]),
   .I3(level4_in[1857]),
   .I4(level4_in[1858]),
   .I5(level4_in[1859])
);

LUT6 #(
   .INIT(64'h6a4772b86a4772b8)  
) LUT6_inst8086 (
   .O(to_level3[310]),
   .I0(level4_in[1860]),
   .I1(level4_in[1861]),
   .I2(level4_in[1862]),
   .I3(level4_in[1863]),
   .I4(level4_in[1864]),
   .I5(level4_in[1865])
);

LUT6 #(
   .INIT(64'hf4f3a3daf4f3a3da)  
) LUT6_inst8087 (
   .O(to_level3[311]),
   .I0(level4_in[1866]),
   .I1(level4_in[1867]),
   .I2(level4_in[1868]),
   .I3(level4_in[1869]),
   .I4(level4_in[1870]),
   .I5(level4_in[1871])
);

LUT6 #(
   .INIT(64'h44cb411544cb4115)  
) LUT6_inst8088 (
   .O(to_level3[312]),
   .I0(level4_in[1872]),
   .I1(level4_in[1873]),
   .I2(level4_in[1874]),
   .I3(level4_in[1875]),
   .I4(level4_in[1876]),
   .I5(level4_in[1877])
);

LUT6 #(
   .INIT(64'h71eab02571eab025)  
) LUT6_inst8089 (
   .O(to_level3[313]),
   .I0(level4_in[1878]),
   .I1(level4_in[1879]),
   .I2(level4_in[1880]),
   .I3(level4_in[1881]),
   .I4(level4_in[1882]),
   .I5(level4_in[1883])
);

LUT6 #(
   .INIT(64'h4744ff184744ff18)  
) LUT6_inst8090 (
   .O(to_level3[314]),
   .I0(level4_in[1884]),
   .I1(level4_in[1885]),
   .I2(level4_in[1886]),
   .I3(level4_in[1887]),
   .I4(level4_in[1888]),
   .I5(level4_in[1889])
);

LUT6 #(
   .INIT(64'h555c3625555c3625)  
) LUT6_inst8091 (
   .O(to_level3[315]),
   .I0(level4_in[1890]),
   .I1(level4_in[1891]),
   .I2(level4_in[1892]),
   .I3(level4_in[1893]),
   .I4(level4_in[1894]),
   .I5(level4_in[1895])
);

LUT6 #(
   .INIT(64'h00127b8500127b85)  
) LUT6_inst8092 (
   .O(to_level3[316]),
   .I0(level4_in[1896]),
   .I1(level4_in[1897]),
   .I2(level4_in[1898]),
   .I3(level4_in[1899]),
   .I4(level4_in[1900]),
   .I5(level4_in[1901])
);

LUT6 #(
   .INIT(64'h9d7bf0669d7bf066)  
) LUT6_inst8093 (
   .O(to_level3[317]),
   .I0(level4_in[1902]),
   .I1(level4_in[1903]),
   .I2(level4_in[1904]),
   .I3(level4_in[1905]),
   .I4(level4_in[1906]),
   .I5(level4_in[1907])
);

LUT6 #(
   .INIT(64'h635092f6635092f6)  
) LUT6_inst8094 (
   .O(to_level3[318]),
   .I0(level4_in[1908]),
   .I1(level4_in[1909]),
   .I2(level4_in[1910]),
   .I3(level4_in[1911]),
   .I4(level4_in[1912]),
   .I5(level4_in[1913])
);

LUT6 #(
   .INIT(64'h7905ccc57905ccc5)  
) LUT6_inst8095 (
   .O(to_level3[319]),
   .I0(level4_in[1914]),
   .I1(level4_in[1915]),
   .I2(level4_in[1916]),
   .I3(level4_in[1917]),
   .I4(level4_in[1918]),
   .I5(level4_in[1919])
);

LUT6 #(
   .INIT(64'h91ff4dfa91ff4dfa)  
) LUT6_inst8096 (
   .O(to_level3[320]),
   .I0(level4_in[1920]),
   .I1(level4_in[1921]),
   .I2(level4_in[1922]),
   .I3(level4_in[1923]),
   .I4(level4_in[1924]),
   .I5(level4_in[1925])
);

LUT6 #(
   .INIT(64'h9625ccc69625ccc6)  
) LUT6_inst8097 (
   .O(to_level3[321]),
   .I0(level4_in[1926]),
   .I1(level4_in[1927]),
   .I2(level4_in[1928]),
   .I3(level4_in[1929]),
   .I4(level4_in[1930]),
   .I5(level4_in[1931])
);

LUT6 #(
   .INIT(64'h4a1d882d4a1d882d)  
) LUT6_inst8098 (
   .O(to_level3[322]),
   .I0(level4_in[1932]),
   .I1(level4_in[1933]),
   .I2(level4_in[1934]),
   .I3(level4_in[1935]),
   .I4(level4_in[1936]),
   .I5(level4_in[1937])
);

LUT6 #(
   .INIT(64'h299a286f299a286f)  
) LUT6_inst8099 (
   .O(to_level3[323]),
   .I0(level4_in[1938]),
   .I1(level4_in[1939]),
   .I2(level4_in[1940]),
   .I3(level4_in[1941]),
   .I4(level4_in[1942]),
   .I5(level4_in[1943])
);

LUT6 #(
   .INIT(64'hafe10133afe10133)  
) LUT6_inst8100 (
   .O(to_level3[324]),
   .I0(level4_in[1944]),
   .I1(level4_in[1945]),
   .I2(level4_in[1946]),
   .I3(level4_in[1947]),
   .I4(level4_in[1948]),
   .I5(level4_in[1949])
);

LUT6 #(
   .INIT(64'hfabea073fabea073)  
) LUT6_inst8101 (
   .O(to_level3[325]),
   .I0(level4_in[1950]),
   .I1(level4_in[1951]),
   .I2(level4_in[1952]),
   .I3(level4_in[1953]),
   .I4(level4_in[1954]),
   .I5(level4_in[1955])
);

LUT6 #(
   .INIT(64'h92c69e5092c69e50)  
) LUT6_inst8102 (
   .O(to_level3[326]),
   .I0(level4_in[1956]),
   .I1(level4_in[1957]),
   .I2(level4_in[1958]),
   .I3(level4_in[1959]),
   .I4(level4_in[1960]),
   .I5(level4_in[1961])
);

LUT6 #(
   .INIT(64'h79d59e9b79d59e9b)  
) LUT6_inst8103 (
   .O(to_level3[327]),
   .I0(level4_in[1962]),
   .I1(level4_in[1963]),
   .I2(level4_in[1964]),
   .I3(level4_in[1965]),
   .I4(level4_in[1966]),
   .I5(level4_in[1967])
);

LUT6 #(
   .INIT(64'hdda4d7f3dda4d7f3)  
) LUT6_inst8104 (
   .O(to_level3[328]),
   .I0(level4_in[1968]),
   .I1(level4_in[1969]),
   .I2(level4_in[1970]),
   .I3(level4_in[1971]),
   .I4(level4_in[1972]),
   .I5(level4_in[1973])
);

LUT6 #(
   .INIT(64'h3e25d8713e25d871)  
) LUT6_inst8105 (
   .O(to_level3[329]),
   .I0(level4_in[1974]),
   .I1(level4_in[1975]),
   .I2(level4_in[1976]),
   .I3(level4_in[1977]),
   .I4(level4_in[1978]),
   .I5(level4_in[1979])
);

LUT6 #(
   .INIT(64'h0bd723230bd72323)  
) LUT6_inst8106 (
   .O(to_level3[330]),
   .I0(level4_in[1980]),
   .I1(level4_in[1981]),
   .I2(level4_in[1982]),
   .I3(level4_in[1983]),
   .I4(level4_in[1984]),
   .I5(level4_in[1985])
);

LUT6 #(
   .INIT(64'ha21f12c7a21f12c7)  
) LUT6_inst8107 (
   .O(to_level3[331]),
   .I0(level4_in[1986]),
   .I1(level4_in[1987]),
   .I2(level4_in[1988]),
   .I3(level4_in[1989]),
   .I4(level4_in[1990]),
   .I5(level4_in[1991])
);

LUT6 #(
   .INIT(64'hf58fadb3f58fadb3)  
) LUT6_inst8108 (
   .O(to_level3[332]),
   .I0(level4_in[1992]),
   .I1(level4_in[1993]),
   .I2(level4_in[1994]),
   .I3(level4_in[1995]),
   .I4(level4_in[1996]),
   .I5(level4_in[1997])
);

LUT6 #(
   .INIT(64'h430800a5430800a5)  
) LUT6_inst8109 (
   .O(to_level3[333]),
   .I0(level4_in[1998]),
   .I1(level4_in[1999]),
   .I2(level4_in[2000]),
   .I3(level4_in[2001]),
   .I4(level4_in[2002]),
   .I5(level4_in[2003])
);

LUT6 #(
   .INIT(64'h9b5464319b546431)  
) LUT6_inst8110 (
   .O(to_level3[334]),
   .I0(level4_in[2004]),
   .I1(level4_in[2005]),
   .I2(level4_in[2006]),
   .I3(level4_in[2007]),
   .I4(level4_in[2008]),
   .I5(level4_in[2009])
);

LUT6 #(
   .INIT(64'h07f9587207f95872)  
) LUT6_inst8111 (
   .O(to_level3[335]),
   .I0(level4_in[2010]),
   .I1(level4_in[2011]),
   .I2(level4_in[2012]),
   .I3(level4_in[2013]),
   .I4(level4_in[2014]),
   .I5(level4_in[2015])
);

LUT6 #(
   .INIT(64'h3b26c10e3b26c10e)  
) LUT6_inst8112 (
   .O(to_level3[336]),
   .I0(level4_in[2016]),
   .I1(level4_in[2017]),
   .I2(level4_in[2018]),
   .I3(level4_in[2019]),
   .I4(level4_in[2020]),
   .I5(level4_in[2021])
);

LUT6 #(
   .INIT(64'h0f31d50b0f31d50b)  
) LUT6_inst8113 (
   .O(to_level3[337]),
   .I0(level4_in[2022]),
   .I1(level4_in[2023]),
   .I2(level4_in[2024]),
   .I3(level4_in[2025]),
   .I4(level4_in[2026]),
   .I5(level4_in[2027])
);

LUT6 #(
   .INIT(64'h609121d8609121d8)  
) LUT6_inst8114 (
   .O(to_level3[338]),
   .I0(level4_in[2028]),
   .I1(level4_in[2029]),
   .I2(level4_in[2030]),
   .I3(level4_in[2031]),
   .I4(level4_in[2032]),
   .I5(level4_in[2033])
);

LUT6 #(
   .INIT(64'h04a3a6d304a3a6d3)  
) LUT6_inst8115 (
   .O(to_level3[339]),
   .I0(level4_in[2034]),
   .I1(level4_in[2035]),
   .I2(level4_in[2036]),
   .I3(level4_in[2037]),
   .I4(level4_in[2038]),
   .I5(level4_in[2039])
);

LUT6 #(
   .INIT(64'h999b5155999b5155)  
) LUT6_inst8116 (
   .O(to_level3[340]),
   .I0(level4_in[2040]),
   .I1(level4_in[2041]),
   .I2(level4_in[2042]),
   .I3(level4_in[2043]),
   .I4(level4_in[2044]),
   .I5(level4_in[2045])
);

LUT6 #(
   .INIT(64'h71e4543471e45434)  
) LUT6_inst8117 (
   .O(to_level3[341]),
   .I0(level4_in[2046]),
   .I1(level4_in[2047]),
   .I2(level4_in[2048]),
   .I3(level4_in[2049]),
   .I4(level4_in[2050]),
   .I5(level4_in[2051])
);

LUT6 #(
   .INIT(64'ha46cb98ca46cb98c)  
) LUT6_inst8118 (
   .O(to_level3[342]),
   .I0(level4_in[2052]),
   .I1(level4_in[2053]),
   .I2(level4_in[2054]),
   .I3(level4_in[2055]),
   .I4(level4_in[2056]),
   .I5(level4_in[2057])
);

LUT6 #(
   .INIT(64'h7d8af0347d8af034)  
) LUT6_inst8119 (
   .O(to_level3[343]),
   .I0(level4_in[2058]),
   .I1(level4_in[2059]),
   .I2(level4_in[2060]),
   .I3(level4_in[2061]),
   .I4(level4_in[2062]),
   .I5(level4_in[2063])
);

LUT6 #(
   .INIT(64'h756a1fef756a1fef)  
) LUT6_inst8120 (
   .O(to_level3[344]),
   .I0(level4_in[2064]),
   .I1(level4_in[2065]),
   .I2(level4_in[2066]),
   .I3(level4_in[2067]),
   .I4(level4_in[2068]),
   .I5(level4_in[2069])
);

LUT6 #(
   .INIT(64'hf3e45be4f3e45be4)  
) LUT6_inst8121 (
   .O(to_level3[345]),
   .I0(level4_in[2070]),
   .I1(level4_in[2071]),
   .I2(level4_in[2072]),
   .I3(level4_in[2073]),
   .I4(level4_in[2074]),
   .I5(level4_in[2075])
);

LUT6 #(
   .INIT(64'hc6d13c65c6d13c65)  
) LUT6_inst8122 (
   .O(to_level3[346]),
   .I0(level4_in[2076]),
   .I1(level4_in[2077]),
   .I2(level4_in[2078]),
   .I3(level4_in[2079]),
   .I4(level4_in[2080]),
   .I5(level4_in[2081])
);

LUT6 #(
   .INIT(64'h1e97ee941e97ee94)  
) LUT6_inst8123 (
   .O(to_level3[347]),
   .I0(level4_in[2082]),
   .I1(level4_in[2083]),
   .I2(level4_in[2084]),
   .I3(level4_in[2085]),
   .I4(level4_in[2086]),
   .I5(level4_in[2087])
);

LUT6 #(
   .INIT(64'h6b6d8be46b6d8be4)  
) LUT6_inst8124 (
   .O(to_level3[348]),
   .I0(level4_in[2088]),
   .I1(level4_in[2089]),
   .I2(level4_in[2090]),
   .I3(level4_in[2091]),
   .I4(level4_in[2092]),
   .I5(level4_in[2093])
);

LUT6 #(
   .INIT(64'he44139b4e44139b4)  
) LUT6_inst8125 (
   .O(to_level3[349]),
   .I0(level4_in[2094]),
   .I1(level4_in[2095]),
   .I2(level4_in[2096]),
   .I3(level4_in[2097]),
   .I4(level4_in[2098]),
   .I5(level4_in[2099])
);

LUT6 #(
   .INIT(64'h50987acd50987acd)  
) LUT6_inst8126 (
   .O(to_level3[350]),
   .I0(level4_in[2100]),
   .I1(level4_in[2101]),
   .I2(level4_in[2102]),
   .I3(level4_in[2103]),
   .I4(level4_in[2104]),
   .I5(level4_in[2105])
);

LUT6 #(
   .INIT(64'hdd1ec615dd1ec615)  
) LUT6_inst8127 (
   .O(to_level3[351]),
   .I0(level4_in[2106]),
   .I1(level4_in[2107]),
   .I2(level4_in[2108]),
   .I3(level4_in[2109]),
   .I4(level4_in[2110]),
   .I5(level4_in[2111])
);

LUT6 #(
   .INIT(64'hf0ec9473f0ec9473)  
) LUT6_inst8128 (
   .O(to_level3[352]),
   .I0(level4_in[2112]),
   .I1(level4_in[2113]),
   .I2(level4_in[2114]),
   .I3(level4_in[2115]),
   .I4(level4_in[2116]),
   .I5(level4_in[2117])
);

LUT6 #(
   .INIT(64'hbf953b01bf953b01)  
) LUT6_inst8129 (
   .O(to_level3[353]),
   .I0(level4_in[2118]),
   .I1(level4_in[2119]),
   .I2(level4_in[2120]),
   .I3(level4_in[2121]),
   .I4(level4_in[2122]),
   .I5(level4_in[2123])
);

LUT6 #(
   .INIT(64'h12a5b59612a5b596)  
) LUT6_inst8130 (
   .O(to_level3[354]),
   .I0(level4_in[2124]),
   .I1(level4_in[2125]),
   .I2(level4_in[2126]),
   .I3(level4_in[2127]),
   .I4(level4_in[2128]),
   .I5(level4_in[2129])
);

LUT6 #(
   .INIT(64'he7d18f81e7d18f81)  
) LUT6_inst8131 (
   .O(to_level3[355]),
   .I0(level4_in[2130]),
   .I1(level4_in[2131]),
   .I2(level4_in[2132]),
   .I3(level4_in[2133]),
   .I4(level4_in[2134]),
   .I5(level4_in[2135])
);

LUT6 #(
   .INIT(64'h02871cbf02871cbf)  
) LUT6_inst8132 (
   .O(to_level3[356]),
   .I0(level4_in[2136]),
   .I1(level4_in[2137]),
   .I2(level4_in[2138]),
   .I3(level4_in[2139]),
   .I4(level4_in[2140]),
   .I5(level4_in[2141])
);

LUT6 #(
   .INIT(64'h45a9033d45a9033d)  
) LUT6_inst8133 (
   .O(to_level3[357]),
   .I0(level4_in[2142]),
   .I1(level4_in[2143]),
   .I2(level4_in[2144]),
   .I3(level4_in[2145]),
   .I4(level4_in[2146]),
   .I5(level4_in[2147])
);

LUT6 #(
   .INIT(64'hd85a3fd6d85a3fd6)  
) LUT6_inst8134 (
   .O(to_level3[358]),
   .I0(level4_in[2148]),
   .I1(level4_in[2149]),
   .I2(level4_in[2150]),
   .I3(level4_in[2151]),
   .I4(level4_in[2152]),
   .I5(level4_in[2153])
);

LUT6 #(
   .INIT(64'h92deb0c392deb0c3)  
) LUT6_inst8135 (
   .O(to_level3[359]),
   .I0(level4_in[2154]),
   .I1(level4_in[2155]),
   .I2(level4_in[2156]),
   .I3(level4_in[2157]),
   .I4(level4_in[2158]),
   .I5(level4_in[2159])
);

LUT6 #(
   .INIT(64'h7660566f7660566f)  
) LUT6_inst8136 (
   .O(to_level3[360]),
   .I0(level4_in[2160]),
   .I1(level4_in[2161]),
   .I2(level4_in[2162]),
   .I3(level4_in[2163]),
   .I4(level4_in[2164]),
   .I5(level4_in[2165])
);

LUT6 #(
   .INIT(64'h5fe11eaf5fe11eaf)  
) LUT6_inst8137 (
   .O(to_level3[361]),
   .I0(level4_in[2166]),
   .I1(level4_in[2167]),
   .I2(level4_in[2168]),
   .I3(level4_in[2169]),
   .I4(level4_in[2170]),
   .I5(level4_in[2171])
);

LUT6 #(
   .INIT(64'hb2848875b2848875)  
) LUT6_inst8138 (
   .O(to_level3[362]),
   .I0(level4_in[2172]),
   .I1(level4_in[2173]),
   .I2(level4_in[2174]),
   .I3(level4_in[2175]),
   .I4(level4_in[2176]),
   .I5(level4_in[2177])
);

LUT6 #(
   .INIT(64'h4ca0919b4ca0919b)  
) LUT6_inst8139 (
   .O(to_level3[363]),
   .I0(level4_in[2178]),
   .I1(level4_in[2179]),
   .I2(level4_in[2180]),
   .I3(level4_in[2181]),
   .I4(level4_in[2182]),
   .I5(level4_in[2183])
);

LUT6 #(
   .INIT(64'h6c1172806c117280)  
) LUT6_inst8140 (
   .O(to_level3[364]),
   .I0(level4_in[2184]),
   .I1(level4_in[2185]),
   .I2(level4_in[2186]),
   .I3(level4_in[2187]),
   .I4(level4_in[2188]),
   .I5(level4_in[2189])
);

LUT6 #(
   .INIT(64'h020e7f72020e7f72)  
) LUT6_inst8141 (
   .O(to_level3[365]),
   .I0(level4_in[2190]),
   .I1(level4_in[2191]),
   .I2(level4_in[2192]),
   .I3(level4_in[2193]),
   .I4(level4_in[2194]),
   .I5(level4_in[2195])
);

LUT6 #(
   .INIT(64'hcc5d0332cc5d0332)  
) LUT6_inst8142 (
   .O(to_level3[366]),
   .I0(level4_in[2196]),
   .I1(level4_in[2197]),
   .I2(level4_in[2198]),
   .I3(level4_in[2199]),
   .I4(level4_in[2200]),
   .I5(level4_in[2201])
);

LUT6 #(
   .INIT(64'h9d3e1c9f9d3e1c9f)  
) LUT6_inst8143 (
   .O(to_level3[367]),
   .I0(level4_in[2202]),
   .I1(level4_in[2203]),
   .I2(level4_in[2204]),
   .I3(level4_in[2205]),
   .I4(level4_in[2206]),
   .I5(level4_in[2207])
);

LUT6 #(
   .INIT(64'h2b7314c12b7314c1)  
) LUT6_inst8144 (
   .O(to_level3[368]),
   .I0(level4_in[2208]),
   .I1(level4_in[2209]),
   .I2(level4_in[2210]),
   .I3(level4_in[2211]),
   .I4(level4_in[2212]),
   .I5(level4_in[2213])
);

LUT6 #(
   .INIT(64'h681de5b5681de5b5)  
) LUT6_inst8145 (
   .O(to_level3[369]),
   .I0(level4_in[2214]),
   .I1(level4_in[2215]),
   .I2(level4_in[2216]),
   .I3(level4_in[2217]),
   .I4(level4_in[2218]),
   .I5(level4_in[2219])
);

LUT6 #(
   .INIT(64'h7a8cc4cf7a8cc4cf)  
) LUT6_inst8146 (
   .O(to_level3[370]),
   .I0(level4_in[2220]),
   .I1(level4_in[2221]),
   .I2(level4_in[2222]),
   .I3(level4_in[2223]),
   .I4(level4_in[2224]),
   .I5(level4_in[2225])
);

LUT6 #(
   .INIT(64'h54ecb85954ecb859)  
) LUT6_inst8147 (
   .O(to_level3[371]),
   .I0(level4_in[2226]),
   .I1(level4_in[2227]),
   .I2(level4_in[2228]),
   .I3(level4_in[2229]),
   .I4(level4_in[2230]),
   .I5(level4_in[2231])
);

LUT6 #(
   .INIT(64'h21db9fc721db9fc7)  
) LUT6_inst8148 (
   .O(to_level3[372]),
   .I0(level4_in[2232]),
   .I1(level4_in[2233]),
   .I2(level4_in[2234]),
   .I3(level4_in[2235]),
   .I4(level4_in[2236]),
   .I5(level4_in[2237])
);

LUT6 #(
   .INIT(64'he5c9c17de5c9c17d)  
) LUT6_inst8149 (
   .O(to_level3[373]),
   .I0(level4_in[2238]),
   .I1(level4_in[2239]),
   .I2(level4_in[2240]),
   .I3(level4_in[2241]),
   .I4(level4_in[2242]),
   .I5(level4_in[2243])
);

LUT6 #(
   .INIT(64'h47f47dc447f47dc4)  
) LUT6_inst8150 (
   .O(to_level3[374]),
   .I0(level4_in[2244]),
   .I1(level4_in[2245]),
   .I2(level4_in[2246]),
   .I3(level4_in[2247]),
   .I4(level4_in[2248]),
   .I5(level4_in[2249])
);

LUT6 #(
   .INIT(64'h697ab148697ab148)  
) LUT6_inst8151 (
   .O(to_level3[375]),
   .I0(level4_in[2250]),
   .I1(level4_in[2251]),
   .I2(level4_in[2252]),
   .I3(level4_in[2253]),
   .I4(level4_in[2254]),
   .I5(level4_in[2255])
);

LUT6 #(
   .INIT(64'he9ea072ce9ea072c)  
) LUT6_inst8152 (
   .O(to_level3[376]),
   .I0(level4_in[2256]),
   .I1(level4_in[2257]),
   .I2(level4_in[2258]),
   .I3(level4_in[2259]),
   .I4(level4_in[2260]),
   .I5(level4_in[2261])
);

LUT6 #(
   .INIT(64'h05e8179105e81791)  
) LUT6_inst8153 (
   .O(to_level3[377]),
   .I0(level4_in[2262]),
   .I1(level4_in[2263]),
   .I2(level4_in[2264]),
   .I3(level4_in[2265]),
   .I4(level4_in[2266]),
   .I5(level4_in[2267])
);

LUT6 #(
   .INIT(64'hd72464bbd72464bb)  
) LUT6_inst8154 (
   .O(to_level3[378]),
   .I0(level4_in[2268]),
   .I1(level4_in[2269]),
   .I2(level4_in[2270]),
   .I3(level4_in[2271]),
   .I4(level4_in[2272]),
   .I5(level4_in[2273])
);

LUT6 #(
   .INIT(64'hdd050fbcdd050fbc)  
) LUT6_inst8155 (
   .O(to_level3[379]),
   .I0(level4_in[2274]),
   .I1(level4_in[2275]),
   .I2(level4_in[2276]),
   .I3(level4_in[2277]),
   .I4(level4_in[2278]),
   .I5(level4_in[2279])
);

LUT6 #(
   .INIT(64'h21dde03d21dde03d)  
) LUT6_inst8156 (
   .O(to_level3[380]),
   .I0(level4_in[2280]),
   .I1(level4_in[2281]),
   .I2(level4_in[2282]),
   .I3(level4_in[2283]),
   .I4(level4_in[2284]),
   .I5(level4_in[2285])
);

LUT6 #(
   .INIT(64'h5eec98ff5eec98ff)  
) LUT6_inst8157 (
   .O(to_level3[381]),
   .I0(level4_in[2286]),
   .I1(level4_in[2287]),
   .I2(level4_in[2288]),
   .I3(level4_in[2289]),
   .I4(level4_in[2290]),
   .I5(level4_in[2291])
);

LUT6 #(
   .INIT(64'hf9e89b06f9e89b06)  
) LUT6_inst8158 (
   .O(to_level3[382]),
   .I0(level4_in[2292]),
   .I1(level4_in[2293]),
   .I2(level4_in[2294]),
   .I3(level4_in[2295]),
   .I4(level4_in[2296]),
   .I5(level4_in[2297])
);

LUT6 #(
   .INIT(64'hf8160e0ff8160e0f)  
) LUT6_inst8159 (
   .O(to_level3[383]),
   .I0(level4_in[2298]),
   .I1(level4_in[2299]),
   .I2(level4_in[2300]),
   .I3(level4_in[2301]),
   .I4(level4_in[2302]),
   .I5(level4_in[2303])
);

LUT6 #(
   .INIT(64'hd320be7ed320be7e)  
) LUT6_inst8160 (
   .O(to_level3[384]),
   .I0(level4_in[2304]),
   .I1(level4_in[2305]),
   .I2(level4_in[2306]),
   .I3(level4_in[2307]),
   .I4(level4_in[2308]),
   .I5(level4_in[2309])
);

LUT6 #(
   .INIT(64'hbb85a638bb85a638)  
) LUT6_inst8161 (
   .O(to_level3[385]),
   .I0(level4_in[2310]),
   .I1(level4_in[2311]),
   .I2(level4_in[2312]),
   .I3(level4_in[2313]),
   .I4(level4_in[2314]),
   .I5(level4_in[2315])
);

LUT6 #(
   .INIT(64'hb07ab909b07ab909)  
) LUT6_inst8162 (
   .O(to_level3[386]),
   .I0(level4_in[2316]),
   .I1(level4_in[2317]),
   .I2(level4_in[2318]),
   .I3(level4_in[2319]),
   .I4(level4_in[2320]),
   .I5(level4_in[2321])
);

LUT6 #(
   .INIT(64'h0db2185b0db2185b)  
) LUT6_inst8163 (
   .O(to_level3[387]),
   .I0(level4_in[2322]),
   .I1(level4_in[2323]),
   .I2(level4_in[2324]),
   .I3(level4_in[2325]),
   .I4(level4_in[2326]),
   .I5(level4_in[2327])
);

LUT6 #(
   .INIT(64'h01c8582401c85824)  
) LUT6_inst8164 (
   .O(to_level3[388]),
   .I0(level4_in[2328]),
   .I1(level4_in[2329]),
   .I2(level4_in[2330]),
   .I3(level4_in[2331]),
   .I4(level4_in[2332]),
   .I5(level4_in[2333])
);

LUT6 #(
   .INIT(64'h04e046f304e046f3)  
) LUT6_inst8165 (
   .O(to_level3[389]),
   .I0(level4_in[2334]),
   .I1(level4_in[2335]),
   .I2(level4_in[2336]),
   .I3(level4_in[2337]),
   .I4(level4_in[2338]),
   .I5(level4_in[2339])
);

LUT6 #(
   .INIT(64'h1b7df2ed1b7df2ed)  
) LUT6_inst8166 (
   .O(to_level3[390]),
   .I0(level4_in[2340]),
   .I1(level4_in[2341]),
   .I2(level4_in[2342]),
   .I3(level4_in[2343]),
   .I4(level4_in[2344]),
   .I5(level4_in[2345])
);

LUT6 #(
   .INIT(64'ha43ce9a1a43ce9a1)  
) LUT6_inst8167 (
   .O(to_level3[391]),
   .I0(level4_in[2346]),
   .I1(level4_in[2347]),
   .I2(level4_in[2348]),
   .I3(level4_in[2349]),
   .I4(level4_in[2350]),
   .I5(level4_in[2351])
);

LUT6 #(
   .INIT(64'hd62a617cd62a617c)  
) LUT6_inst8168 (
   .O(to_level3[392]),
   .I0(level4_in[2352]),
   .I1(level4_in[2353]),
   .I2(level4_in[2354]),
   .I3(level4_in[2355]),
   .I4(level4_in[2356]),
   .I5(level4_in[2357])
);

LUT6 #(
   .INIT(64'h86a42ad986a42ad9)  
) LUT6_inst8169 (
   .O(to_level3[393]),
   .I0(level4_in[2358]),
   .I1(level4_in[2359]),
   .I2(level4_in[2360]),
   .I3(level4_in[2361]),
   .I4(level4_in[2362]),
   .I5(level4_in[2363])
);

LUT6 #(
   .INIT(64'h60f46dcf60f46dcf)  
) LUT6_inst8170 (
   .O(to_level3[394]),
   .I0(level4_in[2364]),
   .I1(level4_in[2365]),
   .I2(level4_in[2366]),
   .I3(level4_in[2367]),
   .I4(level4_in[2368]),
   .I5(level4_in[2369])
);

LUT6 #(
   .INIT(64'h82620d1682620d16)  
) LUT6_inst8171 (
   .O(to_level3[395]),
   .I0(level4_in[2370]),
   .I1(level4_in[2371]),
   .I2(level4_in[2372]),
   .I3(level4_in[2373]),
   .I4(level4_in[2374]),
   .I5(level4_in[2375])
);

LUT6 #(
   .INIT(64'hb3e44274b3e44274)  
) LUT6_inst8172 (
   .O(to_level3[396]),
   .I0(level4_in[2376]),
   .I1(level4_in[2377]),
   .I2(level4_in[2378]),
   .I3(level4_in[2379]),
   .I4(level4_in[2380]),
   .I5(level4_in[2381])
);

LUT6 #(
   .INIT(64'h78c6893a78c6893a)  
) LUT6_inst8173 (
   .O(to_level3[397]),
   .I0(level4_in[2382]),
   .I1(level4_in[2383]),
   .I2(level4_in[2384]),
   .I3(level4_in[2385]),
   .I4(level4_in[2386]),
   .I5(level4_in[2387])
);

LUT6 #(
   .INIT(64'h2e7d90c22e7d90c2)  
) LUT6_inst8174 (
   .O(to_level3[398]),
   .I0(level4_in[2388]),
   .I1(level4_in[2389]),
   .I2(level4_in[2390]),
   .I3(level4_in[2391]),
   .I4(level4_in[2392]),
   .I5(level4_in[2393])
);

LUT6 #(
   .INIT(64'h8070a1738070a173)  
) LUT6_inst8175 (
   .O(to_level3[399]),
   .I0(level4_in[2394]),
   .I1(level4_in[2395]),
   .I2(level4_in[2396]),
   .I3(level4_in[2397]),
   .I4(level4_in[2398]),
   .I5(level4_in[2399])
);

LUT6 #(
   .INIT(64'h2334c0122334c012)  
) LUT6_inst8176 (
   .O(to_level3[400]),
   .I0(level4_in[2400]),
   .I1(level4_in[2401]),
   .I2(level4_in[2402]),
   .I3(level4_in[2403]),
   .I4(level4_in[2404]),
   .I5(level4_in[2405])
);

LUT6 #(
   .INIT(64'h3a9875793a987579)  
) LUT6_inst8177 (
   .O(to_level3[401]),
   .I0(level4_in[2406]),
   .I1(level4_in[2407]),
   .I2(level4_in[2408]),
   .I3(level4_in[2409]),
   .I4(level4_in[2410]),
   .I5(level4_in[2411])
);

LUT6 #(
   .INIT(64'hedc1c2ccedc1c2cc)  
) LUT6_inst8178 (
   .O(to_level3[402]),
   .I0(level4_in[2412]),
   .I1(level4_in[2413]),
   .I2(level4_in[2414]),
   .I3(level4_in[2415]),
   .I4(level4_in[2416]),
   .I5(level4_in[2417])
);

LUT6 #(
   .INIT(64'h92fd828592fd8285)  
) LUT6_inst8179 (
   .O(to_level3[403]),
   .I0(level4_in[2418]),
   .I1(level4_in[2419]),
   .I2(level4_in[2420]),
   .I3(level4_in[2421]),
   .I4(level4_in[2422]),
   .I5(level4_in[2423])
);

LUT6 #(
   .INIT(64'hdbb2a35edbb2a35e)  
) LUT6_inst8180 (
   .O(to_level3[404]),
   .I0(level4_in[2424]),
   .I1(level4_in[2425]),
   .I2(level4_in[2426]),
   .I3(level4_in[2427]),
   .I4(level4_in[2428]),
   .I5(level4_in[2429])
);

LUT6 #(
   .INIT(64'h53f895ce53f895ce)  
) LUT6_inst8181 (
   .O(to_level3[405]),
   .I0(level4_in[2430]),
   .I1(level4_in[2431]),
   .I2(level4_in[2432]),
   .I3(level4_in[2433]),
   .I4(level4_in[2434]),
   .I5(level4_in[2435])
);

LUT6 #(
   .INIT(64'h5c29faa95c29faa9)  
) LUT6_inst8182 (
   .O(to_level3[406]),
   .I0(level4_in[2436]),
   .I1(level4_in[2437]),
   .I2(level4_in[2438]),
   .I3(level4_in[2439]),
   .I4(level4_in[2440]),
   .I5(level4_in[2441])
);

LUT6 #(
   .INIT(64'hf4ed2e10f4ed2e10)  
) LUT6_inst8183 (
   .O(to_level3[407]),
   .I0(level4_in[2442]),
   .I1(level4_in[2443]),
   .I2(level4_in[2444]),
   .I3(level4_in[2445]),
   .I4(level4_in[2446]),
   .I5(level4_in[2447])
);

LUT6 #(
   .INIT(64'h976402f6976402f6)  
) LUT6_inst8184 (
   .O(to_level3[408]),
   .I0(level4_in[2448]),
   .I1(level4_in[2449]),
   .I2(level4_in[2450]),
   .I3(level4_in[2451]),
   .I4(level4_in[2452]),
   .I5(level4_in[2453])
);

LUT6 #(
   .INIT(64'ha3002e56a3002e56)  
) LUT6_inst8185 (
   .O(to_level3[409]),
   .I0(level4_in[2454]),
   .I1(level4_in[2455]),
   .I2(level4_in[2456]),
   .I3(level4_in[2457]),
   .I4(level4_in[2458]),
   .I5(level4_in[2459])
);

LUT6 #(
   .INIT(64'h8558b1278558b127)  
) LUT6_inst8186 (
   .O(to_level3[410]),
   .I0(level4_in[2460]),
   .I1(level4_in[2461]),
   .I2(level4_in[2462]),
   .I3(level4_in[2463]),
   .I4(level4_in[2464]),
   .I5(level4_in[2465])
);

LUT6 #(
   .INIT(64'heba291a8eba291a8)  
) LUT6_inst8187 (
   .O(to_level3[411]),
   .I0(level4_in[2466]),
   .I1(level4_in[2467]),
   .I2(level4_in[2468]),
   .I3(level4_in[2469]),
   .I4(level4_in[2470]),
   .I5(level4_in[2471])
);

LUT6 #(
   .INIT(64'h5b8ae5bb5b8ae5bb)  
) LUT6_inst8188 (
   .O(to_level3[412]),
   .I0(level4_in[2472]),
   .I1(level4_in[2473]),
   .I2(level4_in[2474]),
   .I3(level4_in[2475]),
   .I4(level4_in[2476]),
   .I5(level4_in[2477])
);

LUT6 #(
   .INIT(64'h0367274203672742)  
) LUT6_inst8189 (
   .O(to_level3[413]),
   .I0(level4_in[2478]),
   .I1(level4_in[2479]),
   .I2(level4_in[2480]),
   .I3(level4_in[2481]),
   .I4(level4_in[2482]),
   .I5(level4_in[2483])
);

LUT6 #(
   .INIT(64'h665d4efc665d4efc)  
) LUT6_inst8190 (
   .O(to_level3[414]),
   .I0(level4_in[2484]),
   .I1(level4_in[2485]),
   .I2(level4_in[2486]),
   .I3(level4_in[2487]),
   .I4(level4_in[2488]),
   .I5(level4_in[2489])
);

LUT6 #(
   .INIT(64'he417bcdbe417bcdb)  
) LUT6_inst8191 (
   .O(to_level3[415]),
   .I0(level4_in[2490]),
   .I1(level4_in[2491]),
   .I2(level4_in[2492]),
   .I3(level4_in[2493]),
   .I4(level4_in[2494]),
   .I5(level4_in[2495])
);

LUT6 #(
   .INIT(64'h44f4c62544f4c625)  
) LUT6_inst8192 (
   .O(to_level3[416]),
   .I0(level4_in[2496]),
   .I1(level4_in[2497]),
   .I2(level4_in[2498]),
   .I3(level4_in[2499]),
   .I4(level4_in[2500]),
   .I5(level4_in[2501])
);

LUT6 #(
   .INIT(64'h9511367695113676)  
) LUT6_inst8193 (
   .O(to_level3[417]),
   .I0(level4_in[2502]),
   .I1(level4_in[2503]),
   .I2(level4_in[2504]),
   .I3(level4_in[2505]),
   .I4(level4_in[2506]),
   .I5(level4_in[2507])
);

LUT6 #(
   .INIT(64'h3ba58c9f3ba58c9f)  
) LUT6_inst8194 (
   .O(to_level3[418]),
   .I0(level4_in[2508]),
   .I1(level4_in[2509]),
   .I2(level4_in[2510]),
   .I3(level4_in[2511]),
   .I4(level4_in[2512]),
   .I5(level4_in[2513])
);

LUT6 #(
   .INIT(64'ha468edf7a468edf7)  
) LUT6_inst8195 (
   .O(to_level3[419]),
   .I0(level4_in[2514]),
   .I1(level4_in[2515]),
   .I2(level4_in[2516]),
   .I3(level4_in[2517]),
   .I4(level4_in[2518]),
   .I5(level4_in[2519])
);

LUT6 #(
   .INIT(64'hb8edeedcb8edeedc)  
) LUT6_inst8196 (
   .O(to_level3[420]),
   .I0(level4_in[2520]),
   .I1(level4_in[2521]),
   .I2(level4_in[2522]),
   .I3(level4_in[2523]),
   .I4(level4_in[2524]),
   .I5(level4_in[2525])
);

LUT6 #(
   .INIT(64'h629d84de629d84de)  
) LUT6_inst8197 (
   .O(to_level3[421]),
   .I0(level4_in[2526]),
   .I1(level4_in[2527]),
   .I2(level4_in[2528]),
   .I3(level4_in[2529]),
   .I4(level4_in[2530]),
   .I5(level4_in[2531])
);

LUT6 #(
   .INIT(64'h554af39e554af39e)  
) LUT6_inst8198 (
   .O(to_level3[422]),
   .I0(level4_in[2532]),
   .I1(level4_in[2533]),
   .I2(level4_in[2534]),
   .I3(level4_in[2535]),
   .I4(level4_in[2536]),
   .I5(level4_in[2537])
);

LUT6 #(
   .INIT(64'hea3a4471ea3a4471)  
) LUT6_inst8199 (
   .O(to_level3[423]),
   .I0(level4_in[2538]),
   .I1(level4_in[2539]),
   .I2(level4_in[2540]),
   .I3(level4_in[2541]),
   .I4(level4_in[2542]),
   .I5(level4_in[2543])
);

LUT6 #(
   .INIT(64'h26eb352226eb3522)  
) LUT6_inst8200 (
   .O(to_level3[424]),
   .I0(level4_in[2544]),
   .I1(level4_in[2545]),
   .I2(level4_in[2546]),
   .I3(level4_in[2547]),
   .I4(level4_in[2548]),
   .I5(level4_in[2549])
);

LUT6 #(
   .INIT(64'hfda80728fda80728)  
) LUT6_inst8201 (
   .O(to_level3[425]),
   .I0(level4_in[2550]),
   .I1(level4_in[2551]),
   .I2(level4_in[2552]),
   .I3(level4_in[2553]),
   .I4(level4_in[2554]),
   .I5(level4_in[2555])
);

LUT6 #(
   .INIT(64'h4f61ec4b4f61ec4b)  
) LUT6_inst8202 (
   .O(to_level3[426]),
   .I0(level4_in[2556]),
   .I1(level4_in[2557]),
   .I2(level4_in[2558]),
   .I3(level4_in[2559]),
   .I4(level4_in[2560]),
   .I5(level4_in[2561])
);

LUT6 #(
   .INIT(64'h9b7f90729b7f9072)  
) LUT6_inst8203 (
   .O(to_level3[427]),
   .I0(level4_in[2562]),
   .I1(level4_in[2563]),
   .I2(level4_in[2564]),
   .I3(level4_in[2565]),
   .I4(level4_in[2566]),
   .I5(level4_in[2567])
);

LUT6 #(
   .INIT(64'h13f2278a13f2278a)  
) LUT6_inst8204 (
   .O(to_level3[428]),
   .I0(level4_in[2568]),
   .I1(level4_in[2569]),
   .I2(level4_in[2570]),
   .I3(level4_in[2571]),
   .I4(level4_in[2572]),
   .I5(level4_in[2573])
);

LUT6 #(
   .INIT(64'hcf8b6816cf8b6816)  
) LUT6_inst8205 (
   .O(to_level3[429]),
   .I0(level4_in[2574]),
   .I1(level4_in[2575]),
   .I2(level4_in[2576]),
   .I3(level4_in[2577]),
   .I4(level4_in[2578]),
   .I5(level4_in[2579])
);

LUT6 #(
   .INIT(64'hdacc240bdacc240b)  
) LUT6_inst8206 (
   .O(to_level3[430]),
   .I0(level4_in[2580]),
   .I1(level4_in[2581]),
   .I2(level4_in[2582]),
   .I3(level4_in[2583]),
   .I4(level4_in[2584]),
   .I5(level4_in[2585])
);

LUT6 #(
   .INIT(64'hd7c72327d7c72327)  
) LUT6_inst8207 (
   .O(to_level3[431]),
   .I0(level4_in[2586]),
   .I1(level4_in[2587]),
   .I2(level4_in[2588]),
   .I3(level4_in[2589]),
   .I4(level4_in[2590]),
   .I5(level4_in[2591])
);

LUT6 #(
   .INIT(64'h5f930e1c5f930e1c)  
) LUT6_inst8208 (
   .O(to_level3[432]),
   .I0(level4_in[2592]),
   .I1(level4_in[2593]),
   .I2(level4_in[2594]),
   .I3(level4_in[2595]),
   .I4(level4_in[2596]),
   .I5(level4_in[2597])
);

LUT6 #(
   .INIT(64'h7edbb0407edbb040)  
) LUT6_inst8209 (
   .O(to_level3[433]),
   .I0(level4_in[2598]),
   .I1(level4_in[2599]),
   .I2(level4_in[2600]),
   .I3(level4_in[2601]),
   .I4(level4_in[2602]),
   .I5(level4_in[2603])
);

LUT6 #(
   .INIT(64'hc47a34fac47a34fa)  
) LUT6_inst8210 (
   .O(to_level3[434]),
   .I0(level4_in[2604]),
   .I1(level4_in[2605]),
   .I2(level4_in[2606]),
   .I3(level4_in[2607]),
   .I4(level4_in[2608]),
   .I5(level4_in[2609])
);

LUT6 #(
   .INIT(64'he6df2da0e6df2da0)  
) LUT6_inst8211 (
   .O(to_level3[435]),
   .I0(level4_in[2610]),
   .I1(level4_in[2611]),
   .I2(level4_in[2612]),
   .I3(level4_in[2613]),
   .I4(level4_in[2614]),
   .I5(level4_in[2615])
);

LUT6 #(
   .INIT(64'hd28b9616d28b9616)  
) LUT6_inst8212 (
   .O(to_level3[436]),
   .I0(level4_in[2616]),
   .I1(level4_in[2617]),
   .I2(level4_in[2618]),
   .I3(level4_in[2619]),
   .I4(level4_in[2620]),
   .I5(level4_in[2621])
);

LUT6 #(
   .INIT(64'he39af832e39af832)  
) LUT6_inst8213 (
   .O(to_level3[437]),
   .I0(level4_in[2622]),
   .I1(level4_in[2623]),
   .I2(level4_in[2624]),
   .I3(level4_in[2625]),
   .I4(level4_in[2626]),
   .I5(level4_in[2627])
);

LUT6 #(
   .INIT(64'h1f1559351f155935)  
) LUT6_inst8214 (
   .O(to_level3[438]),
   .I0(level4_in[2628]),
   .I1(level4_in[2629]),
   .I2(level4_in[2630]),
   .I3(level4_in[2631]),
   .I4(level4_in[2632]),
   .I5(level4_in[2633])
);

LUT6 #(
   .INIT(64'h27ec41c627ec41c6)  
) LUT6_inst8215 (
   .O(to_level3[439]),
   .I0(level4_in[2634]),
   .I1(level4_in[2635]),
   .I2(level4_in[2636]),
   .I3(level4_in[2637]),
   .I4(level4_in[2638]),
   .I5(level4_in[2639])
);

LUT6 #(
   .INIT(64'hbbf25988bbf25988)  
) LUT6_inst8216 (
   .O(to_level3[440]),
   .I0(level4_in[2640]),
   .I1(level4_in[2641]),
   .I2(level4_in[2642]),
   .I3(level4_in[2643]),
   .I4(level4_in[2644]),
   .I5(level4_in[2645])
);

LUT6 #(
   .INIT(64'h1557ba4d1557ba4d)  
) LUT6_inst8217 (
   .O(to_level3[441]),
   .I0(level4_in[2646]),
   .I1(level4_in[2647]),
   .I2(level4_in[2648]),
   .I3(level4_in[2649]),
   .I4(level4_in[2650]),
   .I5(level4_in[2651])
);

LUT6 #(
   .INIT(64'he8754dc2e8754dc2)  
) LUT6_inst8218 (
   .O(to_level3[442]),
   .I0(level4_in[2652]),
   .I1(level4_in[2653]),
   .I2(level4_in[2654]),
   .I3(level4_in[2655]),
   .I4(level4_in[2656]),
   .I5(level4_in[2657])
);

LUT6 #(
   .INIT(64'h43b6df8243b6df82)  
) LUT6_inst8219 (
   .O(to_level3[443]),
   .I0(level4_in[2658]),
   .I1(level4_in[2659]),
   .I2(level4_in[2660]),
   .I3(level4_in[2661]),
   .I4(level4_in[2662]),
   .I5(level4_in[2663])
);

LUT6 #(
   .INIT(64'h149f8568149f8568)  
) LUT6_inst8220 (
   .O(to_level3[444]),
   .I0(level4_in[2664]),
   .I1(level4_in[2665]),
   .I2(level4_in[2666]),
   .I3(level4_in[2667]),
   .I4(level4_in[2668]),
   .I5(level4_in[2669])
);

LUT6 #(
   .INIT(64'h3eec11c53eec11c5)  
) LUT6_inst8221 (
   .O(to_level3[445]),
   .I0(level4_in[2670]),
   .I1(level4_in[2671]),
   .I2(level4_in[2672]),
   .I3(level4_in[2673]),
   .I4(level4_in[2674]),
   .I5(level4_in[2675])
);

LUT6 #(
   .INIT(64'ha40f8e97a40f8e97)  
) LUT6_inst8222 (
   .O(to_level3[446]),
   .I0(level4_in[2676]),
   .I1(level4_in[2677]),
   .I2(level4_in[2678]),
   .I3(level4_in[2679]),
   .I4(level4_in[2680]),
   .I5(level4_in[2681])
);

LUT6 #(
   .INIT(64'hea3cec84ea3cec84)  
) LUT6_inst8223 (
   .O(to_level3[447]),
   .I0(level4_in[2682]),
   .I1(level4_in[2683]),
   .I2(level4_in[2684]),
   .I3(level4_in[2685]),
   .I4(level4_in[2686]),
   .I5(level4_in[2687])
);

LUT6 #(
   .INIT(64'h7d64e5817d64e581)  
) LUT6_inst8224 (
   .O(to_level3[448]),
   .I0(level4_in[2688]),
   .I1(level4_in[2689]),
   .I2(level4_in[2690]),
   .I3(level4_in[2691]),
   .I4(level4_in[2692]),
   .I5(level4_in[2693])
);

LUT6 #(
   .INIT(64'h8671f6e58671f6e5)  
) LUT6_inst8225 (
   .O(to_level3[449]),
   .I0(level4_in[2694]),
   .I1(level4_in[2695]),
   .I2(level4_in[2696]),
   .I3(level4_in[2697]),
   .I4(level4_in[2698]),
   .I5(level4_in[2699])
);

LUT6 #(
   .INIT(64'hb0625973b0625973)  
) LUT6_inst8226 (
   .O(to_level3[450]),
   .I0(level4_in[2700]),
   .I1(level4_in[2701]),
   .I2(level4_in[2702]),
   .I3(level4_in[2703]),
   .I4(level4_in[2704]),
   .I5(level4_in[2705])
);

LUT6 #(
   .INIT(64'he8fc2990e8fc2990)  
) LUT6_inst8227 (
   .O(to_level3[451]),
   .I0(level4_in[2706]),
   .I1(level4_in[2707]),
   .I2(level4_in[2708]),
   .I3(level4_in[2709]),
   .I4(level4_in[2710]),
   .I5(level4_in[2711])
);

LUT6 #(
   .INIT(64'h50e0f8b250e0f8b2)  
) LUT6_inst8228 (
   .O(to_level3[452]),
   .I0(level4_in[2712]),
   .I1(level4_in[2713]),
   .I2(level4_in[2714]),
   .I3(level4_in[2715]),
   .I4(level4_in[2716]),
   .I5(level4_in[2717])
);

LUT6 #(
   .INIT(64'h78cad7e978cad7e9)  
) LUT6_inst8229 (
   .O(to_level3[453]),
   .I0(level4_in[2718]),
   .I1(level4_in[2719]),
   .I2(level4_in[2720]),
   .I3(level4_in[2721]),
   .I4(level4_in[2722]),
   .I5(level4_in[2723])
);

LUT6 #(
   .INIT(64'hc2dc6a14c2dc6a14)  
) LUT6_inst8230 (
   .O(to_level3[454]),
   .I0(level4_in[2724]),
   .I1(level4_in[2725]),
   .I2(level4_in[2726]),
   .I3(level4_in[2727]),
   .I4(level4_in[2728]),
   .I5(level4_in[2729])
);

LUT6 #(
   .INIT(64'h6cd1fa2d6cd1fa2d)  
) LUT6_inst8231 (
   .O(to_level3[455]),
   .I0(level4_in[2730]),
   .I1(level4_in[2731]),
   .I2(level4_in[2732]),
   .I3(level4_in[2733]),
   .I4(level4_in[2734]),
   .I5(level4_in[2735])
);

LUT6 #(
   .INIT(64'h60dedbad60dedbad)  
) LUT6_inst8232 (
   .O(to_level3[456]),
   .I0(level4_in[2736]),
   .I1(level4_in[2737]),
   .I2(level4_in[2738]),
   .I3(level4_in[2739]),
   .I4(level4_in[2740]),
   .I5(level4_in[2741])
);

LUT6 #(
   .INIT(64'hbde8fda5bde8fda5)  
) LUT6_inst8233 (
   .O(to_level3[457]),
   .I0(level4_in[2742]),
   .I1(level4_in[2743]),
   .I2(level4_in[2744]),
   .I3(level4_in[2745]),
   .I4(level4_in[2746]),
   .I5(level4_in[2747])
);

LUT6 #(
   .INIT(64'h89d6311389d63113)  
) LUT6_inst8234 (
   .O(to_level3[458]),
   .I0(level4_in[2748]),
   .I1(level4_in[2749]),
   .I2(level4_in[2750]),
   .I3(level4_in[2751]),
   .I4(level4_in[2752]),
   .I5(level4_in[2753])
);

LUT6 #(
   .INIT(64'h830144d9830144d9)  
) LUT6_inst8235 (
   .O(to_level3[459]),
   .I0(level4_in[2754]),
   .I1(level4_in[2755]),
   .I2(level4_in[2756]),
   .I3(level4_in[2757]),
   .I4(level4_in[2758]),
   .I5(level4_in[2759])
);

LUT6 #(
   .INIT(64'h87854bec87854bec)  
) LUT6_inst8236 (
   .O(to_level3[460]),
   .I0(level4_in[2760]),
   .I1(level4_in[2761]),
   .I2(level4_in[2762]),
   .I3(level4_in[2763]),
   .I4(level4_in[2764]),
   .I5(level4_in[2765])
);

LUT6 #(
   .INIT(64'h0146163001461630)  
) LUT6_inst8237 (
   .O(to_level3[461]),
   .I0(level4_in[2766]),
   .I1(level4_in[2767]),
   .I2(level4_in[2768]),
   .I3(level4_in[2769]),
   .I4(level4_in[2770]),
   .I5(level4_in[2771])
);

LUT6 #(
   .INIT(64'hfb57ea18fb57ea18)  
) LUT6_inst8238 (
   .O(to_level3[462]),
   .I0(level4_in[2772]),
   .I1(level4_in[2773]),
   .I2(level4_in[2774]),
   .I3(level4_in[2775]),
   .I4(level4_in[2776]),
   .I5(level4_in[2777])
);

LUT6 #(
   .INIT(64'hbf4fcbe4bf4fcbe4)  
) LUT6_inst8239 (
   .O(to_level3[463]),
   .I0(level4_in[2778]),
   .I1(level4_in[2779]),
   .I2(level4_in[2780]),
   .I3(level4_in[2781]),
   .I4(level4_in[2782]),
   .I5(level4_in[2783])
);

LUT6 #(
   .INIT(64'hc7abd9e9c7abd9e9)  
) LUT6_inst8240 (
   .O(to_level3[464]),
   .I0(level4_in[2784]),
   .I1(level4_in[2785]),
   .I2(level4_in[2786]),
   .I3(level4_in[2787]),
   .I4(level4_in[2788]),
   .I5(level4_in[2789])
);

LUT6 #(
   .INIT(64'h5edfcf655edfcf65)  
) LUT6_inst8241 (
   .O(to_level3[465]),
   .I0(level4_in[2790]),
   .I1(level4_in[2791]),
   .I2(level4_in[2792]),
   .I3(level4_in[2793]),
   .I4(level4_in[2794]),
   .I5(level4_in[2795])
);

LUT6 #(
   .INIT(64'h38c0368138c03681)  
) LUT6_inst8242 (
   .O(to_level3[466]),
   .I0(level4_in[2796]),
   .I1(level4_in[2797]),
   .I2(level4_in[2798]),
   .I3(level4_in[2799]),
   .I4(level4_in[2800]),
   .I5(level4_in[2801])
);

LUT6 #(
   .INIT(64'h6bacc4c56bacc4c5)  
) LUT6_inst8243 (
   .O(to_level3[467]),
   .I0(level4_in[2802]),
   .I1(level4_in[2803]),
   .I2(level4_in[2804]),
   .I3(level4_in[2805]),
   .I4(level4_in[2806]),
   .I5(level4_in[2807])
);

LUT6 #(
   .INIT(64'h4e4f72374e4f7237)  
) LUT6_inst8244 (
   .O(to_level3[468]),
   .I0(level4_in[2808]),
   .I1(level4_in[2809]),
   .I2(level4_in[2810]),
   .I3(level4_in[2811]),
   .I4(level4_in[2812]),
   .I5(level4_in[2813])
);

LUT6 #(
   .INIT(64'hc2e905e3c2e905e3)  
) LUT6_inst8245 (
   .O(to_level3[469]),
   .I0(level4_in[2814]),
   .I1(level4_in[2815]),
   .I2(level4_in[2816]),
   .I3(level4_in[2817]),
   .I4(level4_in[2818]),
   .I5(level4_in[2819])
);

LUT6 #(
   .INIT(64'h88d294a388d294a3)  
) LUT6_inst8246 (
   .O(to_level3[470]),
   .I0(level4_in[2820]),
   .I1(level4_in[2821]),
   .I2(level4_in[2822]),
   .I3(level4_in[2823]),
   .I4(level4_in[2824]),
   .I5(level4_in[2825])
);

LUT6 #(
   .INIT(64'h3ba345953ba34595)  
) LUT6_inst8247 (
   .O(to_level3[471]),
   .I0(level4_in[2826]),
   .I1(level4_in[2827]),
   .I2(level4_in[2828]),
   .I3(level4_in[2829]),
   .I4(level4_in[2830]),
   .I5(level4_in[2831])
);

LUT6 #(
   .INIT(64'h5ec017fa5ec017fa)  
) LUT6_inst8248 (
   .O(to_level3[472]),
   .I0(level4_in[2832]),
   .I1(level4_in[2833]),
   .I2(level4_in[2834]),
   .I3(level4_in[2835]),
   .I4(level4_in[2836]),
   .I5(level4_in[2837])
);

LUT6 #(
   .INIT(64'h7616c5707616c570)  
) LUT6_inst8249 (
   .O(to_level3[473]),
   .I0(level4_in[2838]),
   .I1(level4_in[2839]),
   .I2(level4_in[2840]),
   .I3(level4_in[2841]),
   .I4(level4_in[2842]),
   .I5(level4_in[2843])
);

LUT6 #(
   .INIT(64'h3bc723c53bc723c5)  
) LUT6_inst8250 (
   .O(to_level3[474]),
   .I0(level4_in[2844]),
   .I1(level4_in[2845]),
   .I2(level4_in[2846]),
   .I3(level4_in[2847]),
   .I4(level4_in[2848]),
   .I5(level4_in[2849])
);

LUT6 #(
   .INIT(64'h1d3cc3641d3cc364)  
) LUT6_inst8251 (
   .O(to_level3[475]),
   .I0(level4_in[2850]),
   .I1(level4_in[2851]),
   .I2(level4_in[2852]),
   .I3(level4_in[2853]),
   .I4(level4_in[2854]),
   .I5(level4_in[2855])
);

LUT6 #(
   .INIT(64'h8526f87d8526f87d)  
) LUT6_inst8252 (
   .O(to_level3[476]),
   .I0(level4_in[2856]),
   .I1(level4_in[2857]),
   .I2(level4_in[2858]),
   .I3(level4_in[2859]),
   .I4(level4_in[2860]),
   .I5(level4_in[2861])
);

LUT6 #(
   .INIT(64'hea846f85ea846f85)  
) LUT6_inst8253 (
   .O(to_level3[477]),
   .I0(level4_in[2862]),
   .I1(level4_in[2863]),
   .I2(level4_in[2864]),
   .I3(level4_in[2865]),
   .I4(level4_in[2866]),
   .I5(level4_in[2867])
);

LUT6 #(
   .INIT(64'hfa189513fa189513)  
) LUT6_inst8254 (
   .O(to_level3[478]),
   .I0(level4_in[2868]),
   .I1(level4_in[2869]),
   .I2(level4_in[2870]),
   .I3(level4_in[2871]),
   .I4(level4_in[2872]),
   .I5(level4_in[2873])
);

LUT6 #(
   .INIT(64'hf5aeb654f5aeb654)  
) LUT6_inst8255 (
   .O(to_level3[479]),
   .I0(level4_in[2874]),
   .I1(level4_in[2875]),
   .I2(level4_in[2876]),
   .I3(level4_in[2877]),
   .I4(level4_in[2878]),
   .I5(level4_in[2879])
);

LUT6 #(
   .INIT(64'h78a936cd78a936cd)  
) LUT6_inst8256 (
   .O(to_level3[480]),
   .I0(level4_in[2880]),
   .I1(level4_in[2881]),
   .I2(level4_in[2882]),
   .I3(level4_in[2883]),
   .I4(level4_in[2884]),
   .I5(level4_in[2885])
);

LUT6 #(
   .INIT(64'ha8b000bea8b000be)  
) LUT6_inst8257 (
   .O(to_level3[481]),
   .I0(level4_in[2886]),
   .I1(level4_in[2887]),
   .I2(level4_in[2888]),
   .I3(level4_in[2889]),
   .I4(level4_in[2890]),
   .I5(level4_in[2891])
);

LUT6 #(
   .INIT(64'h66d94aad66d94aad)  
) LUT6_inst8258 (
   .O(to_level3[482]),
   .I0(level4_in[2892]),
   .I1(level4_in[2893]),
   .I2(level4_in[2894]),
   .I3(level4_in[2895]),
   .I4(level4_in[2896]),
   .I5(level4_in[2897])
);

LUT6 #(
   .INIT(64'he199f44ee199f44e)  
) LUT6_inst8259 (
   .O(to_level3[483]),
   .I0(level4_in[2898]),
   .I1(level4_in[2899]),
   .I2(level4_in[2900]),
   .I3(level4_in[2901]),
   .I4(level4_in[2902]),
   .I5(level4_in[2903])
);

LUT6 #(
   .INIT(64'hd3eb910ed3eb910e)  
) LUT6_inst8260 (
   .O(to_level3[484]),
   .I0(level4_in[2904]),
   .I1(level4_in[2905]),
   .I2(level4_in[2906]),
   .I3(level4_in[2907]),
   .I4(level4_in[2908]),
   .I5(level4_in[2909])
);

LUT6 #(
   .INIT(64'h51a2684e51a2684e)  
) LUT6_inst8261 (
   .O(to_level3[485]),
   .I0(level4_in[2910]),
   .I1(level4_in[2911]),
   .I2(level4_in[2912]),
   .I3(level4_in[2913]),
   .I4(level4_in[2914]),
   .I5(level4_in[2915])
);

LUT6 #(
   .INIT(64'h7a5b53797a5b5379)  
) LUT6_inst8262 (
   .O(to_level3[486]),
   .I0(level4_in[2916]),
   .I1(level4_in[2917]),
   .I2(level4_in[2918]),
   .I3(level4_in[2919]),
   .I4(level4_in[2920]),
   .I5(level4_in[2921])
);

LUT6 #(
   .INIT(64'h463c06fe463c06fe)  
) LUT6_inst8263 (
   .O(to_level3[487]),
   .I0(level4_in[2922]),
   .I1(level4_in[2923]),
   .I2(level4_in[2924]),
   .I3(level4_in[2925]),
   .I4(level4_in[2926]),
   .I5(level4_in[2927])
);

LUT6 #(
   .INIT(64'hcf1c6c06cf1c6c06)  
) LUT6_inst8264 (
   .O(to_level3[488]),
   .I0(level4_in[2928]),
   .I1(level4_in[2929]),
   .I2(level4_in[2930]),
   .I3(level4_in[2931]),
   .I4(level4_in[2932]),
   .I5(level4_in[2933])
);

LUT6 #(
   .INIT(64'hf19d089cf19d089c)  
) LUT6_inst8265 (
   .O(to_level3[489]),
   .I0(level4_in[2934]),
   .I1(level4_in[2935]),
   .I2(level4_in[2936]),
   .I3(level4_in[2937]),
   .I4(level4_in[2938]),
   .I5(level4_in[2939])
);

LUT6 #(
   .INIT(64'h287c6350287c6350)  
) LUT6_inst8266 (
   .O(to_level3[490]),
   .I0(level4_in[2940]),
   .I1(level4_in[2941]),
   .I2(level4_in[2942]),
   .I3(level4_in[2943]),
   .I4(level4_in[2944]),
   .I5(level4_in[2945])
);

LUT6 #(
   .INIT(64'h8312424483124244)  
) LUT6_inst8267 (
   .O(to_level3[491]),
   .I0(level4_in[2946]),
   .I1(level4_in[2947]),
   .I2(level4_in[2948]),
   .I3(level4_in[2949]),
   .I4(level4_in[2950]),
   .I5(level4_in[2951])
);

LUT6 #(
   .INIT(64'h48a7c8a348a7c8a3)  
) LUT6_inst8268 (
   .O(to_level3[492]),
   .I0(level4_in[2952]),
   .I1(level4_in[2953]),
   .I2(level4_in[2954]),
   .I3(level4_in[2955]),
   .I4(level4_in[2956]),
   .I5(level4_in[2957])
);

LUT6 #(
   .INIT(64'h7842deb27842deb2)  
) LUT6_inst8269 (
   .O(to_level3[493]),
   .I0(level4_in[2958]),
   .I1(level4_in[2959]),
   .I2(level4_in[2960]),
   .I3(level4_in[2961]),
   .I4(level4_in[2962]),
   .I5(level4_in[2963])
);

LUT6 #(
   .INIT(64'hba75fc11ba75fc11)  
) LUT6_inst8270 (
   .O(to_level3[494]),
   .I0(level4_in[2964]),
   .I1(level4_in[2965]),
   .I2(level4_in[2966]),
   .I3(level4_in[2967]),
   .I4(level4_in[2968]),
   .I5(level4_in[2969])
);

LUT6 #(
   .INIT(64'h4f1292c54f1292c5)  
) LUT6_inst8271 (
   .O(to_level3[495]),
   .I0(level4_in[2970]),
   .I1(level4_in[2971]),
   .I2(level4_in[2972]),
   .I3(level4_in[2973]),
   .I4(level4_in[2974]),
   .I5(level4_in[2975])
);

LUT6 #(
   .INIT(64'h979469b3979469b3)  
) LUT6_inst8272 (
   .O(to_level3[496]),
   .I0(level4_in[2976]),
   .I1(level4_in[2977]),
   .I2(level4_in[2978]),
   .I3(level4_in[2979]),
   .I4(level4_in[2980]),
   .I5(level4_in[2981])
);

LUT6 #(
   .INIT(64'hf4d0ade1f4d0ade1)  
) LUT6_inst8273 (
   .O(to_level3[497]),
   .I0(level4_in[2982]),
   .I1(level4_in[2983]),
   .I2(level4_in[2984]),
   .I3(level4_in[2985]),
   .I4(level4_in[2986]),
   .I5(level4_in[2987])
);

LUT6 #(
   .INIT(64'h64cee17d64cee17d)  
) LUT6_inst8274 (
   .O(to_level3[498]),
   .I0(level4_in[2988]),
   .I1(level4_in[2989]),
   .I2(level4_in[2990]),
   .I3(level4_in[2991]),
   .I4(level4_in[2992]),
   .I5(level4_in[2993])
);

LUT6 #(
   .INIT(64'h2b9f8f0c2b9f8f0c)  
) LUT6_inst8275 (
   .O(to_level3[499]),
   .I0(level4_in[2994]),
   .I1(level4_in[2995]),
   .I2(level4_in[2996]),
   .I3(level4_in[2997]),
   .I4(level4_in[2998]),
   .I5(level4_in[2999])
);

LUT6 #(
   .INIT(64'h3a1882bc3a1882bc)  
) LUT6_inst8276 (
   .O(to_level3[500]),
   .I0(level4_in[3000]),
   .I1(level4_in[3001]),
   .I2(level4_in[3002]),
   .I3(level4_in[3003]),
   .I4(level4_in[3004]),
   .I5(level4_in[3005])
);

LUT6 #(
   .INIT(64'hf8efe60bf8efe60b)  
) LUT6_inst8277 (
   .O(to_level3[501]),
   .I0(level4_in[3006]),
   .I1(level4_in[3007]),
   .I2(level4_in[3008]),
   .I3(level4_in[3009]),
   .I4(level4_in[3010]),
   .I5(level4_in[3011])
);

LUT6 #(
   .INIT(64'hc29af50dc29af50d)  
) LUT6_inst8278 (
   .O(to_level3[502]),
   .I0(level4_in[3012]),
   .I1(level4_in[3013]),
   .I2(level4_in[3014]),
   .I3(level4_in[3015]),
   .I4(level4_in[3016]),
   .I5(level4_in[3017])
);

LUT6 #(
   .INIT(64'h4c4933764c493376)  
) LUT6_inst8279 (
   .O(to_level3[503]),
   .I0(level4_in[3018]),
   .I1(level4_in[3019]),
   .I2(level4_in[3020]),
   .I3(level4_in[3021]),
   .I4(level4_in[3022]),
   .I5(level4_in[3023])
);

LUT6 #(
   .INIT(64'hbbf64658bbf64658)  
) LUT6_inst8280 (
   .O(to_level3[504]),
   .I0(level4_in[3024]),
   .I1(level4_in[3025]),
   .I2(level4_in[3026]),
   .I3(level4_in[3027]),
   .I4(level4_in[3028]),
   .I5(level4_in[3029])
);

LUT6 #(
   .INIT(64'hdf478a09df478a09)  
) LUT6_inst8281 (
   .O(to_level3[505]),
   .I0(level4_in[3030]),
   .I1(level4_in[3031]),
   .I2(level4_in[3032]),
   .I3(level4_in[3033]),
   .I4(level4_in[3034]),
   .I5(level4_in[3035])
);

LUT6 #(
   .INIT(64'h88477d4b88477d4b)  
) LUT6_inst8282 (
   .O(to_level3[506]),
   .I0(level4_in[3036]),
   .I1(level4_in[3037]),
   .I2(level4_in[3038]),
   .I3(level4_in[3039]),
   .I4(level4_in[3040]),
   .I5(level4_in[3041])
);

LUT6 #(
   .INIT(64'h856ea777856ea777)  
) LUT6_inst8283 (
   .O(to_level3[507]),
   .I0(level4_in[3042]),
   .I1(level4_in[3043]),
   .I2(level4_in[3044]),
   .I3(level4_in[3045]),
   .I4(level4_in[3046]),
   .I5(level4_in[3047])
);

LUT6 #(
   .INIT(64'hc9594904c9594904)  
) LUT6_inst8284 (
   .O(to_level3[508]),
   .I0(level4_in[3048]),
   .I1(level4_in[3049]),
   .I2(level4_in[3050]),
   .I3(level4_in[3051]),
   .I4(level4_in[3052]),
   .I5(level4_in[3053])
);

LUT6 #(
   .INIT(64'h4f6a5bc94f6a5bc9)  
) LUT6_inst8285 (
   .O(to_level3[509]),
   .I0(level4_in[3054]),
   .I1(level4_in[3055]),
   .I2(level4_in[3056]),
   .I3(level4_in[3057]),
   .I4(level4_in[3058]),
   .I5(level4_in[3059])
);

LUT6 #(
   .INIT(64'h64a26ca964a26ca9)  
) LUT6_inst8286 (
   .O(to_level3[510]),
   .I0(level4_in[3060]),
   .I1(level4_in[3061]),
   .I2(level4_in[3062]),
   .I3(level4_in[3063]),
   .I4(level4_in[3064]),
   .I5(level4_in[3065])
);

LUT6 #(
   .INIT(64'h4f6755554f675555)  
) LUT6_inst8287 (
   .O(to_level3[511]),
   .I0(level4_in[3066]),
   .I1(level4_in[3067]),
   .I2(level4_in[3068]),
   .I3(level4_in[3069]),
   .I4(level4_in[3070]),
   .I5(level4_in[3071])
);

LUT6 #(
   .INIT(64'h6ebdc1136ebdc113)  
) LUT6_inst8288 (
   .O(to_level3[512]),
   .I0(level4_in[3072]),
   .I1(level4_in[3073]),
   .I2(level4_in[3074]),
   .I3(level4_in[3075]),
   .I4(level4_in[3076]),
   .I5(level4_in[3077])
);

LUT6 #(
   .INIT(64'h15089dfb15089dfb)  
) LUT6_inst8289 (
   .O(to_level3[513]),
   .I0(level4_in[3078]),
   .I1(level4_in[3079]),
   .I2(level4_in[3080]),
   .I3(level4_in[3081]),
   .I4(level4_in[3082]),
   .I5(level4_in[3083])
);

LUT6 #(
   .INIT(64'h6a0479696a047969)  
) LUT6_inst8290 (
   .O(to_level3[514]),
   .I0(level4_in[3084]),
   .I1(level4_in[3085]),
   .I2(level4_in[3086]),
   .I3(level4_in[3087]),
   .I4(level4_in[3088]),
   .I5(level4_in[3089])
);

LUT6 #(
   .INIT(64'hca586a2dca586a2d)  
) LUT6_inst8291 (
   .O(to_level3[515]),
   .I0(level4_in[3090]),
   .I1(level4_in[3091]),
   .I2(level4_in[3092]),
   .I3(level4_in[3093]),
   .I4(level4_in[3094]),
   .I5(level4_in[3095])
);

LUT6 #(
   .INIT(64'h8c19d2db8c19d2db)  
) LUT6_inst8292 (
   .O(to_level3[516]),
   .I0(level4_in[3096]),
   .I1(level4_in[3097]),
   .I2(level4_in[3098]),
   .I3(level4_in[3099]),
   .I4(level4_in[3100]),
   .I5(level4_in[3101])
);

LUT6 #(
   .INIT(64'h365d5327365d5327)  
) LUT6_inst8293 (
   .O(to_level3[517]),
   .I0(level4_in[3102]),
   .I1(level4_in[3103]),
   .I2(level4_in[3104]),
   .I3(level4_in[3105]),
   .I4(level4_in[3106]),
   .I5(level4_in[3107])
);

LUT6 #(
   .INIT(64'h98e2e7d698e2e7d6)  
) LUT6_inst8294 (
   .O(to_level3[518]),
   .I0(level4_in[3108]),
   .I1(level4_in[3109]),
   .I2(level4_in[3110]),
   .I3(level4_in[3111]),
   .I4(level4_in[3112]),
   .I5(level4_in[3113])
);

LUT6 #(
   .INIT(64'hb095b10eb095b10e)  
) LUT6_inst8295 (
   .O(to_level3[519]),
   .I0(level4_in[3114]),
   .I1(level4_in[3115]),
   .I2(level4_in[3116]),
   .I3(level4_in[3117]),
   .I4(level4_in[3118]),
   .I5(level4_in[3119])
);

LUT6 #(
   .INIT(64'h6cc013776cc01377)  
) LUT6_inst8296 (
   .O(to_level3[520]),
   .I0(level4_in[3120]),
   .I1(level4_in[3121]),
   .I2(level4_in[3122]),
   .I3(level4_in[3123]),
   .I4(level4_in[3124]),
   .I5(level4_in[3125])
);

LUT6 #(
   .INIT(64'hc2d140e6c2d140e6)  
) LUT6_inst8297 (
   .O(to_level3[521]),
   .I0(level4_in[3126]),
   .I1(level4_in[3127]),
   .I2(level4_in[3128]),
   .I3(level4_in[3129]),
   .I4(level4_in[3130]),
   .I5(level4_in[3131])
);

LUT6 #(
   .INIT(64'h667cae1e667cae1e)  
) LUT6_inst8298 (
   .O(to_level3[522]),
   .I0(level4_in[3132]),
   .I1(level4_in[3133]),
   .I2(level4_in[3134]),
   .I3(level4_in[3135]),
   .I4(level4_in[3136]),
   .I5(level4_in[3137])
);

LUT6 #(
   .INIT(64'hb5dcc50db5dcc50d)  
) LUT6_inst8299 (
   .O(to_level3[523]),
   .I0(level4_in[3138]),
   .I1(level4_in[3139]),
   .I2(level4_in[3140]),
   .I3(level4_in[3141]),
   .I4(level4_in[3142]),
   .I5(level4_in[3143])
);

LUT6 #(
   .INIT(64'h5171c9095171c909)  
) LUT6_inst8300 (
   .O(to_level3[524]),
   .I0(level4_in[3144]),
   .I1(level4_in[3145]),
   .I2(level4_in[3146]),
   .I3(level4_in[3147]),
   .I4(level4_in[3148]),
   .I5(level4_in[3149])
);

LUT6 #(
   .INIT(64'h0e99bab70e99bab7)  
) LUT6_inst8301 (
   .O(to_level3[525]),
   .I0(level4_in[3150]),
   .I1(level4_in[3151]),
   .I2(level4_in[3152]),
   .I3(level4_in[3153]),
   .I4(level4_in[3154]),
   .I5(level4_in[3155])
);

LUT6 #(
   .INIT(64'h2112632121126321)  
) LUT6_inst8302 (
   .O(to_level3[526]),
   .I0(level4_in[3156]),
   .I1(level4_in[3157]),
   .I2(level4_in[3158]),
   .I3(level4_in[3159]),
   .I4(level4_in[3160]),
   .I5(level4_in[3161])
);

LUT6 #(
   .INIT(64'h9468c4e49468c4e4)  
) LUT6_inst8303 (
   .O(to_level3[527]),
   .I0(level4_in[3162]),
   .I1(level4_in[3163]),
   .I2(level4_in[3164]),
   .I3(level4_in[3165]),
   .I4(level4_in[3166]),
   .I5(level4_in[3167])
);

LUT6 #(
   .INIT(64'hf769da83f769da83)  
) LUT6_inst8304 (
   .O(to_level3[528]),
   .I0(level4_in[3168]),
   .I1(level4_in[3169]),
   .I2(level4_in[3170]),
   .I3(level4_in[3171]),
   .I4(level4_in[3172]),
   .I5(level4_in[3173])
);

LUT6 #(
   .INIT(64'h8bf6a4ee8bf6a4ee)  
) LUT6_inst8305 (
   .O(to_level3[529]),
   .I0(level4_in[3174]),
   .I1(level4_in[3175]),
   .I2(level4_in[3176]),
   .I3(level4_in[3177]),
   .I4(level4_in[3178]),
   .I5(level4_in[3179])
);

LUT6 #(
   .INIT(64'h71ae6e0871ae6e08)  
) LUT6_inst8306 (
   .O(to_level3[530]),
   .I0(level4_in[3180]),
   .I1(level4_in[3181]),
   .I2(level4_in[3182]),
   .I3(level4_in[3183]),
   .I4(level4_in[3184]),
   .I5(level4_in[3185])
);

LUT6 #(
   .INIT(64'h6fb17a906fb17a90)  
) LUT6_inst8307 (
   .O(to_level3[531]),
   .I0(level4_in[3186]),
   .I1(level4_in[3187]),
   .I2(level4_in[3188]),
   .I3(level4_in[3189]),
   .I4(level4_in[3190]),
   .I5(level4_in[3191])
);

LUT6 #(
   .INIT(64'hd121e0d0d121e0d0)  
) LUT6_inst8308 (
   .O(to_level3[532]),
   .I0(level4_in[3192]),
   .I1(level4_in[3193]),
   .I2(level4_in[3194]),
   .I3(level4_in[3195]),
   .I4(level4_in[3196]),
   .I5(level4_in[3197])
);

LUT6 #(
   .INIT(64'hbfb6a4a3bfb6a4a3)  
) LUT6_inst8309 (
   .O(to_level3[533]),
   .I0(level4_in[3198]),
   .I1(level4_in[3199]),
   .I2(level4_in[3200]),
   .I3(level4_in[3201]),
   .I4(level4_in[3202]),
   .I5(level4_in[3203])
);

LUT6 #(
   .INIT(64'h1676878c1676878c)  
) LUT6_inst8310 (
   .O(to_level3[534]),
   .I0(level4_in[3204]),
   .I1(level4_in[3205]),
   .I2(level4_in[3206]),
   .I3(level4_in[3207]),
   .I4(level4_in[3208]),
   .I5(level4_in[3209])
);

LUT6 #(
   .INIT(64'h53eb56b453eb56b4)  
) LUT6_inst8311 (
   .O(to_level3[535]),
   .I0(level4_in[3210]),
   .I1(level4_in[3211]),
   .I2(level4_in[3212]),
   .I3(level4_in[3213]),
   .I4(level4_in[3214]),
   .I5(level4_in[3215])
);

LUT6 #(
   .INIT(64'hebae30dbebae30db)  
) LUT6_inst8312 (
   .O(to_level3[536]),
   .I0(level4_in[3216]),
   .I1(level4_in[3217]),
   .I2(level4_in[3218]),
   .I3(level4_in[3219]),
   .I4(level4_in[3220]),
   .I5(level4_in[3221])
);

LUT6 #(
   .INIT(64'h5b1521325b152132)  
) LUT6_inst8313 (
   .O(to_level3[537]),
   .I0(level4_in[3222]),
   .I1(level4_in[3223]),
   .I2(level4_in[3224]),
   .I3(level4_in[3225]),
   .I4(level4_in[3226]),
   .I5(level4_in[3227])
);

LUT6 #(
   .INIT(64'hf93f645ef93f645e)  
) LUT6_inst8314 (
   .O(to_level3[538]),
   .I0(level4_in[3228]),
   .I1(level4_in[3229]),
   .I2(level4_in[3230]),
   .I3(level4_in[3231]),
   .I4(level4_in[3232]),
   .I5(level4_in[3233])
);

LUT6 #(
   .INIT(64'hb54684d6b54684d6)  
) LUT6_inst8315 (
   .O(to_level3[539]),
   .I0(level4_in[3234]),
   .I1(level4_in[3235]),
   .I2(level4_in[3236]),
   .I3(level4_in[3237]),
   .I4(level4_in[3238]),
   .I5(level4_in[3239])
);

LUT6 #(
   .INIT(64'h0a42a3380a42a338)  
) LUT6_inst8316 (
   .O(to_level3[540]),
   .I0(level4_in[3240]),
   .I1(level4_in[3241]),
   .I2(level4_in[3242]),
   .I3(level4_in[3243]),
   .I4(level4_in[3244]),
   .I5(level4_in[3245])
);

LUT6 #(
   .INIT(64'h68a8f09c68a8f09c)  
) LUT6_inst8317 (
   .O(to_level3[541]),
   .I0(level4_in[3246]),
   .I1(level4_in[3247]),
   .I2(level4_in[3248]),
   .I3(level4_in[3249]),
   .I4(level4_in[3250]),
   .I5(level4_in[3251])
);

LUT6 #(
   .INIT(64'h1be84e421be84e42)  
) LUT6_inst8318 (
   .O(to_level3[542]),
   .I0(level4_in[3252]),
   .I1(level4_in[3253]),
   .I2(level4_in[3254]),
   .I3(level4_in[3255]),
   .I4(level4_in[3256]),
   .I5(level4_in[3257])
);

LUT6 #(
   .INIT(64'he1b1c491e1b1c491)  
) LUT6_inst8319 (
   .O(to_level3[543]),
   .I0(level4_in[3258]),
   .I1(level4_in[3259]),
   .I2(level4_in[3260]),
   .I3(level4_in[3261]),
   .I4(level4_in[3262]),
   .I5(level4_in[3263])
);

LUT6 #(
   .INIT(64'h6bdad28c6bdad28c)  
) LUT6_inst8320 (
   .O(to_level3[544]),
   .I0(level4_in[3264]),
   .I1(level4_in[3265]),
   .I2(level4_in[3266]),
   .I3(level4_in[3267]),
   .I4(level4_in[3268]),
   .I5(level4_in[3269])
);

LUT6 #(
   .INIT(64'hf773b8b8f773b8b8)  
) LUT6_inst8321 (
   .O(to_level3[545]),
   .I0(level4_in[3270]),
   .I1(level4_in[3271]),
   .I2(level4_in[3272]),
   .I3(level4_in[3273]),
   .I4(level4_in[3274]),
   .I5(level4_in[3275])
);

LUT6 #(
   .INIT(64'hc31e00d0c31e00d0)  
) LUT6_inst8322 (
   .O(to_level3[546]),
   .I0(level4_in[3276]),
   .I1(level4_in[3277]),
   .I2(level4_in[3278]),
   .I3(level4_in[3279]),
   .I4(level4_in[3280]),
   .I5(level4_in[3281])
);

LUT6 #(
   .INIT(64'hbc649556bc649556)  
) LUT6_inst8323 (
   .O(to_level3[547]),
   .I0(level4_in[3282]),
   .I1(level4_in[3283]),
   .I2(level4_in[3284]),
   .I3(level4_in[3285]),
   .I4(level4_in[3286]),
   .I5(level4_in[3287])
);

LUT6 #(
   .INIT(64'h6393f7536393f753)  
) LUT6_inst8324 (
   .O(to_level3[548]),
   .I0(level4_in[3288]),
   .I1(level4_in[3289]),
   .I2(level4_in[3290]),
   .I3(level4_in[3291]),
   .I4(level4_in[3292]),
   .I5(level4_in[3293])
);

LUT6 #(
   .INIT(64'h12e7c09d12e7c09d)  
) LUT6_inst8325 (
   .O(to_level3[549]),
   .I0(level4_in[3294]),
   .I1(level4_in[3295]),
   .I2(level4_in[3296]),
   .I3(level4_in[3297]),
   .I4(level4_in[3298]),
   .I5(level4_in[3299])
);

LUT6 #(
   .INIT(64'h56ab317656ab3176)  
) LUT6_inst8326 (
   .O(to_level3[550]),
   .I0(level4_in[3300]),
   .I1(level4_in[3301]),
   .I2(level4_in[3302]),
   .I3(level4_in[3303]),
   .I4(level4_in[3304]),
   .I5(level4_in[3305])
);

LUT6 #(
   .INIT(64'hc6f60678c6f60678)  
) LUT6_inst8327 (
   .O(to_level3[551]),
   .I0(level4_in[3306]),
   .I1(level4_in[3307]),
   .I2(level4_in[3308]),
   .I3(level4_in[3309]),
   .I4(level4_in[3310]),
   .I5(level4_in[3311])
);

LUT6 #(
   .INIT(64'h51f3fa0b51f3fa0b)  
) LUT6_inst8328 (
   .O(to_level3[552]),
   .I0(level4_in[3312]),
   .I1(level4_in[3313]),
   .I2(level4_in[3314]),
   .I3(level4_in[3315]),
   .I4(level4_in[3316]),
   .I5(level4_in[3317])
);

LUT6 #(
   .INIT(64'h4bcef1ed4bcef1ed)  
) LUT6_inst8329 (
   .O(to_level3[553]),
   .I0(level4_in[3318]),
   .I1(level4_in[3319]),
   .I2(level4_in[3320]),
   .I3(level4_in[3321]),
   .I4(level4_in[3322]),
   .I5(level4_in[3323])
);

LUT6 #(
   .INIT(64'h4dd21b854dd21b85)  
) LUT6_inst8330 (
   .O(to_level3[554]),
   .I0(level4_in[3324]),
   .I1(level4_in[3325]),
   .I2(level4_in[3326]),
   .I3(level4_in[3327]),
   .I4(level4_in[3328]),
   .I5(level4_in[3329])
);

LUT6 #(
   .INIT(64'h2479d7102479d710)  
) LUT6_inst8331 (
   .O(to_level3[555]),
   .I0(level4_in[3330]),
   .I1(level4_in[3331]),
   .I2(level4_in[3332]),
   .I3(level4_in[3333]),
   .I4(level4_in[3334]),
   .I5(level4_in[3335])
);

LUT6 #(
   .INIT(64'hfc1e5608fc1e5608)  
) LUT6_inst8332 (
   .O(to_level3[556]),
   .I0(level4_in[3336]),
   .I1(level4_in[3337]),
   .I2(level4_in[3338]),
   .I3(level4_in[3339]),
   .I4(level4_in[3340]),
   .I5(level4_in[3341])
);

LUT6 #(
   .INIT(64'h0d54d2580d54d258)  
) LUT6_inst8333 (
   .O(to_level3[557]),
   .I0(level4_in[3342]),
   .I1(level4_in[3343]),
   .I2(level4_in[3344]),
   .I3(level4_in[3345]),
   .I4(level4_in[3346]),
   .I5(level4_in[3347])
);

LUT6 #(
   .INIT(64'h6a687b736a687b73)  
) LUT6_inst8334 (
   .O(to_level3[558]),
   .I0(level4_in[3348]),
   .I1(level4_in[3349]),
   .I2(level4_in[3350]),
   .I3(level4_in[3351]),
   .I4(level4_in[3352]),
   .I5(level4_in[3353])
);

LUT6 #(
   .INIT(64'he63d5a6be63d5a6b)  
) LUT6_inst8335 (
   .O(to_level3[559]),
   .I0(level4_in[3354]),
   .I1(level4_in[3355]),
   .I2(level4_in[3356]),
   .I3(level4_in[3357]),
   .I4(level4_in[3358]),
   .I5(level4_in[3359])
);

LUT6 #(
   .INIT(64'hf2544684f2544684)  
) LUT6_inst8336 (
   .O(to_level3[560]),
   .I0(level4_in[3360]),
   .I1(level4_in[3361]),
   .I2(level4_in[3362]),
   .I3(level4_in[3363]),
   .I4(level4_in[3364]),
   .I5(level4_in[3365])
);

LUT6 #(
   .INIT(64'h0b4ccd870b4ccd87)  
) LUT6_inst8337 (
   .O(to_level3[561]),
   .I0(level4_in[3366]),
   .I1(level4_in[3367]),
   .I2(level4_in[3368]),
   .I3(level4_in[3369]),
   .I4(level4_in[3370]),
   .I5(level4_in[3371])
);

LUT6 #(
   .INIT(64'h7a89d94a7a89d94a)  
) LUT6_inst8338 (
   .O(to_level3[562]),
   .I0(level4_in[3372]),
   .I1(level4_in[3373]),
   .I2(level4_in[3374]),
   .I3(level4_in[3375]),
   .I4(level4_in[3376]),
   .I5(level4_in[3377])
);

LUT6 #(
   .INIT(64'h433dbe8c433dbe8c)  
) LUT6_inst8339 (
   .O(to_level3[563]),
   .I0(level4_in[3378]),
   .I1(level4_in[3379]),
   .I2(level4_in[3380]),
   .I3(level4_in[3381]),
   .I4(level4_in[3382]),
   .I5(level4_in[3383])
);

LUT6 #(
   .INIT(64'h4c9395bb4c9395bb)  
) LUT6_inst8340 (
   .O(to_level3[564]),
   .I0(level4_in[3384]),
   .I1(level4_in[3385]),
   .I2(level4_in[3386]),
   .I3(level4_in[3387]),
   .I4(level4_in[3388]),
   .I5(level4_in[3389])
);

LUT6 #(
   .INIT(64'h02897bf602897bf6)  
) LUT6_inst8341 (
   .O(to_level3[565]),
   .I0(level4_in[3390]),
   .I1(level4_in[3391]),
   .I2(level4_in[3392]),
   .I3(level4_in[3393]),
   .I4(level4_in[3394]),
   .I5(level4_in[3395])
);

LUT6 #(
   .INIT(64'h7092623b7092623b)  
) LUT6_inst8342 (
   .O(to_level3[566]),
   .I0(level4_in[3396]),
   .I1(level4_in[3397]),
   .I2(level4_in[3398]),
   .I3(level4_in[3399]),
   .I4(level4_in[3400]),
   .I5(level4_in[3401])
);

LUT6 #(
   .INIT(64'haa91a748aa91a748)  
) LUT6_inst8343 (
   .O(to_level3[567]),
   .I0(level4_in[3402]),
   .I1(level4_in[3403]),
   .I2(level4_in[3404]),
   .I3(level4_in[3405]),
   .I4(level4_in[3406]),
   .I5(level4_in[3407])
);

LUT6 #(
   .INIT(64'hf8f3de9df8f3de9d)  
) LUT6_inst8344 (
   .O(to_level3[568]),
   .I0(level4_in[3408]),
   .I1(level4_in[3409]),
   .I2(level4_in[3410]),
   .I3(level4_in[3411]),
   .I4(level4_in[3412]),
   .I5(level4_in[3413])
);

LUT6 #(
   .INIT(64'h24a9a50524a9a505)  
) LUT6_inst8345 (
   .O(to_level3[569]),
   .I0(level4_in[3414]),
   .I1(level4_in[3415]),
   .I2(level4_in[3416]),
   .I3(level4_in[3417]),
   .I4(level4_in[3418]),
   .I5(level4_in[3419])
);

LUT6 #(
   .INIT(64'h9999123899991238)  
) LUT6_inst8346 (
   .O(to_level3[570]),
   .I0(level4_in[3420]),
   .I1(level4_in[3421]),
   .I2(level4_in[3422]),
   .I3(level4_in[3423]),
   .I4(level4_in[3424]),
   .I5(level4_in[3425])
);

LUT6 #(
   .INIT(64'hb51f85aab51f85aa)  
) LUT6_inst8347 (
   .O(to_level3[571]),
   .I0(level4_in[3426]),
   .I1(level4_in[3427]),
   .I2(level4_in[3428]),
   .I3(level4_in[3429]),
   .I4(level4_in[3430]),
   .I5(level4_in[3431])
);

LUT6 #(
   .INIT(64'h412a3f12412a3f12)  
) LUT6_inst8348 (
   .O(to_level3[572]),
   .I0(level4_in[3432]),
   .I1(level4_in[3433]),
   .I2(level4_in[3434]),
   .I3(level4_in[3435]),
   .I4(level4_in[3436]),
   .I5(level4_in[3437])
);

LUT6 #(
   .INIT(64'h8f7767098f776709)  
) LUT6_inst8349 (
   .O(to_level3[573]),
   .I0(level4_in[3438]),
   .I1(level4_in[3439]),
   .I2(level4_in[3440]),
   .I3(level4_in[3441]),
   .I4(level4_in[3442]),
   .I5(level4_in[3443])
);

LUT6 #(
   .INIT(64'h29e4452a29e4452a)  
) LUT6_inst8350 (
   .O(to_level3[574]),
   .I0(level4_in[3444]),
   .I1(level4_in[3445]),
   .I2(level4_in[3446]),
   .I3(level4_in[3447]),
   .I4(level4_in[3448]),
   .I5(level4_in[3449])
);

LUT6 #(
   .INIT(64'h15a65b5215a65b52)  
) LUT6_inst8351 (
   .O(to_level3[575]),
   .I0(level4_in[3450]),
   .I1(level4_in[3451]),
   .I2(level4_in[3452]),
   .I3(level4_in[3453]),
   .I4(level4_in[3454]),
   .I5(level4_in[3455])
);

LUT6 #(
   .INIT(64'ha72a7223a72a7223)  
) LUT6_inst8352 (
   .O(to_level3[576]),
   .I0(level4_in[3456]),
   .I1(level4_in[3457]),
   .I2(level4_in[3458]),
   .I3(level4_in[3459]),
   .I4(level4_in[3460]),
   .I5(level4_in[3461])
);

LUT6 #(
   .INIT(64'h592b9a4c592b9a4c)  
) LUT6_inst8353 (
   .O(to_level3[577]),
   .I0(level4_in[3462]),
   .I1(level4_in[3463]),
   .I2(level4_in[3464]),
   .I3(level4_in[3465]),
   .I4(level4_in[3466]),
   .I5(level4_in[3467])
);

LUT6 #(
   .INIT(64'hae3128fdae3128fd)  
) LUT6_inst8354 (
   .O(to_level3[578]),
   .I0(level4_in[3468]),
   .I1(level4_in[3469]),
   .I2(level4_in[3470]),
   .I3(level4_in[3471]),
   .I4(level4_in[3472]),
   .I5(level4_in[3473])
);

LUT6 #(
   .INIT(64'hb3e6cd02b3e6cd02)  
) LUT6_inst8355 (
   .O(to_level3[579]),
   .I0(level4_in[3474]),
   .I1(level4_in[3475]),
   .I2(level4_in[3476]),
   .I3(level4_in[3477]),
   .I4(level4_in[3478]),
   .I5(level4_in[3479])
);

LUT6 #(
   .INIT(64'h9473179f9473179f)  
) LUT6_inst8356 (
   .O(to_level3[580]),
   .I0(level4_in[3480]),
   .I1(level4_in[3481]),
   .I2(level4_in[3482]),
   .I3(level4_in[3483]),
   .I4(level4_in[3484]),
   .I5(level4_in[3485])
);

LUT6 #(
   .INIT(64'h3e88cacc3e88cacc)  
) LUT6_inst8357 (
   .O(to_level3[581]),
   .I0(level4_in[3486]),
   .I1(level4_in[3487]),
   .I2(level4_in[3488]),
   .I3(level4_in[3489]),
   .I4(level4_in[3490]),
   .I5(level4_in[3491])
);

LUT6 #(
   .INIT(64'haeaf7942aeaf7942)  
) LUT6_inst8358 (
   .O(to_level3[582]),
   .I0(level4_in[3492]),
   .I1(level4_in[3493]),
   .I2(level4_in[3494]),
   .I3(level4_in[3495]),
   .I4(level4_in[3496]),
   .I5(level4_in[3497])
);

LUT6 #(
   .INIT(64'ha1882e44a1882e44)  
) LUT6_inst8359 (
   .O(to_level3[583]),
   .I0(level4_in[3498]),
   .I1(level4_in[3499]),
   .I2(level4_in[3500]),
   .I3(level4_in[3501]),
   .I4(level4_in[3502]),
   .I5(level4_in[3503])
);

LUT6 #(
   .INIT(64'hd9d03aead9d03aea)  
) LUT6_inst8360 (
   .O(to_level3[584]),
   .I0(level4_in[3504]),
   .I1(level4_in[3505]),
   .I2(level4_in[3506]),
   .I3(level4_in[3507]),
   .I4(level4_in[3508]),
   .I5(level4_in[3509])
);

LUT6 #(
   .INIT(64'ha68f149aa68f149a)  
) LUT6_inst8361 (
   .O(to_level3[585]),
   .I0(level4_in[3510]),
   .I1(level4_in[3511]),
   .I2(level4_in[3512]),
   .I3(level4_in[3513]),
   .I4(level4_in[3514]),
   .I5(level4_in[3515])
);

LUT6 #(
   .INIT(64'h07c7c5c007c7c5c0)  
) LUT6_inst8362 (
   .O(to_level3[586]),
   .I0(level4_in[3516]),
   .I1(level4_in[3517]),
   .I2(level4_in[3518]),
   .I3(level4_in[3519]),
   .I4(level4_in[3520]),
   .I5(level4_in[3521])
);

LUT6 #(
   .INIT(64'h09f382a509f382a5)  
) LUT6_inst8363 (
   .O(to_level3[587]),
   .I0(level4_in[3522]),
   .I1(level4_in[3523]),
   .I2(level4_in[3524]),
   .I3(level4_in[3525]),
   .I4(level4_in[3526]),
   .I5(level4_in[3527])
);

LUT6 #(
   .INIT(64'h32a8aaec32a8aaec)  
) LUT6_inst8364 (
   .O(to_level3[588]),
   .I0(level4_in[3528]),
   .I1(level4_in[3529]),
   .I2(level4_in[3530]),
   .I3(level4_in[3531]),
   .I4(level4_in[3532]),
   .I5(level4_in[3533])
);

LUT6 #(
   .INIT(64'h7fbd62bf7fbd62bf)  
) LUT6_inst8365 (
   .O(to_level3[589]),
   .I0(level4_in[3534]),
   .I1(level4_in[3535]),
   .I2(level4_in[3536]),
   .I3(level4_in[3537]),
   .I4(level4_in[3538]),
   .I5(level4_in[3539])
);

LUT6 #(
   .INIT(64'h909f2b0f909f2b0f)  
) LUT6_inst8366 (
   .O(to_level3[590]),
   .I0(level4_in[3540]),
   .I1(level4_in[3541]),
   .I2(level4_in[3542]),
   .I3(level4_in[3543]),
   .I4(level4_in[3544]),
   .I5(level4_in[3545])
);

LUT6 #(
   .INIT(64'h30da8d6430da8d64)  
) LUT6_inst8367 (
   .O(to_level3[591]),
   .I0(level4_in[3546]),
   .I1(level4_in[3547]),
   .I2(level4_in[3548]),
   .I3(level4_in[3549]),
   .I4(level4_in[3550]),
   .I5(level4_in[3551])
);

LUT6 #(
   .INIT(64'hb280c5e0b280c5e0)  
) LUT6_inst8368 (
   .O(to_level3[592]),
   .I0(level4_in[3552]),
   .I1(level4_in[3553]),
   .I2(level4_in[3554]),
   .I3(level4_in[3555]),
   .I4(level4_in[3556]),
   .I5(level4_in[3557])
);

LUT6 #(
   .INIT(64'ha0ec23e6a0ec23e6)  
) LUT6_inst8369 (
   .O(to_level3[593]),
   .I0(level4_in[3558]),
   .I1(level4_in[3559]),
   .I2(level4_in[3560]),
   .I3(level4_in[3561]),
   .I4(level4_in[3562]),
   .I5(level4_in[3563])
);

LUT6 #(
   .INIT(64'h886a5a50886a5a50)  
) LUT6_inst8370 (
   .O(to_level3[594]),
   .I0(level4_in[3564]),
   .I1(level4_in[3565]),
   .I2(level4_in[3566]),
   .I3(level4_in[3567]),
   .I4(level4_in[3568]),
   .I5(level4_in[3569])
);

LUT6 #(
   .INIT(64'hcf2c86f9cf2c86f9)  
) LUT6_inst8371 (
   .O(to_level3[595]),
   .I0(level4_in[3570]),
   .I1(level4_in[3571]),
   .I2(level4_in[3572]),
   .I3(level4_in[3573]),
   .I4(level4_in[3574]),
   .I5(level4_in[3575])
);

LUT6 #(
   .INIT(64'h9478cb689478cb68)  
) LUT6_inst8372 (
   .O(to_level3[596]),
   .I0(level4_in[3576]),
   .I1(level4_in[3577]),
   .I2(level4_in[3578]),
   .I3(level4_in[3579]),
   .I4(level4_in[3580]),
   .I5(level4_in[3581])
);

LUT6 #(
   .INIT(64'h3a70730e3a70730e)  
) LUT6_inst8373 (
   .O(to_level3[597]),
   .I0(level4_in[3582]),
   .I1(level4_in[3583]),
   .I2(level4_in[3584]),
   .I3(level4_in[3585]),
   .I4(level4_in[3586]),
   .I5(level4_in[3587])
);

LUT6 #(
   .INIT(64'h1806c2331806c233)  
) LUT6_inst8374 (
   .O(to_level3[598]),
   .I0(level4_in[3588]),
   .I1(level4_in[3589]),
   .I2(level4_in[3590]),
   .I3(level4_in[3591]),
   .I4(level4_in[3592]),
   .I5(level4_in[3593])
);

LUT6 #(
   .INIT(64'h4b96607c4b96607c)  
) LUT6_inst8375 (
   .O(to_level3[599]),
   .I0(level4_in[3594]),
   .I1(level4_in[3595]),
   .I2(level4_in[3596]),
   .I3(level4_in[3597]),
   .I4(level4_in[3598]),
   .I5(level4_in[3599])
);

LUT6 #(
   .INIT(64'h1dfe6ba91dfe6ba9)  
) LUT6_inst8376 (
   .O(to_level3[600]),
   .I0(level4_in[3600]),
   .I1(level4_in[3601]),
   .I2(level4_in[3602]),
   .I3(level4_in[3603]),
   .I4(level4_in[3604]),
   .I5(level4_in[3605])
);

LUT6 #(
   .INIT(64'h631d31ac631d31ac)  
) LUT6_inst8377 (
   .O(to_level3[601]),
   .I0(level4_in[3606]),
   .I1(level4_in[3607]),
   .I2(level4_in[3608]),
   .I3(level4_in[3609]),
   .I4(level4_in[3610]),
   .I5(level4_in[3611])
);

LUT6 #(
   .INIT(64'ha0a092e3a0a092e3)  
) LUT6_inst8378 (
   .O(to_level3[602]),
   .I0(level4_in[3612]),
   .I1(level4_in[3613]),
   .I2(level4_in[3614]),
   .I3(level4_in[3615]),
   .I4(level4_in[3616]),
   .I5(level4_in[3617])
);

LUT6 #(
   .INIT(64'ha1d1c40ea1d1c40e)  
) LUT6_inst8379 (
   .O(to_level3[603]),
   .I0(level4_in[3618]),
   .I1(level4_in[3619]),
   .I2(level4_in[3620]),
   .I3(level4_in[3621]),
   .I4(level4_in[3622]),
   .I5(level4_in[3623])
);

LUT6 #(
   .INIT(64'hc9fc06edc9fc06ed)  
) LUT6_inst8380 (
   .O(to_level3[604]),
   .I0(level4_in[3624]),
   .I1(level4_in[3625]),
   .I2(level4_in[3626]),
   .I3(level4_in[3627]),
   .I4(level4_in[3628]),
   .I5(level4_in[3629])
);

LUT6 #(
   .INIT(64'haed2ca59aed2ca59)  
) LUT6_inst8381 (
   .O(to_level3[605]),
   .I0(level4_in[3630]),
   .I1(level4_in[3631]),
   .I2(level4_in[3632]),
   .I3(level4_in[3633]),
   .I4(level4_in[3634]),
   .I5(level4_in[3635])
);

LUT6 #(
   .INIT(64'hc8ce7b7ac8ce7b7a)  
) LUT6_inst8382 (
   .O(to_level3[606]),
   .I0(level4_in[3636]),
   .I1(level4_in[3637]),
   .I2(level4_in[3638]),
   .I3(level4_in[3639]),
   .I4(level4_in[3640]),
   .I5(level4_in[3641])
);

LUT6 #(
   .INIT(64'hd661f6a1d661f6a1)  
) LUT6_inst8383 (
   .O(to_level3[607]),
   .I0(level4_in[3642]),
   .I1(level4_in[3643]),
   .I2(level4_in[3644]),
   .I3(level4_in[3645]),
   .I4(level4_in[3646]),
   .I5(level4_in[3647])
);

LUT6 #(
   .INIT(64'h4db8bc324db8bc32)  
) LUT6_inst8384 (
   .O(to_level3[608]),
   .I0(level4_in[3648]),
   .I1(level4_in[3649]),
   .I2(level4_in[3650]),
   .I3(level4_in[3651]),
   .I4(level4_in[3652]),
   .I5(level4_in[3653])
);

LUT6 #(
   .INIT(64'h74494e9374494e93)  
) LUT6_inst8385 (
   .O(to_level3[609]),
   .I0(level4_in[3654]),
   .I1(level4_in[3655]),
   .I2(level4_in[3656]),
   .I3(level4_in[3657]),
   .I4(level4_in[3658]),
   .I5(level4_in[3659])
);

LUT6 #(
   .INIT(64'h3377dd093377dd09)  
) LUT6_inst8386 (
   .O(to_level3[610]),
   .I0(level4_in[3660]),
   .I1(level4_in[3661]),
   .I2(level4_in[3662]),
   .I3(level4_in[3663]),
   .I4(level4_in[3664]),
   .I5(level4_in[3665])
);

LUT6 #(
   .INIT(64'hf7e9ee4df7e9ee4d)  
) LUT6_inst8387 (
   .O(to_level3[611]),
   .I0(level4_in[3666]),
   .I1(level4_in[3667]),
   .I2(level4_in[3668]),
   .I3(level4_in[3669]),
   .I4(level4_in[3670]),
   .I5(level4_in[3671])
);

LUT6 #(
   .INIT(64'h57d43ebb57d43ebb)  
) LUT6_inst8388 (
   .O(to_level3[612]),
   .I0(level4_in[3672]),
   .I1(level4_in[3673]),
   .I2(level4_in[3674]),
   .I3(level4_in[3675]),
   .I4(level4_in[3676]),
   .I5(level4_in[3677])
);

LUT6 #(
   .INIT(64'ha54c8ccca54c8ccc)  
) LUT6_inst8389 (
   .O(to_level3[613]),
   .I0(level4_in[3678]),
   .I1(level4_in[3679]),
   .I2(level4_in[3680]),
   .I3(level4_in[3681]),
   .I4(level4_in[3682]),
   .I5(level4_in[3683])
);

LUT6 #(
   .INIT(64'hd91abb85d91abb85)  
) LUT6_inst8390 (
   .O(to_level3[614]),
   .I0(level4_in[3684]),
   .I1(level4_in[3685]),
   .I2(level4_in[3686]),
   .I3(level4_in[3687]),
   .I4(level4_in[3688]),
   .I5(level4_in[3689])
);

LUT6 #(
   .INIT(64'h5b6634cf5b6634cf)  
) LUT6_inst8391 (
   .O(to_level3[615]),
   .I0(level4_in[3690]),
   .I1(level4_in[3691]),
   .I2(level4_in[3692]),
   .I3(level4_in[3693]),
   .I4(level4_in[3694]),
   .I5(level4_in[3695])
);

LUT6 #(
   .INIT(64'hed90ef30ed90ef30)  
) LUT6_inst8392 (
   .O(to_level3[616]),
   .I0(level4_in[3696]),
   .I1(level4_in[3697]),
   .I2(level4_in[3698]),
   .I3(level4_in[3699]),
   .I4(level4_in[3700]),
   .I5(level4_in[3701])
);

LUT6 #(
   .INIT(64'hfd2ed329fd2ed329)  
) LUT6_inst8393 (
   .O(to_level3[617]),
   .I0(level4_in[3702]),
   .I1(level4_in[3703]),
   .I2(level4_in[3704]),
   .I3(level4_in[3705]),
   .I4(level4_in[3706]),
   .I5(level4_in[3707])
);

LUT6 #(
   .INIT(64'hae66e5f9ae66e5f9)  
) LUT6_inst8394 (
   .O(to_level3[618]),
   .I0(level4_in[3708]),
   .I1(level4_in[3709]),
   .I2(level4_in[3710]),
   .I3(level4_in[3711]),
   .I4(level4_in[3712]),
   .I5(level4_in[3713])
);

LUT6 #(
   .INIT(64'h6f841fc66f841fc6)  
) LUT6_inst8395 (
   .O(to_level3[619]),
   .I0(level4_in[3714]),
   .I1(level4_in[3715]),
   .I2(level4_in[3716]),
   .I3(level4_in[3717]),
   .I4(level4_in[3718]),
   .I5(level4_in[3719])
);

LUT6 #(
   .INIT(64'h3e49c0ac3e49c0ac)  
) LUT6_inst8396 (
   .O(to_level3[620]),
   .I0(level4_in[3720]),
   .I1(level4_in[3721]),
   .I2(level4_in[3722]),
   .I3(level4_in[3723]),
   .I4(level4_in[3724]),
   .I5(level4_in[3725])
);

LUT6 #(
   .INIT(64'h8eb064e78eb064e7)  
) LUT6_inst8397 (
   .O(to_level3[621]),
   .I0(level4_in[3726]),
   .I1(level4_in[3727]),
   .I2(level4_in[3728]),
   .I3(level4_in[3729]),
   .I4(level4_in[3730]),
   .I5(level4_in[3731])
);

LUT6 #(
   .INIT(64'hecb4a001ecb4a001)  
) LUT6_inst8398 (
   .O(to_level3[622]),
   .I0(level4_in[3732]),
   .I1(level4_in[3733]),
   .I2(level4_in[3734]),
   .I3(level4_in[3735]),
   .I4(level4_in[3736]),
   .I5(level4_in[3737])
);

LUT6 #(
   .INIT(64'hbb397909bb397909)  
) LUT6_inst8399 (
   .O(to_level3[623]),
   .I0(level4_in[3738]),
   .I1(level4_in[3739]),
   .I2(level4_in[3740]),
   .I3(level4_in[3741]),
   .I4(level4_in[3742]),
   .I5(level4_in[3743])
);

LUT6 #(
   .INIT(64'h61f593b061f593b0)  
) LUT6_inst8400 (
   .O(to_level3[624]),
   .I0(level4_in[3744]),
   .I1(level4_in[3745]),
   .I2(level4_in[3746]),
   .I3(level4_in[3747]),
   .I4(level4_in[3748]),
   .I5(level4_in[3749])
);

LUT6 #(
   .INIT(64'h840fe034840fe034)  
) LUT6_inst8401 (
   .O(to_level3[625]),
   .I0(level4_in[3750]),
   .I1(level4_in[3751]),
   .I2(level4_in[3752]),
   .I3(level4_in[3753]),
   .I4(level4_in[3754]),
   .I5(level4_in[3755])
);

LUT6 #(
   .INIT(64'hd68b0d61d68b0d61)  
) LUT6_inst8402 (
   .O(to_level3[626]),
   .I0(level4_in[3756]),
   .I1(level4_in[3757]),
   .I2(level4_in[3758]),
   .I3(level4_in[3759]),
   .I4(level4_in[3760]),
   .I5(level4_in[3761])
);

LUT6 #(
   .INIT(64'h1eb9ea001eb9ea00)  
) LUT6_inst8403 (
   .O(to_level3[627]),
   .I0(level4_in[3762]),
   .I1(level4_in[3763]),
   .I2(level4_in[3764]),
   .I3(level4_in[3765]),
   .I4(level4_in[3766]),
   .I5(level4_in[3767])
);

LUT6 #(
   .INIT(64'hf5fbae01f5fbae01)  
) LUT6_inst8404 (
   .O(to_level3[628]),
   .I0(level4_in[3768]),
   .I1(level4_in[3769]),
   .I2(level4_in[3770]),
   .I3(level4_in[3771]),
   .I4(level4_in[3772]),
   .I5(level4_in[3773])
);

LUT6 #(
   .INIT(64'h31a7c8f431a7c8f4)  
) LUT6_inst8405 (
   .O(to_level3[629]),
   .I0(level4_in[3774]),
   .I1(level4_in[3775]),
   .I2(level4_in[3776]),
   .I3(level4_in[3777]),
   .I4(level4_in[3778]),
   .I5(level4_in[3779])
);

LUT6 #(
   .INIT(64'h19feb0bf19feb0bf)  
) LUT6_inst8406 (
   .O(to_level3[630]),
   .I0(level4_in[3780]),
   .I1(level4_in[3781]),
   .I2(level4_in[3782]),
   .I3(level4_in[3783]),
   .I4(level4_in[3784]),
   .I5(level4_in[3785])
);

LUT6 #(
   .INIT(64'h60e49d4b60e49d4b)  
) LUT6_inst8407 (
   .O(to_level3[631]),
   .I0(level4_in[3786]),
   .I1(level4_in[3787]),
   .I2(level4_in[3788]),
   .I3(level4_in[3789]),
   .I4(level4_in[3790]),
   .I5(level4_in[3791])
);

LUT6 #(
   .INIT(64'h63ea023763ea0237)  
) LUT6_inst8408 (
   .O(to_level3[632]),
   .I0(level4_in[3792]),
   .I1(level4_in[3793]),
   .I2(level4_in[3794]),
   .I3(level4_in[3795]),
   .I4(level4_in[3796]),
   .I5(level4_in[3797])
);

LUT6 #(
   .INIT(64'h148cfe21148cfe21)  
) LUT6_inst8409 (
   .O(to_level3[633]),
   .I0(level4_in[3798]),
   .I1(level4_in[3799]),
   .I2(level4_in[3800]),
   .I3(level4_in[3801]),
   .I4(level4_in[3802]),
   .I5(level4_in[3803])
);

LUT6 #(
   .INIT(64'h396c0d88396c0d88)  
) LUT6_inst8410 (
   .O(to_level3[634]),
   .I0(level4_in[3804]),
   .I1(level4_in[3805]),
   .I2(level4_in[3806]),
   .I3(level4_in[3807]),
   .I4(level4_in[3808]),
   .I5(level4_in[3809])
);

LUT6 #(
   .INIT(64'hc3c76a0cc3c76a0c)  
) LUT6_inst8411 (
   .O(to_level3[635]),
   .I0(level4_in[3810]),
   .I1(level4_in[3811]),
   .I2(level4_in[3812]),
   .I3(level4_in[3813]),
   .I4(level4_in[3814]),
   .I5(level4_in[3815])
);

LUT6 #(
   .INIT(64'h9ce244a29ce244a2)  
) LUT6_inst8412 (
   .O(to_level3[636]),
   .I0(level4_in[3816]),
   .I1(level4_in[3817]),
   .I2(level4_in[3818]),
   .I3(level4_in[3819]),
   .I4(level4_in[3820]),
   .I5(level4_in[3821])
);

LUT6 #(
   .INIT(64'hef023486ef023486)  
) LUT6_inst8413 (
   .O(to_level3[637]),
   .I0(level4_in[3822]),
   .I1(level4_in[3823]),
   .I2(level4_in[3824]),
   .I3(level4_in[3825]),
   .I4(level4_in[3826]),
   .I5(level4_in[3827])
);

LUT6 #(
   .INIT(64'h03a3093c03a3093c)  
) LUT6_inst8414 (
   .O(to_level3[638]),
   .I0(level4_in[3828]),
   .I1(level4_in[3829]),
   .I2(level4_in[3830]),
   .I3(level4_in[3831]),
   .I4(level4_in[3832]),
   .I5(level4_in[3833])
);

LUT6 #(
   .INIT(64'h6e0bedaa6e0bedaa)  
) LUT6_inst8415 (
   .O(to_level3[639]),
   .I0(level4_in[3834]),
   .I1(level4_in[3835]),
   .I2(level4_in[3836]),
   .I3(level4_in[3837]),
   .I4(level4_in[3838]),
   .I5(level4_in[3839])
);

LUT6 #(
   .INIT(64'h47acc9c247acc9c2)  
) LUT6_inst8416 (
   .O(to_level3[640]),
   .I0(level4_in[3840]),
   .I1(level4_in[3841]),
   .I2(level4_in[3842]),
   .I3(level4_in[3843]),
   .I4(level4_in[3844]),
   .I5(level4_in[3845])
);

LUT6 #(
   .INIT(64'h62e9fed762e9fed7)  
) LUT6_inst8417 (
   .O(to_level3[641]),
   .I0(level4_in[3846]),
   .I1(level4_in[3847]),
   .I2(level4_in[3848]),
   .I3(level4_in[3849]),
   .I4(level4_in[3850]),
   .I5(level4_in[3851])
);

LUT6 #(
   .INIT(64'h9cf9481e9cf9481e)  
) LUT6_inst8418 (
   .O(to_level3[642]),
   .I0(level4_in[3852]),
   .I1(level4_in[3853]),
   .I2(level4_in[3854]),
   .I3(level4_in[3855]),
   .I4(level4_in[3856]),
   .I5(level4_in[3857])
);

LUT6 #(
   .INIT(64'ha4864141a4864141)  
) LUT6_inst8419 (
   .O(to_level3[643]),
   .I0(level4_in[3858]),
   .I1(level4_in[3859]),
   .I2(level4_in[3860]),
   .I3(level4_in[3861]),
   .I4(level4_in[3862]),
   .I5(level4_in[3863])
);

LUT6 #(
   .INIT(64'h98ff86d098ff86d0)  
) LUT6_inst8420 (
   .O(to_level3[644]),
   .I0(level4_in[3864]),
   .I1(level4_in[3865]),
   .I2(level4_in[3866]),
   .I3(level4_in[3867]),
   .I4(level4_in[3868]),
   .I5(level4_in[3869])
);

LUT6 #(
   .INIT(64'h805c1eb7805c1eb7)  
) LUT6_inst8421 (
   .O(to_level3[645]),
   .I0(level4_in[3870]),
   .I1(level4_in[3871]),
   .I2(level4_in[3872]),
   .I3(level4_in[3873]),
   .I4(level4_in[3874]),
   .I5(level4_in[3875])
);

LUT6 #(
   .INIT(64'he2052f59e2052f59)  
) LUT6_inst8422 (
   .O(to_level3[646]),
   .I0(level4_in[3876]),
   .I1(level4_in[3877]),
   .I2(level4_in[3878]),
   .I3(level4_in[3879]),
   .I4(level4_in[3880]),
   .I5(level4_in[3881])
);

LUT6 #(
   .INIT(64'h1eba51f11eba51f1)  
) LUT6_inst8423 (
   .O(to_level3[647]),
   .I0(level4_in[3882]),
   .I1(level4_in[3883]),
   .I2(level4_in[3884]),
   .I3(level4_in[3885]),
   .I4(level4_in[3886]),
   .I5(level4_in[3887])
);

LUT6 #(
   .INIT(64'hc83e2106c83e2106)  
) LUT6_inst8424 (
   .O(to_level3[648]),
   .I0(level4_in[3888]),
   .I1(level4_in[3889]),
   .I2(level4_in[3890]),
   .I3(level4_in[3891]),
   .I4(level4_in[3892]),
   .I5(level4_in[3893])
);

LUT6 #(
   .INIT(64'h69e368a369e368a3)  
) LUT6_inst8425 (
   .O(to_level3[649]),
   .I0(level4_in[3894]),
   .I1(level4_in[3895]),
   .I2(level4_in[3896]),
   .I3(level4_in[3897]),
   .I4(level4_in[3898]),
   .I5(level4_in[3899])
);

LUT6 #(
   .INIT(64'h6cd786296cd78629)  
) LUT6_inst8426 (
   .O(to_level3[650]),
   .I0(level4_in[3900]),
   .I1(level4_in[3901]),
   .I2(level4_in[3902]),
   .I3(level4_in[3903]),
   .I4(level4_in[3904]),
   .I5(level4_in[3905])
);

LUT6 #(
   .INIT(64'h7f5699be7f5699be)  
) LUT6_inst8427 (
   .O(to_level3[651]),
   .I0(level4_in[3906]),
   .I1(level4_in[3907]),
   .I2(level4_in[3908]),
   .I3(level4_in[3909]),
   .I4(level4_in[3910]),
   .I5(level4_in[3911])
);

LUT6 #(
   .INIT(64'h1a2ae0741a2ae074)  
) LUT6_inst8428 (
   .O(to_level3[652]),
   .I0(level4_in[3912]),
   .I1(level4_in[3913]),
   .I2(level4_in[3914]),
   .I3(level4_in[3915]),
   .I4(level4_in[3916]),
   .I5(level4_in[3917])
);

LUT6 #(
   .INIT(64'h5495112854951128)  
) LUT6_inst8429 (
   .O(to_level3[653]),
   .I0(level4_in[3918]),
   .I1(level4_in[3919]),
   .I2(level4_in[3920]),
   .I3(level4_in[3921]),
   .I4(level4_in[3922]),
   .I5(level4_in[3923])
);

LUT6 #(
   .INIT(64'h58ee029258ee0292)  
) LUT6_inst8430 (
   .O(to_level3[654]),
   .I0(level4_in[3924]),
   .I1(level4_in[3925]),
   .I2(level4_in[3926]),
   .I3(level4_in[3927]),
   .I4(level4_in[3928]),
   .I5(level4_in[3929])
);

LUT6 #(
   .INIT(64'h8284377382843773)  
) LUT6_inst8431 (
   .O(to_level3[655]),
   .I0(level4_in[3930]),
   .I1(level4_in[3931]),
   .I2(level4_in[3932]),
   .I3(level4_in[3933]),
   .I4(level4_in[3934]),
   .I5(level4_in[3935])
);

LUT6 #(
   .INIT(64'h19efba0f19efba0f)  
) LUT6_inst8432 (
   .O(to_level3[656]),
   .I0(level4_in[3936]),
   .I1(level4_in[3937]),
   .I2(level4_in[3938]),
   .I3(level4_in[3939]),
   .I4(level4_in[3940]),
   .I5(level4_in[3941])
);

LUT6 #(
   .INIT(64'hcfb14d8bcfb14d8b)  
) LUT6_inst8433 (
   .O(to_level3[657]),
   .I0(level4_in[3942]),
   .I1(level4_in[3943]),
   .I2(level4_in[3944]),
   .I3(level4_in[3945]),
   .I4(level4_in[3946]),
   .I5(level4_in[3947])
);

LUT6 #(
   .INIT(64'h8d050a888d050a88)  
) LUT6_inst8434 (
   .O(to_level3[658]),
   .I0(level4_in[3948]),
   .I1(level4_in[3949]),
   .I2(level4_in[3950]),
   .I3(level4_in[3951]),
   .I4(level4_in[3952]),
   .I5(level4_in[3953])
);

LUT6 #(
   .INIT(64'h5a0df6ed5a0df6ed)  
) LUT6_inst8435 (
   .O(to_level3[659]),
   .I0(level4_in[3954]),
   .I1(level4_in[3955]),
   .I2(level4_in[3956]),
   .I3(level4_in[3957]),
   .I4(level4_in[3958]),
   .I5(level4_in[3959])
);

LUT6 #(
   .INIT(64'h792445b0792445b0)  
) LUT6_inst8436 (
   .O(to_level3[660]),
   .I0(level4_in[3960]),
   .I1(level4_in[3961]),
   .I2(level4_in[3962]),
   .I3(level4_in[3963]),
   .I4(level4_in[3964]),
   .I5(level4_in[3965])
);

LUT6 #(
   .INIT(64'h322672f4322672f4)  
) LUT6_inst8437 (
   .O(to_level3[661]),
   .I0(level4_in[3966]),
   .I1(level4_in[3967]),
   .I2(level4_in[3968]),
   .I3(level4_in[3969]),
   .I4(level4_in[3970]),
   .I5(level4_in[3971])
);

LUT6 #(
   .INIT(64'h8d8256d98d8256d9)  
) LUT6_inst8438 (
   .O(to_level3[662]),
   .I0(level4_in[3972]),
   .I1(level4_in[3973]),
   .I2(level4_in[3974]),
   .I3(level4_in[3975]),
   .I4(level4_in[3976]),
   .I5(level4_in[3977])
);

LUT6 #(
   .INIT(64'h14a465de14a465de)  
) LUT6_inst8439 (
   .O(to_level3[663]),
   .I0(level4_in[3978]),
   .I1(level4_in[3979]),
   .I2(level4_in[3980]),
   .I3(level4_in[3981]),
   .I4(level4_in[3982]),
   .I5(level4_in[3983])
);

LUT6 #(
   .INIT(64'h05c1ba5305c1ba53)  
) LUT6_inst8440 (
   .O(to_level3[664]),
   .I0(level4_in[3984]),
   .I1(level4_in[3985]),
   .I2(level4_in[3986]),
   .I3(level4_in[3987]),
   .I4(level4_in[3988]),
   .I5(level4_in[3989])
);

LUT6 #(
   .INIT(64'h8f1f06be8f1f06be)  
) LUT6_inst8441 (
   .O(to_level3[665]),
   .I0(level4_in[3990]),
   .I1(level4_in[3991]),
   .I2(level4_in[3992]),
   .I3(level4_in[3993]),
   .I4(level4_in[3994]),
   .I5(level4_in[3995])
);

LUT6 #(
   .INIT(64'h5e09ae535e09ae53)  
) LUT6_inst8442 (
   .O(to_level3[666]),
   .I0(level4_in[3996]),
   .I1(level4_in[3997]),
   .I2(level4_in[3998]),
   .I3(level4_in[3999]),
   .I4(level4_in[4000]),
   .I5(level4_in[4001])
);

LUT6 #(
   .INIT(64'h14fb82dd14fb82dd)  
) LUT6_inst8443 (
   .O(to_level3[667]),
   .I0(level4_in[4002]),
   .I1(level4_in[4003]),
   .I2(level4_in[4004]),
   .I3(level4_in[4005]),
   .I4(level4_in[4006]),
   .I5(level4_in[4007])
);

LUT6 #(
   .INIT(64'hd325128bd325128b)  
) LUT6_inst8444 (
   .O(to_level3[668]),
   .I0(level4_in[4008]),
   .I1(level4_in[4009]),
   .I2(level4_in[4010]),
   .I3(level4_in[4011]),
   .I4(level4_in[4012]),
   .I5(level4_in[4013])
);

LUT6 #(
   .INIT(64'h7c12eecb7c12eecb)  
) LUT6_inst8445 (
   .O(to_level3[669]),
   .I0(level4_in[4014]),
   .I1(level4_in[4015]),
   .I2(level4_in[4016]),
   .I3(level4_in[4017]),
   .I4(level4_in[4018]),
   .I5(level4_in[4019])
);

LUT6 #(
   .INIT(64'h03aa199a03aa199a)  
) LUT6_inst8446 (
   .O(to_level3[670]),
   .I0(level4_in[4020]),
   .I1(level4_in[4021]),
   .I2(level4_in[4022]),
   .I3(level4_in[4023]),
   .I4(level4_in[4024]),
   .I5(level4_in[4025])
);

LUT6 #(
   .INIT(64'hc6ae3b75c6ae3b75)  
) LUT6_inst8447 (
   .O(to_level3[671]),
   .I0(level4_in[4026]),
   .I1(level4_in[4027]),
   .I2(level4_in[4028]),
   .I3(level4_in[4029]),
   .I4(level4_in[4030]),
   .I5(level4_in[4031])
);

LUT6 #(
   .INIT(64'hef11d3feef11d3fe)  
) LUT6_inst8448 (
   .O(to_level3[672]),
   .I0(level4_in[4032]),
   .I1(level4_in[4033]),
   .I2(level4_in[4034]),
   .I3(level4_in[4035]),
   .I4(level4_in[4036]),
   .I5(level4_in[4037])
);

LUT6 #(
   .INIT(64'h3d33b3313d33b331)  
) LUT6_inst8449 (
   .O(to_level3[673]),
   .I0(level4_in[4038]),
   .I1(level4_in[4039]),
   .I2(level4_in[4040]),
   .I3(level4_in[4041]),
   .I4(level4_in[4042]),
   .I5(level4_in[4043])
);

LUT6 #(
   .INIT(64'hd4e29247d4e29247)  
) LUT6_inst8450 (
   .O(to_level3[674]),
   .I0(level4_in[4044]),
   .I1(level4_in[4045]),
   .I2(level4_in[4046]),
   .I3(level4_in[4047]),
   .I4(level4_in[4048]),
   .I5(level4_in[4049])
);

LUT6 #(
   .INIT(64'hc2f8e006c2f8e006)  
) LUT6_inst8451 (
   .O(to_level3[675]),
   .I0(level4_in[4050]),
   .I1(level4_in[4051]),
   .I2(level4_in[4052]),
   .I3(level4_in[4053]),
   .I4(level4_in[4054]),
   .I5(level4_in[4055])
);

LUT6 #(
   .INIT(64'ha0ce3828a0ce3828)  
) LUT6_inst8452 (
   .O(to_level3[676]),
   .I0(level4_in[4056]),
   .I1(level4_in[4057]),
   .I2(level4_in[4058]),
   .I3(level4_in[4059]),
   .I4(level4_in[4060]),
   .I5(level4_in[4061])
);

LUT6 #(
   .INIT(64'hfad2bac9fad2bac9)  
) LUT6_inst8453 (
   .O(to_level3[677]),
   .I0(level4_in[4062]),
   .I1(level4_in[4063]),
   .I2(level4_in[4064]),
   .I3(level4_in[4065]),
   .I4(level4_in[4066]),
   .I5(level4_in[4067])
);

LUT6 #(
   .INIT(64'h03a9c1c703a9c1c7)  
) LUT6_inst8454 (
   .O(to_level3[678]),
   .I0(level4_in[4068]),
   .I1(level4_in[4069]),
   .I2(level4_in[4070]),
   .I3(level4_in[4071]),
   .I4(level4_in[4072]),
   .I5(level4_in[4073])
);

LUT6 #(
   .INIT(64'hf48e90f4f48e90f4)  
) LUT6_inst8455 (
   .O(to_level3[679]),
   .I0(level4_in[4074]),
   .I1(level4_in[4075]),
   .I2(level4_in[4076]),
   .I3(level4_in[4077]),
   .I4(level4_in[4078]),
   .I5(level4_in[4079])
);

LUT6 #(
   .INIT(64'h73d42b8673d42b86)  
) LUT6_inst8456 (
   .O(to_level3[680]),
   .I0(level4_in[4080]),
   .I1(level4_in[4081]),
   .I2(level4_in[4082]),
   .I3(level4_in[4083]),
   .I4(level4_in[4084]),
   .I5(level4_in[4085])
);

LUT6 #(
   .INIT(64'h05cacd4105cacd41)  
) LUT6_inst8457 (
   .O(to_level3[681]),
   .I0(level4_in[4086]),
   .I1(level4_in[4087]),
   .I2(level4_in[4088]),
   .I3(level4_in[4089]),
   .I4(level4_in[4090]),
   .I5(level4_in[4091])
);

LUT6 #(
   .INIT(64'h4b36c18c4b36c18c)  
) LUT6_inst8458 (
   .O(to_level3[682]),
   .I0(level4_in[4092]),
   .I1(level4_in[4093]),
   .I2(level4_in[4094]),
   .I3(level4_in[4095]),
   .I4(level4_in[4096]),
   .I5(level4_in[4097])
);

LUT6 #(
   .INIT(64'h43622a7743622a77)  
) LUT6_inst8459 (
   .O(to_level3[683]),
   .I0(level4_in[4098]),
   .I1(level4_in[4099]),
   .I2(level4_in[4100]),
   .I3(level4_in[4101]),
   .I4(level4_in[4102]),
   .I5(level4_in[4103])
);

LUT6 #(
   .INIT(64'hff46267eff46267e)  
) LUT6_inst8460 (
   .O(to_level3[684]),
   .I0(level4_in[4104]),
   .I1(level4_in[4105]),
   .I2(level4_in[4106]),
   .I3(level4_in[4107]),
   .I4(level4_in[4108]),
   .I5(level4_in[4109])
);

LUT6 #(
   .INIT(64'hfa56837efa56837e)  
) LUT6_inst8461 (
   .O(to_level3[685]),
   .I0(level4_in[4110]),
   .I1(level4_in[4111]),
   .I2(level4_in[4112]),
   .I3(level4_in[4113]),
   .I4(level4_in[4114]),
   .I5(level4_in[4115])
);

LUT6 #(
   .INIT(64'h3e498cdb3e498cdb)  
) LUT6_inst8462 (
   .O(to_level3[686]),
   .I0(level4_in[4116]),
   .I1(level4_in[4117]),
   .I2(level4_in[4118]),
   .I3(level4_in[4119]),
   .I4(level4_in[4120]),
   .I5(level4_in[4121])
);

LUT6 #(
   .INIT(64'hbef5e0bebef5e0be)  
) LUT6_inst8463 (
   .O(to_level3[687]),
   .I0(level4_in[4122]),
   .I1(level4_in[4123]),
   .I2(level4_in[4124]),
   .I3(level4_in[4125]),
   .I4(level4_in[4126]),
   .I5(level4_in[4127])
);

LUT6 #(
   .INIT(64'he4766217e4766217)  
) LUT6_inst8464 (
   .O(to_level3[688]),
   .I0(level4_in[4128]),
   .I1(level4_in[4129]),
   .I2(level4_in[4130]),
   .I3(level4_in[4131]),
   .I4(level4_in[4132]),
   .I5(level4_in[4133])
);

LUT6 #(
   .INIT(64'h7c1a35e67c1a35e6)  
) LUT6_inst8465 (
   .O(to_level3[689]),
   .I0(level4_in[4134]),
   .I1(level4_in[4135]),
   .I2(level4_in[4136]),
   .I3(level4_in[4137]),
   .I4(level4_in[4138]),
   .I5(level4_in[4139])
);

LUT6 #(
   .INIT(64'ha8f37cd0a8f37cd0)  
) LUT6_inst8466 (
   .O(to_level3[690]),
   .I0(level4_in[4140]),
   .I1(level4_in[4141]),
   .I2(level4_in[4142]),
   .I3(level4_in[4143]),
   .I4(level4_in[4144]),
   .I5(level4_in[4145])
);

LUT6 #(
   .INIT(64'had22e3a9ad22e3a9)  
) LUT6_inst8467 (
   .O(to_level3[691]),
   .I0(level4_in[4146]),
   .I1(level4_in[4147]),
   .I2(level4_in[4148]),
   .I3(level4_in[4149]),
   .I4(level4_in[4150]),
   .I5(level4_in[4151])
);

LUT6 #(
   .INIT(64'h483fcdaf483fcdaf)  
) LUT6_inst8468 (
   .O(to_level3[692]),
   .I0(level4_in[4152]),
   .I1(level4_in[4153]),
   .I2(level4_in[4154]),
   .I3(level4_in[4155]),
   .I4(level4_in[4156]),
   .I5(level4_in[4157])
);

LUT6 #(
   .INIT(64'h6729bc166729bc16)  
) LUT6_inst8469 (
   .O(to_level3[693]),
   .I0(level4_in[4158]),
   .I1(level4_in[4159]),
   .I2(level4_in[4160]),
   .I3(level4_in[4161]),
   .I4(level4_in[4162]),
   .I5(level4_in[4163])
);

LUT6 #(
   .INIT(64'h9dcddeaa9dcddeaa)  
) LUT6_inst8470 (
   .O(to_level3[694]),
   .I0(level4_in[4164]),
   .I1(level4_in[4165]),
   .I2(level4_in[4166]),
   .I3(level4_in[4167]),
   .I4(level4_in[4168]),
   .I5(level4_in[4169])
);

LUT6 #(
   .INIT(64'h7f11e5507f11e550)  
) LUT6_inst8471 (
   .O(to_level3[695]),
   .I0(level4_in[4170]),
   .I1(level4_in[4171]),
   .I2(level4_in[4172]),
   .I3(level4_in[4173]),
   .I4(level4_in[4174]),
   .I5(level4_in[4175])
);

LUT6 #(
   .INIT(64'h1cccc0361cccc036)  
) LUT6_inst8472 (
   .O(to_level3[696]),
   .I0(level4_in[4176]),
   .I1(level4_in[4177]),
   .I2(level4_in[4178]),
   .I3(level4_in[4179]),
   .I4(level4_in[4180]),
   .I5(level4_in[4181])
);

LUT6 #(
   .INIT(64'haed0837daed0837d)  
) LUT6_inst8473 (
   .O(to_level3[697]),
   .I0(level4_in[4182]),
   .I1(level4_in[4183]),
   .I2(level4_in[4184]),
   .I3(level4_in[4185]),
   .I4(level4_in[4186]),
   .I5(level4_in[4187])
);

LUT6 #(
   .INIT(64'h4aa06e5c4aa06e5c)  
) LUT6_inst8474 (
   .O(to_level3[698]),
   .I0(level4_in[4188]),
   .I1(level4_in[4189]),
   .I2(level4_in[4190]),
   .I3(level4_in[4191]),
   .I4(level4_in[4192]),
   .I5(level4_in[4193])
);

LUT6 #(
   .INIT(64'hbe77469cbe77469c)  
) LUT6_inst8475 (
   .O(to_level3[699]),
   .I0(level4_in[4194]),
   .I1(level4_in[4195]),
   .I2(level4_in[4196]),
   .I3(level4_in[4197]),
   .I4(level4_in[4198]),
   .I5(level4_in[4199])
);

LUT6 #(
   .INIT(64'ha9c189a3a9c189a3)  
) LUT6_inst8476 (
   .O(to_level3[700]),
   .I0(level4_in[4200]),
   .I1(level4_in[4201]),
   .I2(level4_in[4202]),
   .I3(level4_in[4203]),
   .I4(level4_in[4204]),
   .I5(level4_in[4205])
);

LUT6 #(
   .INIT(64'h7f2ce3417f2ce341)  
) LUT6_inst8477 (
   .O(to_level3[701]),
   .I0(level4_in[4206]),
   .I1(level4_in[4207]),
   .I2(level4_in[4208]),
   .I3(level4_in[4209]),
   .I4(level4_in[4210]),
   .I5(level4_in[4211])
);

LUT6 #(
   .INIT(64'hf2ffb7bef2ffb7be)  
) LUT6_inst8478 (
   .O(to_level3[702]),
   .I0(level4_in[4212]),
   .I1(level4_in[4213]),
   .I2(level4_in[4214]),
   .I3(level4_in[4215]),
   .I4(level4_in[4216]),
   .I5(level4_in[4217])
);

LUT6 #(
   .INIT(64'h19651b3d19651b3d)  
) LUT6_inst8479 (
   .O(to_level3[703]),
   .I0(level4_in[4218]),
   .I1(level4_in[4219]),
   .I2(level4_in[4220]),
   .I3(level4_in[4221]),
   .I4(level4_in[4222]),
   .I5(level4_in[4223])
);

LUT6 #(
   .INIT(64'h4f31e5e04f31e5e0)  
) LUT6_inst8480 (
   .O(to_level3[704]),
   .I0(level4_in[4224]),
   .I1(level4_in[4225]),
   .I2(level4_in[4226]),
   .I3(level4_in[4227]),
   .I4(level4_in[4228]),
   .I5(level4_in[4229])
);

LUT6 #(
   .INIT(64'h2f42b8bb2f42b8bb)  
) LUT6_inst8481 (
   .O(to_level3[705]),
   .I0(level4_in[4230]),
   .I1(level4_in[4231]),
   .I2(level4_in[4232]),
   .I3(level4_in[4233]),
   .I4(level4_in[4234]),
   .I5(level4_in[4235])
);

LUT6 #(
   .INIT(64'h146bf6bd146bf6bd)  
) LUT6_inst8482 (
   .O(to_level3[706]),
   .I0(level4_in[4236]),
   .I1(level4_in[4237]),
   .I2(level4_in[4238]),
   .I3(level4_in[4239]),
   .I4(level4_in[4240]),
   .I5(level4_in[4241])
);

LUT6 #(
   .INIT(64'h9c48e5c79c48e5c7)  
) LUT6_inst8483 (
   .O(to_level3[707]),
   .I0(level4_in[4242]),
   .I1(level4_in[4243]),
   .I2(level4_in[4244]),
   .I3(level4_in[4245]),
   .I4(level4_in[4246]),
   .I5(level4_in[4247])
);

LUT6 #(
   .INIT(64'h899b5fcc899b5fcc)  
) LUT6_inst8484 (
   .O(to_level3[708]),
   .I0(level4_in[4248]),
   .I1(level4_in[4249]),
   .I2(level4_in[4250]),
   .I3(level4_in[4251]),
   .I4(level4_in[4252]),
   .I5(level4_in[4253])
);

LUT6 #(
   .INIT(64'h1cd86c0a1cd86c0a)  
) LUT6_inst8485 (
   .O(to_level3[709]),
   .I0(level4_in[4254]),
   .I1(level4_in[4255]),
   .I2(level4_in[4256]),
   .I3(level4_in[4257]),
   .I4(level4_in[4258]),
   .I5(level4_in[4259])
);

LUT6 #(
   .INIT(64'h5612da0a5612da0a)  
) LUT6_inst8486 (
   .O(to_level3[710]),
   .I0(level4_in[4260]),
   .I1(level4_in[4261]),
   .I2(level4_in[4262]),
   .I3(level4_in[4263]),
   .I4(level4_in[4264]),
   .I5(level4_in[4265])
);

LUT6 #(
   .INIT(64'h270b3af2270b3af2)  
) LUT6_inst8487 (
   .O(to_level3[711]),
   .I0(level4_in[4266]),
   .I1(level4_in[4267]),
   .I2(level4_in[4268]),
   .I3(level4_in[4269]),
   .I4(level4_in[4270]),
   .I5(level4_in[4271])
);

LUT6 #(
   .INIT(64'h29bbf7da29bbf7da)  
) LUT6_inst8488 (
   .O(to_level3[712]),
   .I0(level4_in[4272]),
   .I1(level4_in[4273]),
   .I2(level4_in[4274]),
   .I3(level4_in[4275]),
   .I4(level4_in[4276]),
   .I5(level4_in[4277])
);

LUT6 #(
   .INIT(64'h0b0d2c2f0b0d2c2f)  
) LUT6_inst8489 (
   .O(to_level3[713]),
   .I0(level4_in[4278]),
   .I1(level4_in[4279]),
   .I2(level4_in[4280]),
   .I3(level4_in[4281]),
   .I4(level4_in[4282]),
   .I5(level4_in[4283])
);

LUT6 #(
   .INIT(64'h75abd13a75abd13a)  
) LUT6_inst8490 (
   .O(to_level3[714]),
   .I0(level4_in[4284]),
   .I1(level4_in[4285]),
   .I2(level4_in[4286]),
   .I3(level4_in[4287]),
   .I4(level4_in[4288]),
   .I5(level4_in[4289])
);

LUT6 #(
   .INIT(64'h05e4ec3b05e4ec3b)  
) LUT6_inst8491 (
   .O(to_level3[715]),
   .I0(level4_in[4290]),
   .I1(level4_in[4291]),
   .I2(level4_in[4292]),
   .I3(level4_in[4293]),
   .I4(level4_in[4294]),
   .I5(level4_in[4295])
);

LUT6 #(
   .INIT(64'hf8d89ab3f8d89ab3)  
) LUT6_inst8492 (
   .O(to_level3[716]),
   .I0(level4_in[4296]),
   .I1(level4_in[4297]),
   .I2(level4_in[4298]),
   .I3(level4_in[4299]),
   .I4(level4_in[4300]),
   .I5(level4_in[4301])
);

LUT6 #(
   .INIT(64'h9c3ee4129c3ee412)  
) LUT6_inst8493 (
   .O(to_level3[717]),
   .I0(level4_in[4302]),
   .I1(level4_in[4303]),
   .I2(level4_in[4304]),
   .I3(level4_in[4305]),
   .I4(level4_in[4306]),
   .I5(level4_in[4307])
);

LUT6 #(
   .INIT(64'h790f27e8790f27e8)  
) LUT6_inst8494 (
   .O(to_level3[718]),
   .I0(level4_in[4308]),
   .I1(level4_in[4309]),
   .I2(level4_in[4310]),
   .I3(level4_in[4311]),
   .I4(level4_in[4312]),
   .I5(level4_in[4313])
);

LUT6 #(
   .INIT(64'h8a97a0f28a97a0f2)  
) LUT6_inst8495 (
   .O(to_level3[719]),
   .I0(level4_in[4314]),
   .I1(level4_in[4315]),
   .I2(level4_in[4316]),
   .I3(level4_in[4317]),
   .I4(level4_in[4318]),
   .I5(level4_in[4319])
);

LUT6 #(
   .INIT(64'h0ba5a7f10ba5a7f1)  
) LUT6_inst8496 (
   .O(to_level3[720]),
   .I0(level4_in[4320]),
   .I1(level4_in[4321]),
   .I2(level4_in[4322]),
   .I3(level4_in[4323]),
   .I4(level4_in[4324]),
   .I5(level4_in[4325])
);

LUT6 #(
   .INIT(64'hd656f19fd656f19f)  
) LUT6_inst8497 (
   .O(to_level3[721]),
   .I0(level4_in[4326]),
   .I1(level4_in[4327]),
   .I2(level4_in[4328]),
   .I3(level4_in[4329]),
   .I4(level4_in[4330]),
   .I5(level4_in[4331])
);

LUT6 #(
   .INIT(64'h517e7e73517e7e73)  
) LUT6_inst8498 (
   .O(to_level3[722]),
   .I0(level4_in[4332]),
   .I1(level4_in[4333]),
   .I2(level4_in[4334]),
   .I3(level4_in[4335]),
   .I4(level4_in[4336]),
   .I5(level4_in[4337])
);

LUT6 #(
   .INIT(64'h3033dc7e3033dc7e)  
) LUT6_inst8499 (
   .O(to_level3[723]),
   .I0(level4_in[4338]),
   .I1(level4_in[4339]),
   .I2(level4_in[4340]),
   .I3(level4_in[4341]),
   .I4(level4_in[4342]),
   .I5(level4_in[4343])
);

LUT6 #(
   .INIT(64'h8d364df78d364df7)  
) LUT6_inst8500 (
   .O(to_level3[724]),
   .I0(level4_in[4344]),
   .I1(level4_in[4345]),
   .I2(level4_in[4346]),
   .I3(level4_in[4347]),
   .I4(level4_in[4348]),
   .I5(level4_in[4349])
);

LUT6 #(
   .INIT(64'hc9b9a084c9b9a084)  
) LUT6_inst8501 (
   .O(to_level3[725]),
   .I0(level4_in[4350]),
   .I1(level4_in[4351]),
   .I2(level4_in[4352]),
   .I3(level4_in[4353]),
   .I4(level4_in[4354]),
   .I5(level4_in[4355])
);

LUT6 #(
   .INIT(64'h65e9335d65e9335d)  
) LUT6_inst8502 (
   .O(to_level3[726]),
   .I0(level4_in[4356]),
   .I1(level4_in[4357]),
   .I2(level4_in[4358]),
   .I3(level4_in[4359]),
   .I4(level4_in[4360]),
   .I5(level4_in[4361])
);

LUT6 #(
   .INIT(64'hbc3554eabc3554ea)  
) LUT6_inst8503 (
   .O(to_level3[727]),
   .I0(level4_in[4362]),
   .I1(level4_in[4363]),
   .I2(level4_in[4364]),
   .I3(level4_in[4365]),
   .I4(level4_in[4366]),
   .I5(level4_in[4367])
);

LUT6 #(
   .INIT(64'hb2f52deab2f52dea)  
) LUT6_inst8504 (
   .O(to_level3[728]),
   .I0(level4_in[4368]),
   .I1(level4_in[4369]),
   .I2(level4_in[4370]),
   .I3(level4_in[4371]),
   .I4(level4_in[4372]),
   .I5(level4_in[4373])
);

LUT6 #(
   .INIT(64'hbd0a9f78bd0a9f78)  
) LUT6_inst8505 (
   .O(to_level3[729]),
   .I0(level4_in[4374]),
   .I1(level4_in[4375]),
   .I2(level4_in[4376]),
   .I3(level4_in[4377]),
   .I4(level4_in[4378]),
   .I5(level4_in[4379])
);

LUT6 #(
   .INIT(64'h157b87be157b87be)  
) LUT6_inst8506 (
   .O(to_level3[730]),
   .I0(level4_in[4380]),
   .I1(level4_in[4381]),
   .I2(level4_in[4382]),
   .I3(level4_in[4383]),
   .I4(level4_in[4384]),
   .I5(level4_in[4385])
);

LUT6 #(
   .INIT(64'hdb85d063db85d063)  
) LUT6_inst8507 (
   .O(to_level3[731]),
   .I0(level4_in[4386]),
   .I1(level4_in[4387]),
   .I2(level4_in[4388]),
   .I3(level4_in[4389]),
   .I4(level4_in[4390]),
   .I5(level4_in[4391])
);

LUT6 #(
   .INIT(64'h27dec52427dec524)  
) LUT6_inst8508 (
   .O(to_level3[732]),
   .I0(level4_in[4392]),
   .I1(level4_in[4393]),
   .I2(level4_in[4394]),
   .I3(level4_in[4395]),
   .I4(level4_in[4396]),
   .I5(level4_in[4397])
);

LUT6 #(
   .INIT(64'h02595c0202595c02)  
) LUT6_inst8509 (
   .O(to_level3[733]),
   .I0(level4_in[4398]),
   .I1(level4_in[4399]),
   .I2(level4_in[4400]),
   .I3(level4_in[4401]),
   .I4(level4_in[4402]),
   .I5(level4_in[4403])
);

LUT6 #(
   .INIT(64'hdbac2bc2dbac2bc2)  
) LUT6_inst8510 (
   .O(to_level3[734]),
   .I0(level4_in[4404]),
   .I1(level4_in[4405]),
   .I2(level4_in[4406]),
   .I3(level4_in[4407]),
   .I4(level4_in[4408]),
   .I5(level4_in[4409])
);

LUT6 #(
   .INIT(64'h9168950c9168950c)  
) LUT6_inst8511 (
   .O(to_level3[735]),
   .I0(level4_in[4410]),
   .I1(level4_in[4411]),
   .I2(level4_in[4412]),
   .I3(level4_in[4413]),
   .I4(level4_in[4414]),
   .I5(level4_in[4415])
);

LUT6 #(
   .INIT(64'h611627c2611627c2)  
) LUT6_inst8512 (
   .O(to_level3[736]),
   .I0(level4_in[4416]),
   .I1(level4_in[4417]),
   .I2(level4_in[4418]),
   .I3(level4_in[4419]),
   .I4(level4_in[4420]),
   .I5(level4_in[4421])
);

LUT6 #(
   .INIT(64'h3330069033300690)  
) LUT6_inst8513 (
   .O(to_level3[737]),
   .I0(level4_in[4422]),
   .I1(level4_in[4423]),
   .I2(level4_in[4424]),
   .I3(level4_in[4425]),
   .I4(level4_in[4426]),
   .I5(level4_in[4427])
);

LUT6 #(
   .INIT(64'h878f6f9a878f6f9a)  
) LUT6_inst8514 (
   .O(to_level3[738]),
   .I0(level4_in[4428]),
   .I1(level4_in[4429]),
   .I2(level4_in[4430]),
   .I3(level4_in[4431]),
   .I4(level4_in[4432]),
   .I5(level4_in[4433])
);

LUT6 #(
   .INIT(64'h2ca08baf2ca08baf)  
) LUT6_inst8515 (
   .O(to_level3[739]),
   .I0(level4_in[4434]),
   .I1(level4_in[4435]),
   .I2(level4_in[4436]),
   .I3(level4_in[4437]),
   .I4(level4_in[4438]),
   .I5(level4_in[4439])
);

LUT6 #(
   .INIT(64'h6d6105b86d6105b8)  
) LUT6_inst8516 (
   .O(to_level3[740]),
   .I0(level4_in[4440]),
   .I1(level4_in[4441]),
   .I2(level4_in[4442]),
   .I3(level4_in[4443]),
   .I4(level4_in[4444]),
   .I5(level4_in[4445])
);

LUT6 #(
   .INIT(64'h10885da510885da5)  
) LUT6_inst8517 (
   .O(to_level3[741]),
   .I0(level4_in[4446]),
   .I1(level4_in[4447]),
   .I2(level4_in[4448]),
   .I3(level4_in[4449]),
   .I4(level4_in[4450]),
   .I5(level4_in[4451])
);

LUT6 #(
   .INIT(64'hf478652bf478652b)  
) LUT6_inst8518 (
   .O(to_level3[742]),
   .I0(level4_in[4452]),
   .I1(level4_in[4453]),
   .I2(level4_in[4454]),
   .I3(level4_in[4455]),
   .I4(level4_in[4456]),
   .I5(level4_in[4457])
);

LUT6 #(
   .INIT(64'hb15c3916b15c3916)  
) LUT6_inst8519 (
   .O(to_level3[743]),
   .I0(level4_in[4458]),
   .I1(level4_in[4459]),
   .I2(level4_in[4460]),
   .I3(level4_in[4461]),
   .I4(level4_in[4462]),
   .I5(level4_in[4463])
);

LUT6 #(
   .INIT(64'hf3ddbf0df3ddbf0d)  
) LUT6_inst8520 (
   .O(to_level3[744]),
   .I0(level4_in[4464]),
   .I1(level4_in[4465]),
   .I2(level4_in[4466]),
   .I3(level4_in[4467]),
   .I4(level4_in[4468]),
   .I5(level4_in[4469])
);

LUT6 #(
   .INIT(64'h75a4b06675a4b066)  
) LUT6_inst8521 (
   .O(to_level3[745]),
   .I0(level4_in[4470]),
   .I1(level4_in[4471]),
   .I2(level4_in[4472]),
   .I3(level4_in[4473]),
   .I4(level4_in[4474]),
   .I5(level4_in[4475])
);

LUT6 #(
   .INIT(64'h2442de4e2442de4e)  
) LUT6_inst8522 (
   .O(to_level3[746]),
   .I0(level4_in[4476]),
   .I1(level4_in[4477]),
   .I2(level4_in[4478]),
   .I3(level4_in[4479]),
   .I4(level4_in[4480]),
   .I5(level4_in[4481])
);

LUT6 #(
   .INIT(64'hc005f813c005f813)  
) LUT6_inst8523 (
   .O(to_level3[747]),
   .I0(level4_in[4482]),
   .I1(level4_in[4483]),
   .I2(level4_in[4484]),
   .I3(level4_in[4485]),
   .I4(level4_in[4486]),
   .I5(level4_in[4487])
);

LUT6 #(
   .INIT(64'h4f07687d4f07687d)  
) LUT6_inst8524 (
   .O(to_level3[748]),
   .I0(level4_in[4488]),
   .I1(level4_in[4489]),
   .I2(level4_in[4490]),
   .I3(level4_in[4491]),
   .I4(level4_in[4492]),
   .I5(level4_in[4493])
);

LUT6 #(
   .INIT(64'h53473f0f53473f0f)  
) LUT6_inst8525 (
   .O(to_level3[749]),
   .I0(level4_in[4494]),
   .I1(level4_in[4495]),
   .I2(level4_in[4496]),
   .I3(level4_in[4497]),
   .I4(level4_in[4498]),
   .I5(level4_in[4499])
);

LUT6 #(
   .INIT(64'h42291ee242291ee2)  
) LUT6_inst8526 (
   .O(to_level3[750]),
   .I0(level4_in[4500]),
   .I1(level4_in[4501]),
   .I2(level4_in[4502]),
   .I3(level4_in[4503]),
   .I4(level4_in[4504]),
   .I5(level4_in[4505])
);

LUT6 #(
   .INIT(64'hff93a05aff93a05a)  
) LUT6_inst8527 (
   .O(to_level3[751]),
   .I0(level4_in[4506]),
   .I1(level4_in[4507]),
   .I2(level4_in[4508]),
   .I3(level4_in[4509]),
   .I4(level4_in[4510]),
   .I5(level4_in[4511])
);

LUT6 #(
   .INIT(64'h9ab7a2c99ab7a2c9)  
) LUT6_inst8528 (
   .O(to_level3[752]),
   .I0(level4_in[4512]),
   .I1(level4_in[4513]),
   .I2(level4_in[4514]),
   .I3(level4_in[4515]),
   .I4(level4_in[4516]),
   .I5(level4_in[4517])
);

LUT6 #(
   .INIT(64'hf68dacbff68dacbf)  
) LUT6_inst8529 (
   .O(to_level3[753]),
   .I0(level4_in[4518]),
   .I1(level4_in[4519]),
   .I2(level4_in[4520]),
   .I3(level4_in[4521]),
   .I4(level4_in[4522]),
   .I5(level4_in[4523])
);

LUT6 #(
   .INIT(64'hc1b22889c1b22889)  
) LUT6_inst8530 (
   .O(to_level3[754]),
   .I0(level4_in[4524]),
   .I1(level4_in[4525]),
   .I2(level4_in[4526]),
   .I3(level4_in[4527]),
   .I4(level4_in[4528]),
   .I5(level4_in[4529])
);

LUT6 #(
   .INIT(64'h0f6ad9570f6ad957)  
) LUT6_inst8531 (
   .O(to_level3[755]),
   .I0(level4_in[4530]),
   .I1(level4_in[4531]),
   .I2(level4_in[4532]),
   .I3(level4_in[4533]),
   .I4(level4_in[4534]),
   .I5(level4_in[4535])
);

LUT6 #(
   .INIT(64'h4351e2a44351e2a4)  
) LUT6_inst8532 (
   .O(to_level3[756]),
   .I0(level4_in[4536]),
   .I1(level4_in[4537]),
   .I2(level4_in[4538]),
   .I3(level4_in[4539]),
   .I4(level4_in[4540]),
   .I5(level4_in[4541])
);

LUT6 #(
   .INIT(64'h9200585a9200585a)  
) LUT6_inst8533 (
   .O(to_level3[757]),
   .I0(level4_in[4542]),
   .I1(level4_in[4543]),
   .I2(level4_in[4544]),
   .I3(level4_in[4545]),
   .I4(level4_in[4546]),
   .I5(level4_in[4547])
);

LUT6 #(
   .INIT(64'h1d00bdfb1d00bdfb)  
) LUT6_inst8534 (
   .O(to_level3[758]),
   .I0(level4_in[4548]),
   .I1(level4_in[4549]),
   .I2(level4_in[4550]),
   .I3(level4_in[4551]),
   .I4(level4_in[4552]),
   .I5(level4_in[4553])
);

LUT6 #(
   .INIT(64'hd63abe96d63abe96)  
) LUT6_inst8535 (
   .O(to_level3[759]),
   .I0(level4_in[4554]),
   .I1(level4_in[4555]),
   .I2(level4_in[4556]),
   .I3(level4_in[4557]),
   .I4(level4_in[4558]),
   .I5(level4_in[4559])
);

LUT6 #(
   .INIT(64'h02971aaa02971aaa)  
) LUT6_inst8536 (
   .O(to_level3[760]),
   .I0(level4_in[4560]),
   .I1(level4_in[4561]),
   .I2(level4_in[4562]),
   .I3(level4_in[4563]),
   .I4(level4_in[4564]),
   .I5(level4_in[4565])
);

LUT6 #(
   .INIT(64'hd4a654e9d4a654e9)  
) LUT6_inst8537 (
   .O(to_level3[761]),
   .I0(level4_in[4566]),
   .I1(level4_in[4567]),
   .I2(level4_in[4568]),
   .I3(level4_in[4569]),
   .I4(level4_in[4570]),
   .I5(level4_in[4571])
);

LUT6 #(
   .INIT(64'hda742482da742482)  
) LUT6_inst8538 (
   .O(to_level3[762]),
   .I0(level4_in[4572]),
   .I1(level4_in[4573]),
   .I2(level4_in[4574]),
   .I3(level4_in[4575]),
   .I4(level4_in[4576]),
   .I5(level4_in[4577])
);

LUT6 #(
   .INIT(64'h862f396b862f396b)  
) LUT6_inst8539 (
   .O(to_level3[763]),
   .I0(level4_in[4578]),
   .I1(level4_in[4579]),
   .I2(level4_in[4580]),
   .I3(level4_in[4581]),
   .I4(level4_in[4582]),
   .I5(level4_in[4583])
);

LUT6 #(
   .INIT(64'h7997ef267997ef26)  
) LUT6_inst8540 (
   .O(to_level3[764]),
   .I0(level4_in[4584]),
   .I1(level4_in[4585]),
   .I2(level4_in[4586]),
   .I3(level4_in[4587]),
   .I4(level4_in[4588]),
   .I5(level4_in[4589])
);

LUT6 #(
   .INIT(64'h3fc363383fc36338)  
) LUT6_inst8541 (
   .O(to_level3[765]),
   .I0(level4_in[4590]),
   .I1(level4_in[4591]),
   .I2(level4_in[4592]),
   .I3(level4_in[4593]),
   .I4(level4_in[4594]),
   .I5(level4_in[4595])
);

LUT6 #(
   .INIT(64'he7d960c0e7d960c0)  
) LUT6_inst8542 (
   .O(to_level3[766]),
   .I0(level4_in[4596]),
   .I1(level4_in[4597]),
   .I2(level4_in[4598]),
   .I3(level4_in[4599]),
   .I4(level4_in[4600]),
   .I5(level4_in[4601])
);

LUT6 #(
   .INIT(64'h57d3d40c57d3d40c)  
) LUT6_inst8543 (
   .O(to_level3[767]),
   .I0(level4_in[4602]),
   .I1(level4_in[4603]),
   .I2(level4_in[4604]),
   .I3(level4_in[4605]),
   .I4(level4_in[4606]),
   .I5(level4_in[4607])
);

LUT6 #(
   .INIT(64'h9fdbb59d9fdbb59d)  
) LUT6_inst8544 (
   .O(to_level3[768]),
   .I0(level4_in[4608]),
   .I1(level4_in[4609]),
   .I2(level4_in[4610]),
   .I3(level4_in[4611]),
   .I4(level4_in[4612]),
   .I5(level4_in[4613])
);

LUT6 #(
   .INIT(64'ha227c8eaa227c8ea)  
) LUT6_inst8545 (
   .O(to_level3[769]),
   .I0(level4_in[4614]),
   .I1(level4_in[4615]),
   .I2(level4_in[4616]),
   .I3(level4_in[4617]),
   .I4(level4_in[4618]),
   .I5(level4_in[4619])
);

LUT6 #(
   .INIT(64'h366815e8366815e8)  
) LUT6_inst8546 (
   .O(to_level3[770]),
   .I0(level4_in[4620]),
   .I1(level4_in[4621]),
   .I2(level4_in[4622]),
   .I3(level4_in[4623]),
   .I4(level4_in[4624]),
   .I5(level4_in[4625])
);

LUT6 #(
   .INIT(64'h8b3bbba68b3bbba6)  
) LUT6_inst8547 (
   .O(to_level3[771]),
   .I0(level4_in[4626]),
   .I1(level4_in[4627]),
   .I2(level4_in[4628]),
   .I3(level4_in[4629]),
   .I4(level4_in[4630]),
   .I5(level4_in[4631])
);

LUT6 #(
   .INIT(64'h5759633457596334)  
) LUT6_inst8548 (
   .O(to_level3[772]),
   .I0(level4_in[4632]),
   .I1(level4_in[4633]),
   .I2(level4_in[4634]),
   .I3(level4_in[4635]),
   .I4(level4_in[4636]),
   .I5(level4_in[4637])
);

LUT6 #(
   .INIT(64'h010c96b3010c96b3)  
) LUT6_inst8549 (
   .O(to_level3[773]),
   .I0(level4_in[4638]),
   .I1(level4_in[4639]),
   .I2(level4_in[4640]),
   .I3(level4_in[4641]),
   .I4(level4_in[4642]),
   .I5(level4_in[4643])
);

LUT6 #(
   .INIT(64'hf8d69a44f8d69a44)  
) LUT6_inst8550 (
   .O(to_level3[774]),
   .I0(level4_in[4644]),
   .I1(level4_in[4645]),
   .I2(level4_in[4646]),
   .I3(level4_in[4647]),
   .I4(level4_in[4648]),
   .I5(level4_in[4649])
);

LUT6 #(
   .INIT(64'hcc9ac869cc9ac869)  
) LUT6_inst8551 (
   .O(to_level3[775]),
   .I0(level4_in[4650]),
   .I1(level4_in[4651]),
   .I2(level4_in[4652]),
   .I3(level4_in[4653]),
   .I4(level4_in[4654]),
   .I5(level4_in[4655])
);

LUT6 #(
   .INIT(64'h0b769c480b769c48)  
) LUT6_inst8552 (
   .O(to_level3[776]),
   .I0(level4_in[4656]),
   .I1(level4_in[4657]),
   .I2(level4_in[4658]),
   .I3(level4_in[4659]),
   .I4(level4_in[4660]),
   .I5(level4_in[4661])
);

LUT6 #(
   .INIT(64'h7cdb71107cdb7110)  
) LUT6_inst8553 (
   .O(to_level3[777]),
   .I0(level4_in[4662]),
   .I1(level4_in[4663]),
   .I2(level4_in[4664]),
   .I3(level4_in[4665]),
   .I4(level4_in[4666]),
   .I5(level4_in[4667])
);

LUT6 #(
   .INIT(64'h5234d5e25234d5e2)  
) LUT6_inst8554 (
   .O(to_level3[778]),
   .I0(level4_in[4668]),
   .I1(level4_in[4669]),
   .I2(level4_in[4670]),
   .I3(level4_in[4671]),
   .I4(level4_in[4672]),
   .I5(level4_in[4673])
);

LUT6 #(
   .INIT(64'hbdcf7939bdcf7939)  
) LUT6_inst8555 (
   .O(to_level3[779]),
   .I0(level4_in[4674]),
   .I1(level4_in[4675]),
   .I2(level4_in[4676]),
   .I3(level4_in[4677]),
   .I4(level4_in[4678]),
   .I5(level4_in[4679])
);

LUT6 #(
   .INIT(64'hedd0b8b7edd0b8b7)  
) LUT6_inst8556 (
   .O(to_level3[780]),
   .I0(level4_in[4680]),
   .I1(level4_in[4681]),
   .I2(level4_in[4682]),
   .I3(level4_in[4683]),
   .I4(level4_in[4684]),
   .I5(level4_in[4685])
);

LUT6 #(
   .INIT(64'h48aabd7d48aabd7d)  
) LUT6_inst8557 (
   .O(to_level3[781]),
   .I0(level4_in[4686]),
   .I1(level4_in[4687]),
   .I2(level4_in[4688]),
   .I3(level4_in[4689]),
   .I4(level4_in[4690]),
   .I5(level4_in[4691])
);

LUT6 #(
   .INIT(64'hd3e17be3d3e17be3)  
) LUT6_inst8558 (
   .O(to_level3[782]),
   .I0(level4_in[4692]),
   .I1(level4_in[4693]),
   .I2(level4_in[4694]),
   .I3(level4_in[4695]),
   .I4(level4_in[4696]),
   .I5(level4_in[4697])
);

LUT6 #(
   .INIT(64'h3903f9f13903f9f1)  
) LUT6_inst8559 (
   .O(to_level3[783]),
   .I0(level4_in[4698]),
   .I1(level4_in[4699]),
   .I2(level4_in[4700]),
   .I3(level4_in[4701]),
   .I4(level4_in[4702]),
   .I5(level4_in[4703])
);

LUT6 #(
   .INIT(64'h99c48ea699c48ea6)  
) LUT6_inst8560 (
   .O(to_level3[784]),
   .I0(level4_in[4704]),
   .I1(level4_in[4705]),
   .I2(level4_in[4706]),
   .I3(level4_in[4707]),
   .I4(level4_in[4708]),
   .I5(level4_in[4709])
);

LUT6 #(
   .INIT(64'he6da5040e6da5040)  
) LUT6_inst8561 (
   .O(to_level3[785]),
   .I0(level4_in[4710]),
   .I1(level4_in[4711]),
   .I2(level4_in[4712]),
   .I3(level4_in[4713]),
   .I4(level4_in[4714]),
   .I5(level4_in[4715])
);

LUT6 #(
   .INIT(64'h02d7a53e02d7a53e)  
) LUT6_inst8562 (
   .O(to_level3[786]),
   .I0(level4_in[4716]),
   .I1(level4_in[4717]),
   .I2(level4_in[4718]),
   .I3(level4_in[4719]),
   .I4(level4_in[4720]),
   .I5(level4_in[4721])
);

LUT6 #(
   .INIT(64'h42c0168c42c0168c)  
) LUT6_inst8563 (
   .O(to_level3[787]),
   .I0(level4_in[4722]),
   .I1(level4_in[4723]),
   .I2(level4_in[4724]),
   .I3(level4_in[4725]),
   .I4(level4_in[4726]),
   .I5(level4_in[4727])
);

LUT6 #(
   .INIT(64'hb3bcc4ffb3bcc4ff)  
) LUT6_inst8564 (
   .O(to_level3[788]),
   .I0(level4_in[4728]),
   .I1(level4_in[4729]),
   .I2(level4_in[4730]),
   .I3(level4_in[4731]),
   .I4(level4_in[4732]),
   .I5(level4_in[4733])
);

LUT6 #(
   .INIT(64'hed38fdb0ed38fdb0)  
) LUT6_inst8565 (
   .O(to_level3[789]),
   .I0(level4_in[4734]),
   .I1(level4_in[4735]),
   .I2(level4_in[4736]),
   .I3(level4_in[4737]),
   .I4(level4_in[4738]),
   .I5(level4_in[4739])
);

LUT6 #(
   .INIT(64'hb03c78afb03c78af)  
) LUT6_inst8566 (
   .O(to_level3[790]),
   .I0(level4_in[4740]),
   .I1(level4_in[4741]),
   .I2(level4_in[4742]),
   .I3(level4_in[4743]),
   .I4(level4_in[4744]),
   .I5(level4_in[4745])
);

LUT6 #(
   .INIT(64'h16394d8f16394d8f)  
) LUT6_inst8567 (
   .O(to_level3[791]),
   .I0(level4_in[4746]),
   .I1(level4_in[4747]),
   .I2(level4_in[4748]),
   .I3(level4_in[4749]),
   .I4(level4_in[4750]),
   .I5(level4_in[4751])
);

LUT6 #(
   .INIT(64'h15bcb26e15bcb26e)  
) LUT6_inst8568 (
   .O(to_level3[792]),
   .I0(level4_in[4752]),
   .I1(level4_in[4753]),
   .I2(level4_in[4754]),
   .I3(level4_in[4755]),
   .I4(level4_in[4756]),
   .I5(level4_in[4757])
);

LUT6 #(
   .INIT(64'h1eefecea1eefecea)  
) LUT6_inst8569 (
   .O(to_level3[793]),
   .I0(level4_in[4758]),
   .I1(level4_in[4759]),
   .I2(level4_in[4760]),
   .I3(level4_in[4761]),
   .I4(level4_in[4762]),
   .I5(level4_in[4763])
);

LUT6 #(
   .INIT(64'hc4d65ef4c4d65ef4)  
) LUT6_inst8570 (
   .O(to_level3[794]),
   .I0(level4_in[4764]),
   .I1(level4_in[4765]),
   .I2(level4_in[4766]),
   .I3(level4_in[4767]),
   .I4(level4_in[4768]),
   .I5(level4_in[4769])
);

LUT6 #(
   .INIT(64'hf89facaef89facae)  
) LUT6_inst8571 (
   .O(to_level3[795]),
   .I0(level4_in[4770]),
   .I1(level4_in[4771]),
   .I2(level4_in[4772]),
   .I3(level4_in[4773]),
   .I4(level4_in[4774]),
   .I5(level4_in[4775])
);

LUT6 #(
   .INIT(64'hb61621c6b61621c6)  
) LUT6_inst8572 (
   .O(to_level3[796]),
   .I0(level4_in[4776]),
   .I1(level4_in[4777]),
   .I2(level4_in[4778]),
   .I3(level4_in[4779]),
   .I4(level4_in[4780]),
   .I5(level4_in[4781])
);

LUT6 #(
   .INIT(64'h30a613fe30a613fe)  
) LUT6_inst8573 (
   .O(to_level3[797]),
   .I0(level4_in[4782]),
   .I1(level4_in[4783]),
   .I2(level4_in[4784]),
   .I3(level4_in[4785]),
   .I4(level4_in[4786]),
   .I5(level4_in[4787])
);

LUT6 #(
   .INIT(64'h30a3afe230a3afe2)  
) LUT6_inst8574 (
   .O(to_level3[798]),
   .I0(level4_in[4788]),
   .I1(level4_in[4789]),
   .I2(level4_in[4790]),
   .I3(level4_in[4791]),
   .I4(level4_in[4792]),
   .I5(level4_in[4793])
);

LUT6 #(
   .INIT(64'h66cff35766cff357)  
) LUT6_inst8575 (
   .O(to_level3[799]),
   .I0(level4_in[4794]),
   .I1(level4_in[4795]),
   .I2(level4_in[4796]),
   .I3(level4_in[4797]),
   .I4(level4_in[4798]),
   .I5(level4_in[4799])
);

LUT6 #(
   .INIT(64'hc2a8a99cc2a8a99c)  
) LUT6_inst8576 (
   .O(to_level3[800]),
   .I0(level4_in[4800]),
   .I1(level4_in[4801]),
   .I2(level4_in[4802]),
   .I3(level4_in[4803]),
   .I4(level4_in[4804]),
   .I5(level4_in[4805])
);

LUT6 #(
   .INIT(64'h765028c2765028c2)  
) LUT6_inst8577 (
   .O(to_level3[801]),
   .I0(level4_in[4806]),
   .I1(level4_in[4807]),
   .I2(level4_in[4808]),
   .I3(level4_in[4809]),
   .I4(level4_in[4810]),
   .I5(level4_in[4811])
);

LUT6 #(
   .INIT(64'h5c3033f25c3033f2)  
) LUT6_inst8578 (
   .O(to_level3[802]),
   .I0(level4_in[4812]),
   .I1(level4_in[4813]),
   .I2(level4_in[4814]),
   .I3(level4_in[4815]),
   .I4(level4_in[4816]),
   .I5(level4_in[4817])
);

LUT6 #(
   .INIT(64'hf503cf08f503cf08)  
) LUT6_inst8579 (
   .O(to_level3[803]),
   .I0(level4_in[4818]),
   .I1(level4_in[4819]),
   .I2(level4_in[4820]),
   .I3(level4_in[4821]),
   .I4(level4_in[4822]),
   .I5(level4_in[4823])
);

LUT6 #(
   .INIT(64'h8fad936c8fad936c)  
) LUT6_inst8580 (
   .O(to_level3[804]),
   .I0(level4_in[4824]),
   .I1(level4_in[4825]),
   .I2(level4_in[4826]),
   .I3(level4_in[4827]),
   .I4(level4_in[4828]),
   .I5(level4_in[4829])
);

LUT6 #(
   .INIT(64'h086e5250086e5250)  
) LUT6_inst8581 (
   .O(to_level3[805]),
   .I0(level4_in[4830]),
   .I1(level4_in[4831]),
   .I2(level4_in[4832]),
   .I3(level4_in[4833]),
   .I4(level4_in[4834]),
   .I5(level4_in[4835])
);

LUT6 #(
   .INIT(64'h8c6695918c669591)  
) LUT6_inst8582 (
   .O(to_level3[806]),
   .I0(level4_in[4836]),
   .I1(level4_in[4837]),
   .I2(level4_in[4838]),
   .I3(level4_in[4839]),
   .I4(level4_in[4840]),
   .I5(level4_in[4841])
);

LUT6 #(
   .INIT(64'h83d1011683d10116)  
) LUT6_inst8583 (
   .O(to_level3[807]),
   .I0(level4_in[4842]),
   .I1(level4_in[4843]),
   .I2(level4_in[4844]),
   .I3(level4_in[4845]),
   .I4(level4_in[4846]),
   .I5(level4_in[4847])
);

LUT6 #(
   .INIT(64'h6b9db9a46b9db9a4)  
) LUT6_inst8584 (
   .O(to_level3[808]),
   .I0(level4_in[4848]),
   .I1(level4_in[4849]),
   .I2(level4_in[4850]),
   .I3(level4_in[4851]),
   .I4(level4_in[4852]),
   .I5(level4_in[4853])
);

LUT6 #(
   .INIT(64'h3bbc9b663bbc9b66)  
) LUT6_inst8585 (
   .O(to_level3[809]),
   .I0(level4_in[4854]),
   .I1(level4_in[4855]),
   .I2(level4_in[4856]),
   .I3(level4_in[4857]),
   .I4(level4_in[4858]),
   .I5(level4_in[4859])
);

LUT6 #(
   .INIT(64'h499c0e30499c0e30)  
) LUT6_inst8586 (
   .O(to_level3[810]),
   .I0(level4_in[4860]),
   .I1(level4_in[4861]),
   .I2(level4_in[4862]),
   .I3(level4_in[4863]),
   .I4(level4_in[4864]),
   .I5(level4_in[4865])
);

LUT6 #(
   .INIT(64'hf76b99a9f76b99a9)  
) LUT6_inst8587 (
   .O(to_level3[811]),
   .I0(level4_in[4866]),
   .I1(level4_in[4867]),
   .I2(level4_in[4868]),
   .I3(level4_in[4869]),
   .I4(level4_in[4870]),
   .I5(level4_in[4871])
);

LUT6 #(
   .INIT(64'h1d8b96ba1d8b96ba)  
) LUT6_inst8588 (
   .O(to_level3[812]),
   .I0(level4_in[4872]),
   .I1(level4_in[4873]),
   .I2(level4_in[4874]),
   .I3(level4_in[4875]),
   .I4(level4_in[4876]),
   .I5(level4_in[4877])
);

LUT6 #(
   .INIT(64'h9772799897727998)  
) LUT6_inst8589 (
   .O(to_level3[813]),
   .I0(level4_in[4878]),
   .I1(level4_in[4879]),
   .I2(level4_in[4880]),
   .I3(level4_in[4881]),
   .I4(level4_in[4882]),
   .I5(level4_in[4883])
);

LUT6 #(
   .INIT(64'h3652582536525825)  
) LUT6_inst8590 (
   .O(to_level3[814]),
   .I0(level4_in[4884]),
   .I1(level4_in[4885]),
   .I2(level4_in[4886]),
   .I3(level4_in[4887]),
   .I4(level4_in[4888]),
   .I5(level4_in[4889])
);

LUT6 #(
   .INIT(64'h6ff2c70f6ff2c70f)  
) LUT6_inst8591 (
   .O(to_level3[815]),
   .I0(level4_in[4890]),
   .I1(level4_in[4891]),
   .I2(level4_in[4892]),
   .I3(level4_in[4893]),
   .I4(level4_in[4894]),
   .I5(level4_in[4895])
);

LUT6 #(
   .INIT(64'h44d874c544d874c5)  
) LUT6_inst8592 (
   .O(to_level3[816]),
   .I0(level4_in[4896]),
   .I1(level4_in[4897]),
   .I2(level4_in[4898]),
   .I3(level4_in[4899]),
   .I4(level4_in[4900]),
   .I5(level4_in[4901])
);

LUT6 #(
   .INIT(64'he156268de156268d)  
) LUT6_inst8593 (
   .O(to_level3[817]),
   .I0(level4_in[4902]),
   .I1(level4_in[4903]),
   .I2(level4_in[4904]),
   .I3(level4_in[4905]),
   .I4(level4_in[4906]),
   .I5(level4_in[4907])
);

LUT6 #(
   .INIT(64'h4fe71f9b4fe71f9b)  
) LUT6_inst8594 (
   .O(to_level3[818]),
   .I0(level4_in[4908]),
   .I1(level4_in[4909]),
   .I2(level4_in[4910]),
   .I3(level4_in[4911]),
   .I4(level4_in[4912]),
   .I5(level4_in[4913])
);

LUT6 #(
   .INIT(64'h248fac19248fac19)  
) LUT6_inst8595 (
   .O(to_level3[819]),
   .I0(level4_in[4914]),
   .I1(level4_in[4915]),
   .I2(level4_in[4916]),
   .I3(level4_in[4917]),
   .I4(level4_in[4918]),
   .I5(level4_in[4919])
);

LUT6 #(
   .INIT(64'he7601df2e7601df2)  
) LUT6_inst8596 (
   .O(to_level3[820]),
   .I0(level4_in[4920]),
   .I1(level4_in[4921]),
   .I2(level4_in[4922]),
   .I3(level4_in[4923]),
   .I4(level4_in[4924]),
   .I5(level4_in[4925])
);

LUT6 #(
   .INIT(64'he45babb1e45babb1)  
) LUT6_inst8597 (
   .O(to_level3[821]),
   .I0(level4_in[4926]),
   .I1(level4_in[4927]),
   .I2(level4_in[4928]),
   .I3(level4_in[4929]),
   .I4(level4_in[4930]),
   .I5(level4_in[4931])
);

LUT6 #(
   .INIT(64'h77b77d9277b77d92)  
) LUT6_inst8598 (
   .O(to_level3[822]),
   .I0(level4_in[4932]),
   .I1(level4_in[4933]),
   .I2(level4_in[4934]),
   .I3(level4_in[4935]),
   .I4(level4_in[4936]),
   .I5(level4_in[4937])
);

LUT6 #(
   .INIT(64'h954d0afe954d0afe)  
) LUT6_inst8599 (
   .O(to_level3[823]),
   .I0(level4_in[4938]),
   .I1(level4_in[4939]),
   .I2(level4_in[4940]),
   .I3(level4_in[4941]),
   .I4(level4_in[4942]),
   .I5(level4_in[4943])
);

LUT6 #(
   .INIT(64'h266d0f72266d0f72)  
) LUT6_inst8600 (
   .O(to_level3[824]),
   .I0(level4_in[4944]),
   .I1(level4_in[4945]),
   .I2(level4_in[4946]),
   .I3(level4_in[4947]),
   .I4(level4_in[4948]),
   .I5(level4_in[4949])
);

LUT6 #(
   .INIT(64'h94fd628594fd6285)  
) LUT6_inst8601 (
   .O(to_level3[825]),
   .I0(level4_in[4950]),
   .I1(level4_in[4951]),
   .I2(level4_in[4952]),
   .I3(level4_in[4953]),
   .I4(level4_in[4954]),
   .I5(level4_in[4955])
);

LUT6 #(
   .INIT(64'hebb9403cebb9403c)  
) LUT6_inst8602 (
   .O(to_level3[826]),
   .I0(level4_in[4956]),
   .I1(level4_in[4957]),
   .I2(level4_in[4958]),
   .I3(level4_in[4959]),
   .I4(level4_in[4960]),
   .I5(level4_in[4961])
);

LUT6 #(
   .INIT(64'h4bef23584bef2358)  
) LUT6_inst8603 (
   .O(to_level3[827]),
   .I0(level4_in[4962]),
   .I1(level4_in[4963]),
   .I2(level4_in[4964]),
   .I3(level4_in[4965]),
   .I4(level4_in[4966]),
   .I5(level4_in[4967])
);

LUT6 #(
   .INIT(64'h1b74751b1b74751b)  
) LUT6_inst8604 (
   .O(to_level3[828]),
   .I0(level4_in[4968]),
   .I1(level4_in[4969]),
   .I2(level4_in[4970]),
   .I3(level4_in[4971]),
   .I4(level4_in[4972]),
   .I5(level4_in[4973])
);

LUT6 #(
   .INIT(64'h2ffaa56d2ffaa56d)  
) LUT6_inst8605 (
   .O(to_level3[829]),
   .I0(level4_in[4974]),
   .I1(level4_in[4975]),
   .I2(level4_in[4976]),
   .I3(level4_in[4977]),
   .I4(level4_in[4978]),
   .I5(level4_in[4979])
);

LUT6 #(
   .INIT(64'hf0310342f0310342)  
) LUT6_inst8606 (
   .O(to_level3[830]),
   .I0(level4_in[4980]),
   .I1(level4_in[4981]),
   .I2(level4_in[4982]),
   .I3(level4_in[4983]),
   .I4(level4_in[4984]),
   .I5(level4_in[4985])
);

LUT6 #(
   .INIT(64'hf7562a17f7562a17)  
) LUT6_inst8607 (
   .O(to_level3[831]),
   .I0(level4_in[4986]),
   .I1(level4_in[4987]),
   .I2(level4_in[4988]),
   .I3(level4_in[4989]),
   .I4(level4_in[4990]),
   .I5(level4_in[4991])
);

LUT6 #(
   .INIT(64'h36983bc836983bc8)  
) LUT6_inst8608 (
   .O(to_level3[832]),
   .I0(level4_in[4992]),
   .I1(level4_in[4993]),
   .I2(level4_in[4994]),
   .I3(level4_in[4995]),
   .I4(level4_in[4996]),
   .I5(level4_in[4997])
);

LUT6 #(
   .INIT(64'hd9b74f62d9b74f62)  
) LUT6_inst8609 (
   .O(to_level3[833]),
   .I0(level4_in[4998]),
   .I1(level4_in[4999]),
   .I2(level4_in[5000]),
   .I3(level4_in[5001]),
   .I4(level4_in[5002]),
   .I5(level4_in[5003])
);

LUT6 #(
   .INIT(64'h0300c3b10300c3b1)  
) LUT6_inst8610 (
   .O(to_level3[834]),
   .I0(level4_in[5004]),
   .I1(level4_in[5005]),
   .I2(level4_in[5006]),
   .I3(level4_in[5007]),
   .I4(level4_in[5008]),
   .I5(level4_in[5009])
);

LUT6 #(
   .INIT(64'h8231b1de8231b1de)  
) LUT6_inst8611 (
   .O(to_level3[835]),
   .I0(level4_in[5010]),
   .I1(level4_in[5011]),
   .I2(level4_in[5012]),
   .I3(level4_in[5013]),
   .I4(level4_in[5014]),
   .I5(level4_in[5015])
);

LUT6 #(
   .INIT(64'h1148b0481148b048)  
) LUT6_inst8612 (
   .O(to_level3[836]),
   .I0(level4_in[5016]),
   .I1(level4_in[5017]),
   .I2(level4_in[5018]),
   .I3(level4_in[5019]),
   .I4(level4_in[5020]),
   .I5(level4_in[5021])
);

LUT6 #(
   .INIT(64'h30d8bcb430d8bcb4)  
) LUT6_inst8613 (
   .O(to_level3[837]),
   .I0(level4_in[5022]),
   .I1(level4_in[5023]),
   .I2(level4_in[5024]),
   .I3(level4_in[5025]),
   .I4(level4_in[5026]),
   .I5(level4_in[5027])
);

LUT6 #(
   .INIT(64'hca427f2aca427f2a)  
) LUT6_inst8614 (
   .O(to_level3[838]),
   .I0(level4_in[5028]),
   .I1(level4_in[5029]),
   .I2(level4_in[5030]),
   .I3(level4_in[5031]),
   .I4(level4_in[5032]),
   .I5(level4_in[5033])
);

LUT6 #(
   .INIT(64'hfe491d36fe491d36)  
) LUT6_inst8615 (
   .O(to_level3[839]),
   .I0(level4_in[5034]),
   .I1(level4_in[5035]),
   .I2(level4_in[5036]),
   .I3(level4_in[5037]),
   .I4(level4_in[5038]),
   .I5(level4_in[5039])
);

LUT6 #(
   .INIT(64'h5e6e205e5e6e205e)  
) LUT6_inst8616 (
   .O(to_level3[840]),
   .I0(level4_in[5040]),
   .I1(level4_in[5041]),
   .I2(level4_in[5042]),
   .I3(level4_in[5043]),
   .I4(level4_in[5044]),
   .I5(level4_in[5045])
);

LUT6 #(
   .INIT(64'hcb6f3664cb6f3664)  
) LUT6_inst8617 (
   .O(to_level3[841]),
   .I0(level4_in[5046]),
   .I1(level4_in[5047]),
   .I2(level4_in[5048]),
   .I3(level4_in[5049]),
   .I4(level4_in[5050]),
   .I5(level4_in[5051])
);

LUT6 #(
   .INIT(64'hf3727351f3727351)  
) LUT6_inst8618 (
   .O(to_level3[842]),
   .I0(level4_in[5052]),
   .I1(level4_in[5053]),
   .I2(level4_in[5054]),
   .I3(level4_in[5055]),
   .I4(level4_in[5056]),
   .I5(level4_in[5057])
);

LUT6 #(
   .INIT(64'h96e551ab96e551ab)  
) LUT6_inst8619 (
   .O(to_level3[843]),
   .I0(level4_in[5058]),
   .I1(level4_in[5059]),
   .I2(level4_in[5060]),
   .I3(level4_in[5061]),
   .I4(level4_in[5062]),
   .I5(level4_in[5063])
);

LUT6 #(
   .INIT(64'he9243b71e9243b71)  
) LUT6_inst8620 (
   .O(to_level3[844]),
   .I0(level4_in[5064]),
   .I1(level4_in[5065]),
   .I2(level4_in[5066]),
   .I3(level4_in[5067]),
   .I4(level4_in[5068]),
   .I5(level4_in[5069])
);

LUT6 #(
   .INIT(64'h68e89c6a68e89c6a)  
) LUT6_inst8621 (
   .O(to_level3[845]),
   .I0(level4_in[5070]),
   .I1(level4_in[5071]),
   .I2(level4_in[5072]),
   .I3(level4_in[5073]),
   .I4(level4_in[5074]),
   .I5(level4_in[5075])
);

LUT6 #(
   .INIT(64'h8695feb28695feb2)  
) LUT6_inst8622 (
   .O(to_level3[846]),
   .I0(level4_in[5076]),
   .I1(level4_in[5077]),
   .I2(level4_in[5078]),
   .I3(level4_in[5079]),
   .I4(level4_in[5080]),
   .I5(level4_in[5081])
);

LUT6 #(
   .INIT(64'hadb8228eadb8228e)  
) LUT6_inst8623 (
   .O(to_level3[847]),
   .I0(level4_in[5082]),
   .I1(level4_in[5083]),
   .I2(level4_in[5084]),
   .I3(level4_in[5085]),
   .I4(level4_in[5086]),
   .I5(level4_in[5087])
);

LUT6 #(
   .INIT(64'hb32c6e2eb32c6e2e)  
) LUT6_inst8624 (
   .O(to_level3[848]),
   .I0(level4_in[5088]),
   .I1(level4_in[5089]),
   .I2(level4_in[5090]),
   .I3(level4_in[5091]),
   .I4(level4_in[5092]),
   .I5(level4_in[5093])
);

LUT6 #(
   .INIT(64'hff2d4970ff2d4970)  
) LUT6_inst8625 (
   .O(to_level3[849]),
   .I0(level4_in[5094]),
   .I1(level4_in[5095]),
   .I2(level4_in[5096]),
   .I3(level4_in[5097]),
   .I4(level4_in[5098]),
   .I5(level4_in[5099])
);

LUT6 #(
   .INIT(64'ha10dafcba10dafcb)  
) LUT6_inst8626 (
   .O(to_level3[850]),
   .I0(level4_in[5100]),
   .I1(level4_in[5101]),
   .I2(level4_in[5102]),
   .I3(level4_in[5103]),
   .I4(level4_in[5104]),
   .I5(level4_in[5105])
);

LUT6 #(
   .INIT(64'hbfc2b536bfc2b536)  
) LUT6_inst8627 (
   .O(to_level3[851]),
   .I0(level4_in[5106]),
   .I1(level4_in[5107]),
   .I2(level4_in[5108]),
   .I3(level4_in[5109]),
   .I4(level4_in[5110]),
   .I5(level4_in[5111])
);

LUT6 #(
   .INIT(64'h1998e8d61998e8d6)  
) LUT6_inst8628 (
   .O(to_level3[852]),
   .I0(level4_in[5112]),
   .I1(level4_in[5113]),
   .I2(level4_in[5114]),
   .I3(level4_in[5115]),
   .I4(level4_in[5116]),
   .I5(level4_in[5117])
);

LUT6 #(
   .INIT(64'h9f937a779f937a77)  
) LUT6_inst8629 (
   .O(to_level3[853]),
   .I0(level4_in[5118]),
   .I1(level4_in[5119]),
   .I2(level4_in[5120]),
   .I3(level4_in[5121]),
   .I4(level4_in[5122]),
   .I5(level4_in[5123])
);

LUT6 #(
   .INIT(64'h7d7bf6df7d7bf6df)  
) LUT6_inst8630 (
   .O(to_level3[854]),
   .I0(level4_in[5124]),
   .I1(level4_in[5125]),
   .I2(level4_in[5126]),
   .I3(level4_in[5127]),
   .I4(level4_in[5128]),
   .I5(level4_in[5129])
);

LUT6 #(
   .INIT(64'h6fa020dd6fa020dd)  
) LUT6_inst8631 (
   .O(to_level3[855]),
   .I0(level4_in[5130]),
   .I1(level4_in[5131]),
   .I2(level4_in[5132]),
   .I3(level4_in[5133]),
   .I4(level4_in[5134]),
   .I5(level4_in[5135])
);

LUT6 #(
   .INIT(64'h3ed55bdf3ed55bdf)  
) LUT6_inst8632 (
   .O(to_level3[856]),
   .I0(level4_in[5136]),
   .I1(level4_in[5137]),
   .I2(level4_in[5138]),
   .I3(level4_in[5139]),
   .I4(level4_in[5140]),
   .I5(level4_in[5141])
);

LUT6 #(
   .INIT(64'h81ddfef481ddfef4)  
) LUT6_inst8633 (
   .O(to_level3[857]),
   .I0(level4_in[5142]),
   .I1(level4_in[5143]),
   .I2(level4_in[5144]),
   .I3(level4_in[5145]),
   .I4(level4_in[5146]),
   .I5(level4_in[5147])
);

LUT6 #(
   .INIT(64'h7b3903357b390335)  
) LUT6_inst8634 (
   .O(to_level3[858]),
   .I0(level4_in[5148]),
   .I1(level4_in[5149]),
   .I2(level4_in[5150]),
   .I3(level4_in[5151]),
   .I4(level4_in[5152]),
   .I5(level4_in[5153])
);

LUT6 #(
   .INIT(64'h8a29f8918a29f891)  
) LUT6_inst8635 (
   .O(to_level3[859]),
   .I0(level4_in[5154]),
   .I1(level4_in[5155]),
   .I2(level4_in[5156]),
   .I3(level4_in[5157]),
   .I4(level4_in[5158]),
   .I5(level4_in[5159])
);

LUT6 #(
   .INIT(64'ha0dd2541a0dd2541)  
) LUT6_inst8636 (
   .O(to_level3[860]),
   .I0(level4_in[5160]),
   .I1(level4_in[5161]),
   .I2(level4_in[5162]),
   .I3(level4_in[5163]),
   .I4(level4_in[5164]),
   .I5(level4_in[5165])
);

LUT6 #(
   .INIT(64'h15f9239f15f9239f)  
) LUT6_inst8637 (
   .O(to_level3[861]),
   .I0(level4_in[5166]),
   .I1(level4_in[5167]),
   .I2(level4_in[5168]),
   .I3(level4_in[5169]),
   .I4(level4_in[5170]),
   .I5(level4_in[5171])
);

LUT6 #(
   .INIT(64'h22bf960b22bf960b)  
) LUT6_inst8638 (
   .O(to_level3[862]),
   .I0(level4_in[5172]),
   .I1(level4_in[5173]),
   .I2(level4_in[5174]),
   .I3(level4_in[5175]),
   .I4(level4_in[5176]),
   .I5(level4_in[5177])
);

LUT6 #(
   .INIT(64'h25b3846525b38465)  
) LUT6_inst8639 (
   .O(to_level3[863]),
   .I0(level4_in[5178]),
   .I1(level4_in[5179]),
   .I2(level4_in[5180]),
   .I3(level4_in[5181]),
   .I4(level4_in[5182]),
   .I5(level4_in[5183])
);

LUT6 #(
   .INIT(64'hf3c6776df3c6776d)  
) LUT6_inst8640 (
   .O(to_level3[864]),
   .I0(level4_in[5184]),
   .I1(level4_in[5185]),
   .I2(level4_in[5186]),
   .I3(level4_in[5187]),
   .I4(level4_in[5188]),
   .I5(level4_in[5189])
);

LUT6 #(
   .INIT(64'he58438c5e58438c5)  
) LUT6_inst8641 (
   .O(to_level3[865]),
   .I0(level4_in[5190]),
   .I1(level4_in[5191]),
   .I2(level4_in[5192]),
   .I3(level4_in[5193]),
   .I4(level4_in[5194]),
   .I5(level4_in[5195])
);

LUT6 #(
   .INIT(64'h5403005054030050)  
) LUT6_inst8642 (
   .O(to_level3[866]),
   .I0(level4_in[5196]),
   .I1(level4_in[5197]),
   .I2(level4_in[5198]),
   .I3(level4_in[5199]),
   .I4(level4_in[5200]),
   .I5(level4_in[5201])
);

LUT6 #(
   .INIT(64'h5dffac325dffac32)  
) LUT6_inst8643 (
   .O(to_level3[867]),
   .I0(level4_in[5202]),
   .I1(level4_in[5203]),
   .I2(level4_in[5204]),
   .I3(level4_in[5205]),
   .I4(level4_in[5206]),
   .I5(level4_in[5207])
);

LUT6 #(
   .INIT(64'h1683f4231683f423)  
) LUT6_inst8644 (
   .O(to_level3[868]),
   .I0(level4_in[5208]),
   .I1(level4_in[5209]),
   .I2(level4_in[5210]),
   .I3(level4_in[5211]),
   .I4(level4_in[5212]),
   .I5(level4_in[5213])
);

LUT6 #(
   .INIT(64'hb265dceab265dcea)  
) LUT6_inst8645 (
   .O(to_level3[869]),
   .I0(level4_in[5214]),
   .I1(level4_in[5215]),
   .I2(level4_in[5216]),
   .I3(level4_in[5217]),
   .I4(level4_in[5218]),
   .I5(level4_in[5219])
);

LUT6 #(
   .INIT(64'hcb945229cb945229)  
) LUT6_inst8646 (
   .O(to_level3[870]),
   .I0(level4_in[5220]),
   .I1(level4_in[5221]),
   .I2(level4_in[5222]),
   .I3(level4_in[5223]),
   .I4(level4_in[5224]),
   .I5(level4_in[5225])
);

LUT6 #(
   .INIT(64'h590d17e3590d17e3)  
) LUT6_inst8647 (
   .O(to_level3[871]),
   .I0(level4_in[5226]),
   .I1(level4_in[5227]),
   .I2(level4_in[5228]),
   .I3(level4_in[5229]),
   .I4(level4_in[5230]),
   .I5(level4_in[5231])
);

LUT6 #(
   .INIT(64'hdef30b6ddef30b6d)  
) LUT6_inst8648 (
   .O(to_level3[872]),
   .I0(level4_in[5232]),
   .I1(level4_in[5233]),
   .I2(level4_in[5234]),
   .I3(level4_in[5235]),
   .I4(level4_in[5236]),
   .I5(level4_in[5237])
);

LUT6 #(
   .INIT(64'h57f07e4357f07e43)  
) LUT6_inst8649 (
   .O(to_level3[873]),
   .I0(level4_in[5238]),
   .I1(level4_in[5239]),
   .I2(level4_in[5240]),
   .I3(level4_in[5241]),
   .I4(level4_in[5242]),
   .I5(level4_in[5243])
);

LUT6 #(
   .INIT(64'h9a115e509a115e50)  
) LUT6_inst8650 (
   .O(to_level3[874]),
   .I0(level4_in[5244]),
   .I1(level4_in[5245]),
   .I2(level4_in[5246]),
   .I3(level4_in[5247]),
   .I4(level4_in[5248]),
   .I5(level4_in[5249])
);

LUT6 #(
   .INIT(64'hc676fc39c676fc39)  
) LUT6_inst8651 (
   .O(to_level3[875]),
   .I0(level4_in[5250]),
   .I1(level4_in[5251]),
   .I2(level4_in[5252]),
   .I3(level4_in[5253]),
   .I4(level4_in[5254]),
   .I5(level4_in[5255])
);

LUT6 #(
   .INIT(64'h7ac2b0257ac2b025)  
) LUT6_inst8652 (
   .O(to_level3[876]),
   .I0(level4_in[5256]),
   .I1(level4_in[5257]),
   .I2(level4_in[5258]),
   .I3(level4_in[5259]),
   .I4(level4_in[5260]),
   .I5(level4_in[5261])
);

LUT6 #(
   .INIT(64'hd7f7301bd7f7301b)  
) LUT6_inst8653 (
   .O(to_level3[877]),
   .I0(level4_in[5262]),
   .I1(level4_in[5263]),
   .I2(level4_in[5264]),
   .I3(level4_in[5265]),
   .I4(level4_in[5266]),
   .I5(level4_in[5267])
);

LUT6 #(
   .INIT(64'hfcd458b4fcd458b4)  
) LUT6_inst8654 (
   .O(to_level3[878]),
   .I0(level4_in[5268]),
   .I1(level4_in[5269]),
   .I2(level4_in[5270]),
   .I3(level4_in[5271]),
   .I4(level4_in[5272]),
   .I5(level4_in[5273])
);

LUT6 #(
   .INIT(64'h0d3136ba0d3136ba)  
) LUT6_inst8655 (
   .O(to_level3[879]),
   .I0(level4_in[5274]),
   .I1(level4_in[5275]),
   .I2(level4_in[5276]),
   .I3(level4_in[5277]),
   .I4(level4_in[5278]),
   .I5(level4_in[5279])
);

LUT6 #(
   .INIT(64'h11c9a60c11c9a60c)  
) LUT6_inst8656 (
   .O(to_level3[880]),
   .I0(level4_in[5280]),
   .I1(level4_in[5281]),
   .I2(level4_in[5282]),
   .I3(level4_in[5283]),
   .I4(level4_in[5284]),
   .I5(level4_in[5285])
);

LUT6 #(
   .INIT(64'h5c77d2525c77d252)  
) LUT6_inst8657 (
   .O(to_level3[881]),
   .I0(level4_in[5286]),
   .I1(level4_in[5287]),
   .I2(level4_in[5288]),
   .I3(level4_in[5289]),
   .I4(level4_in[5290]),
   .I5(level4_in[5291])
);

LUT6 #(
   .INIT(64'h336351f7336351f7)  
) LUT6_inst8658 (
   .O(to_level3[882]),
   .I0(level4_in[5292]),
   .I1(level4_in[5293]),
   .I2(level4_in[5294]),
   .I3(level4_in[5295]),
   .I4(level4_in[5296]),
   .I5(level4_in[5297])
);

LUT6 #(
   .INIT(64'h0d936cff0d936cff)  
) LUT6_inst8659 (
   .O(to_level3[883]),
   .I0(level4_in[5298]),
   .I1(level4_in[5299]),
   .I2(level4_in[5300]),
   .I3(level4_in[5301]),
   .I4(level4_in[5302]),
   .I5(level4_in[5303])
);

LUT6 #(
   .INIT(64'h335c4fa7335c4fa7)  
) LUT6_inst8660 (
   .O(to_level3[884]),
   .I0(level4_in[5304]),
   .I1(level4_in[5305]),
   .I2(level4_in[5306]),
   .I3(level4_in[5307]),
   .I4(level4_in[5308]),
   .I5(level4_in[5309])
);

LUT6 #(
   .INIT(64'h3b1aa52c3b1aa52c)  
) LUT6_inst8661 (
   .O(to_level3[885]),
   .I0(level4_in[5310]),
   .I1(level4_in[5311]),
   .I2(level4_in[5312]),
   .I3(level4_in[5313]),
   .I4(level4_in[5314]),
   .I5(level4_in[5315])
);

LUT6 #(
   .INIT(64'hddc20e9fddc20e9f)  
) LUT6_inst8662 (
   .O(to_level3[886]),
   .I0(level4_in[5316]),
   .I1(level4_in[5317]),
   .I2(level4_in[5318]),
   .I3(level4_in[5319]),
   .I4(level4_in[5320]),
   .I5(level4_in[5321])
);

LUT6 #(
   .INIT(64'had5bc877ad5bc877)  
) LUT6_inst8663 (
   .O(to_level3[887]),
   .I0(level4_in[5322]),
   .I1(level4_in[5323]),
   .I2(level4_in[5324]),
   .I3(level4_in[5325]),
   .I4(level4_in[5326]),
   .I5(level4_in[5327])
);

LUT6 #(
   .INIT(64'h772d9faf772d9faf)  
) LUT6_inst8664 (
   .O(to_level3[888]),
   .I0(level4_in[5328]),
   .I1(level4_in[5329]),
   .I2(level4_in[5330]),
   .I3(level4_in[5331]),
   .I4(level4_in[5332]),
   .I5(level4_in[5333])
);

LUT6 #(
   .INIT(64'hffb6bc51ffb6bc51)  
) LUT6_inst8665 (
   .O(to_level3[889]),
   .I0(level4_in[5334]),
   .I1(level4_in[5335]),
   .I2(level4_in[5336]),
   .I3(level4_in[5337]),
   .I4(level4_in[5338]),
   .I5(level4_in[5339])
);

LUT6 #(
   .INIT(64'h8c7fc2498c7fc249)  
) LUT6_inst8666 (
   .O(to_level3[890]),
   .I0(level4_in[5340]),
   .I1(level4_in[5341]),
   .I2(level4_in[5342]),
   .I3(level4_in[5343]),
   .I4(level4_in[5344]),
   .I5(level4_in[5345])
);

LUT6 #(
   .INIT(64'hee972484ee972484)  
) LUT6_inst8667 (
   .O(to_level3[891]),
   .I0(level4_in[5346]),
   .I1(level4_in[5347]),
   .I2(level4_in[5348]),
   .I3(level4_in[5349]),
   .I4(level4_in[5350]),
   .I5(level4_in[5351])
);

LUT6 #(
   .INIT(64'h70593b8270593b82)  
) LUT6_inst8668 (
   .O(to_level3[892]),
   .I0(level4_in[5352]),
   .I1(level4_in[5353]),
   .I2(level4_in[5354]),
   .I3(level4_in[5355]),
   .I4(level4_in[5356]),
   .I5(level4_in[5357])
);

LUT6 #(
   .INIT(64'h3ebeb8ce3ebeb8ce)  
) LUT6_inst8669 (
   .O(to_level3[893]),
   .I0(level4_in[5358]),
   .I1(level4_in[5359]),
   .I2(level4_in[5360]),
   .I3(level4_in[5361]),
   .I4(level4_in[5362]),
   .I5(level4_in[5363])
);

LUT6 #(
   .INIT(64'h0e3781450e378145)  
) LUT6_inst8670 (
   .O(to_level3[894]),
   .I0(level4_in[5364]),
   .I1(level4_in[5365]),
   .I2(level4_in[5366]),
   .I3(level4_in[5367]),
   .I4(level4_in[5368]),
   .I5(level4_in[5369])
);

LUT6 #(
   .INIT(64'h09fe1c6d09fe1c6d)  
) LUT6_inst8671 (
   .O(to_level3[895]),
   .I0(level4_in[5370]),
   .I1(level4_in[5371]),
   .I2(level4_in[5372]),
   .I3(level4_in[5373]),
   .I4(level4_in[5374]),
   .I5(level4_in[5375])
);

LUT6 #(
   .INIT(64'h356a7783356a7783)  
) LUT6_inst8672 (
   .O(to_level3[896]),
   .I0(level4_in[5376]),
   .I1(level4_in[5377]),
   .I2(level4_in[5378]),
   .I3(level4_in[5379]),
   .I4(level4_in[5380]),
   .I5(level4_in[5381])
);

LUT6 #(
   .INIT(64'hd5d21c25d5d21c25)  
) LUT6_inst8673 (
   .O(to_level3[897]),
   .I0(level4_in[5382]),
   .I1(level4_in[5383]),
   .I2(level4_in[5384]),
   .I3(level4_in[5385]),
   .I4(level4_in[5386]),
   .I5(level4_in[5387])
);

LUT6 #(
   .INIT(64'h6942f2076942f207)  
) LUT6_inst8674 (
   .O(to_level3[898]),
   .I0(level4_in[5388]),
   .I1(level4_in[5389]),
   .I2(level4_in[5390]),
   .I3(level4_in[5391]),
   .I4(level4_in[5392]),
   .I5(level4_in[5393])
);

LUT6 #(
   .INIT(64'h7058c95e7058c95e)  
) LUT6_inst8675 (
   .O(to_level3[899]),
   .I0(level4_in[5394]),
   .I1(level4_in[5395]),
   .I2(level4_in[5396]),
   .I3(level4_in[5397]),
   .I4(level4_in[5398]),
   .I5(level4_in[5399])
);

LUT6 #(
   .INIT(64'hb85858f8b85858f8)  
) LUT6_inst8676 (
   .O(to_level3[900]),
   .I0(level4_in[5400]),
   .I1(level4_in[5401]),
   .I2(level4_in[5402]),
   .I3(level4_in[5403]),
   .I4(level4_in[5404]),
   .I5(level4_in[5405])
);

LUT6 #(
   .INIT(64'hb94ecc1cb94ecc1c)  
) LUT6_inst8677 (
   .O(to_level3[901]),
   .I0(level4_in[5406]),
   .I1(level4_in[5407]),
   .I2(level4_in[5408]),
   .I3(level4_in[5409]),
   .I4(level4_in[5410]),
   .I5(level4_in[5411])
);

LUT6 #(
   .INIT(64'hbb6668b9bb6668b9)  
) LUT6_inst8678 (
   .O(to_level3[902]),
   .I0(level4_in[5412]),
   .I1(level4_in[5413]),
   .I2(level4_in[5414]),
   .I3(level4_in[5415]),
   .I4(level4_in[5416]),
   .I5(level4_in[5417])
);

LUT6 #(
   .INIT(64'hcc361868cc361868)  
) LUT6_inst8679 (
   .O(to_level3[903]),
   .I0(level4_in[5418]),
   .I1(level4_in[5419]),
   .I2(level4_in[5420]),
   .I3(level4_in[5421]),
   .I4(level4_in[5422]),
   .I5(level4_in[5423])
);

LUT6 #(
   .INIT(64'h2485741c2485741c)  
) LUT6_inst8680 (
   .O(to_level3[904]),
   .I0(level4_in[5424]),
   .I1(level4_in[5425]),
   .I2(level4_in[5426]),
   .I3(level4_in[5427]),
   .I4(level4_in[5428]),
   .I5(level4_in[5429])
);

LUT6 #(
   .INIT(64'hf9a97c2df9a97c2d)  
) LUT6_inst8681 (
   .O(to_level3[905]),
   .I0(level4_in[5430]),
   .I1(level4_in[5431]),
   .I2(level4_in[5432]),
   .I3(level4_in[5433]),
   .I4(level4_in[5434]),
   .I5(level4_in[5435])
);

LUT6 #(
   .INIT(64'h5984ba785984ba78)  
) LUT6_inst8682 (
   .O(to_level3[906]),
   .I0(level4_in[5436]),
   .I1(level4_in[5437]),
   .I2(level4_in[5438]),
   .I3(level4_in[5439]),
   .I4(level4_in[5440]),
   .I5(level4_in[5441])
);

LUT6 #(
   .INIT(64'h9147748f9147748f)  
) LUT6_inst8683 (
   .O(to_level3[907]),
   .I0(level4_in[5442]),
   .I1(level4_in[5443]),
   .I2(level4_in[5444]),
   .I3(level4_in[5445]),
   .I4(level4_in[5446]),
   .I5(level4_in[5447])
);

LUT6 #(
   .INIT(64'heba221e0eba221e0)  
) LUT6_inst8684 (
   .O(to_level3[908]),
   .I0(level4_in[5448]),
   .I1(level4_in[5449]),
   .I2(level4_in[5450]),
   .I3(level4_in[5451]),
   .I4(level4_in[5452]),
   .I5(level4_in[5453])
);

LUT6 #(
   .INIT(64'hfce980c7fce980c7)  
) LUT6_inst8685 (
   .O(to_level3[909]),
   .I0(level4_in[5454]),
   .I1(level4_in[5455]),
   .I2(level4_in[5456]),
   .I3(level4_in[5457]),
   .I4(level4_in[5458]),
   .I5(level4_in[5459])
);

LUT6 #(
   .INIT(64'h921aaf45921aaf45)  
) LUT6_inst8686 (
   .O(to_level3[910]),
   .I0(level4_in[5460]),
   .I1(level4_in[5461]),
   .I2(level4_in[5462]),
   .I3(level4_in[5463]),
   .I4(level4_in[5464]),
   .I5(level4_in[5465])
);

LUT6 #(
   .INIT(64'hc9b61b9cc9b61b9c)  
) LUT6_inst8687 (
   .O(to_level3[911]),
   .I0(level4_in[5466]),
   .I1(level4_in[5467]),
   .I2(level4_in[5468]),
   .I3(level4_in[5469]),
   .I4(level4_in[5470]),
   .I5(level4_in[5471])
);

LUT6 #(
   .INIT(64'h78eb476878eb4768)  
) LUT6_inst8688 (
   .O(to_level3[912]),
   .I0(level4_in[5472]),
   .I1(level4_in[5473]),
   .I2(level4_in[5474]),
   .I3(level4_in[5475]),
   .I4(level4_in[5476]),
   .I5(level4_in[5477])
);

LUT6 #(
   .INIT(64'h0150ec3e0150ec3e)  
) LUT6_inst8689 (
   .O(to_level3[913]),
   .I0(level4_in[5478]),
   .I1(level4_in[5479]),
   .I2(level4_in[5480]),
   .I3(level4_in[5481]),
   .I4(level4_in[5482]),
   .I5(level4_in[5483])
);

LUT6 #(
   .INIT(64'h1f135e291f135e29)  
) LUT6_inst8690 (
   .O(to_level3[914]),
   .I0(level4_in[5484]),
   .I1(level4_in[5485]),
   .I2(level4_in[5486]),
   .I3(level4_in[5487]),
   .I4(level4_in[5488]),
   .I5(level4_in[5489])
);

LUT6 #(
   .INIT(64'h571bc97d571bc97d)  
) LUT6_inst8691 (
   .O(to_level3[915]),
   .I0(level4_in[5490]),
   .I1(level4_in[5491]),
   .I2(level4_in[5492]),
   .I3(level4_in[5493]),
   .I4(level4_in[5494]),
   .I5(level4_in[5495])
);

LUT6 #(
   .INIT(64'h9fd87b8d9fd87b8d)  
) LUT6_inst8692 (
   .O(to_level3[916]),
   .I0(level4_in[5496]),
   .I1(level4_in[5497]),
   .I2(level4_in[5498]),
   .I3(level4_in[5499]),
   .I4(level4_in[5500]),
   .I5(level4_in[5501])
);

LUT6 #(
   .INIT(64'hdfea36d9dfea36d9)  
) LUT6_inst8693 (
   .O(to_level3[917]),
   .I0(level4_in[5502]),
   .I1(level4_in[5503]),
   .I2(level4_in[5504]),
   .I3(level4_in[5505]),
   .I4(level4_in[5506]),
   .I5(level4_in[5507])
);

LUT6 #(
   .INIT(64'haea5ddfdaea5ddfd)  
) LUT6_inst8694 (
   .O(to_level3[918]),
   .I0(level4_in[5508]),
   .I1(level4_in[5509]),
   .I2(level4_in[5510]),
   .I3(level4_in[5511]),
   .I4(level4_in[5512]),
   .I5(level4_in[5513])
);

LUT6 #(
   .INIT(64'h7979fcc57979fcc5)  
) LUT6_inst8695 (
   .O(to_level3[919]),
   .I0(level4_in[5514]),
   .I1(level4_in[5515]),
   .I2(level4_in[5516]),
   .I3(level4_in[5517]),
   .I4(level4_in[5518]),
   .I5(level4_in[5519])
);

LUT6 #(
   .INIT(64'h0c70061c0c70061c)  
) LUT6_inst8696 (
   .O(to_level3[920]),
   .I0(level4_in[5520]),
   .I1(level4_in[5521]),
   .I2(level4_in[5522]),
   .I3(level4_in[5523]),
   .I4(level4_in[5524]),
   .I5(level4_in[5525])
);

LUT6 #(
   .INIT(64'h08a4b5b608a4b5b6)  
) LUT6_inst8697 (
   .O(to_level3[921]),
   .I0(level4_in[5526]),
   .I1(level4_in[5527]),
   .I2(level4_in[5528]),
   .I3(level4_in[5529]),
   .I4(level4_in[5530]),
   .I5(level4_in[5531])
);

LUT6 #(
   .INIT(64'h2985966229859662)  
) LUT6_inst8698 (
   .O(to_level3[922]),
   .I0(level4_in[5532]),
   .I1(level4_in[5533]),
   .I2(level4_in[5534]),
   .I3(level4_in[5535]),
   .I4(level4_in[5536]),
   .I5(level4_in[5537])
);

LUT6 #(
   .INIT(64'h7142d23a7142d23a)  
) LUT6_inst8699 (
   .O(to_level3[923]),
   .I0(level4_in[5538]),
   .I1(level4_in[5539]),
   .I2(level4_in[5540]),
   .I3(level4_in[5541]),
   .I4(level4_in[5542]),
   .I5(level4_in[5543])
);

LUT6 #(
   .INIT(64'hc413d1d7c413d1d7)  
) LUT6_inst8700 (
   .O(to_level3[924]),
   .I0(level4_in[5544]),
   .I1(level4_in[5545]),
   .I2(level4_in[5546]),
   .I3(level4_in[5547]),
   .I4(level4_in[5548]),
   .I5(level4_in[5549])
);

LUT6 #(
   .INIT(64'ha3438d04a3438d04)  
) LUT6_inst8701 (
   .O(to_level3[925]),
   .I0(level4_in[5550]),
   .I1(level4_in[5551]),
   .I2(level4_in[5552]),
   .I3(level4_in[5553]),
   .I4(level4_in[5554]),
   .I5(level4_in[5555])
);

LUT6 #(
   .INIT(64'ha1d2ff2ca1d2ff2c)  
) LUT6_inst8702 (
   .O(to_level3[926]),
   .I0(level4_in[5556]),
   .I1(level4_in[5557]),
   .I2(level4_in[5558]),
   .I3(level4_in[5559]),
   .I4(level4_in[5560]),
   .I5(level4_in[5561])
);

LUT6 #(
   .INIT(64'hde331a37de331a37)  
) LUT6_inst8703 (
   .O(to_level3[927]),
   .I0(level4_in[5562]),
   .I1(level4_in[5563]),
   .I2(level4_in[5564]),
   .I3(level4_in[5565]),
   .I4(level4_in[5566]),
   .I5(level4_in[5567])
);

LUT6 #(
   .INIT(64'h048f7344048f7344)  
) LUT6_inst8704 (
   .O(to_level3[928]),
   .I0(level4_in[5568]),
   .I1(level4_in[5569]),
   .I2(level4_in[5570]),
   .I3(level4_in[5571]),
   .I4(level4_in[5572]),
   .I5(level4_in[5573])
);

LUT6 #(
   .INIT(64'ha2db169ba2db169b)  
) LUT6_inst8705 (
   .O(to_level3[929]),
   .I0(level4_in[5574]),
   .I1(level4_in[5575]),
   .I2(level4_in[5576]),
   .I3(level4_in[5577]),
   .I4(level4_in[5578]),
   .I5(level4_in[5579])
);

LUT6 #(
   .INIT(64'h6df8d3d26df8d3d2)  
) LUT6_inst8706 (
   .O(to_level3[930]),
   .I0(level4_in[5580]),
   .I1(level4_in[5581]),
   .I2(level4_in[5582]),
   .I3(level4_in[5583]),
   .I4(level4_in[5584]),
   .I5(level4_in[5585])
);

LUT6 #(
   .INIT(64'h2586324c2586324c)  
) LUT6_inst8707 (
   .O(to_level3[931]),
   .I0(level4_in[5586]),
   .I1(level4_in[5587]),
   .I2(level4_in[5588]),
   .I3(level4_in[5589]),
   .I4(level4_in[5590]),
   .I5(level4_in[5591])
);

LUT6 #(
   .INIT(64'h010116ff010116ff)  
) LUT6_inst8708 (
   .O(to_level3[932]),
   .I0(level4_in[5592]),
   .I1(level4_in[5593]),
   .I2(level4_in[5594]),
   .I3(level4_in[5595]),
   .I4(level4_in[5596]),
   .I5(level4_in[5597])
);

LUT6 #(
   .INIT(64'h3e9cb8533e9cb853)  
) LUT6_inst8709 (
   .O(to_level3[933]),
   .I0(level4_in[5598]),
   .I1(level4_in[5599]),
   .I2(level4_in[5600]),
   .I3(level4_in[5601]),
   .I4(level4_in[5602]),
   .I5(level4_in[5603])
);

LUT6 #(
   .INIT(64'hb2e2bbe4b2e2bbe4)  
) LUT6_inst8710 (
   .O(to_level3[934]),
   .I0(level4_in[5604]),
   .I1(level4_in[5605]),
   .I2(level4_in[5606]),
   .I3(level4_in[5607]),
   .I4(level4_in[5608]),
   .I5(level4_in[5609])
);

LUT6 #(
   .INIT(64'h53e04abe53e04abe)  
) LUT6_inst8711 (
   .O(to_level3[935]),
   .I0(level4_in[5610]),
   .I1(level4_in[5611]),
   .I2(level4_in[5612]),
   .I3(level4_in[5613]),
   .I4(level4_in[5614]),
   .I5(level4_in[5615])
);

LUT6 #(
   .INIT(64'h4a1fa4564a1fa456)  
) LUT6_inst8712 (
   .O(to_level3[936]),
   .I0(level4_in[5616]),
   .I1(level4_in[5617]),
   .I2(level4_in[5618]),
   .I3(level4_in[5619]),
   .I4(level4_in[5620]),
   .I5(level4_in[5621])
);

LUT6 #(
   .INIT(64'hdb835a2bdb835a2b)  
) LUT6_inst8713 (
   .O(to_level3[937]),
   .I0(level4_in[5622]),
   .I1(level4_in[5623]),
   .I2(level4_in[5624]),
   .I3(level4_in[5625]),
   .I4(level4_in[5626]),
   .I5(level4_in[5627])
);

LUT6 #(
   .INIT(64'h38d4c1a138d4c1a1)  
) LUT6_inst8714 (
   .O(to_level3[938]),
   .I0(level4_in[5628]),
   .I1(level4_in[5629]),
   .I2(level4_in[5630]),
   .I3(level4_in[5631]),
   .I4(level4_in[5632]),
   .I5(level4_in[5633])
);

LUT6 #(
   .INIT(64'h305413a4305413a4)  
) LUT6_inst8715 (
   .O(to_level3[939]),
   .I0(level4_in[5634]),
   .I1(level4_in[5635]),
   .I2(level4_in[5636]),
   .I3(level4_in[5637]),
   .I4(level4_in[5638]),
   .I5(level4_in[5639])
);

LUT6 #(
   .INIT(64'h55ddb7cd55ddb7cd)  
) LUT6_inst8716 (
   .O(to_level3[940]),
   .I0(level4_in[5640]),
   .I1(level4_in[5641]),
   .I2(level4_in[5642]),
   .I3(level4_in[5643]),
   .I4(level4_in[5644]),
   .I5(level4_in[5645])
);

LUT6 #(
   .INIT(64'hf3b79587f3b79587)  
) LUT6_inst8717 (
   .O(to_level3[941]),
   .I0(level4_in[5646]),
   .I1(level4_in[5647]),
   .I2(level4_in[5648]),
   .I3(level4_in[5649]),
   .I4(level4_in[5650]),
   .I5(level4_in[5651])
);

LUT6 #(
   .INIT(64'h8390ff808390ff80)  
) LUT6_inst8718 (
   .O(to_level3[942]),
   .I0(level4_in[5652]),
   .I1(level4_in[5653]),
   .I2(level4_in[5654]),
   .I3(level4_in[5655]),
   .I4(level4_in[5656]),
   .I5(level4_in[5657])
);

LUT6 #(
   .INIT(64'hea41fd6dea41fd6d)  
) LUT6_inst8719 (
   .O(to_level3[943]),
   .I0(level4_in[5658]),
   .I1(level4_in[5659]),
   .I2(level4_in[5660]),
   .I3(level4_in[5661]),
   .I4(level4_in[5662]),
   .I5(level4_in[5663])
);

LUT6 #(
   .INIT(64'h029b6a8e029b6a8e)  
) LUT6_inst8720 (
   .O(to_level3[944]),
   .I0(level4_in[5664]),
   .I1(level4_in[5665]),
   .I2(level4_in[5666]),
   .I3(level4_in[5667]),
   .I4(level4_in[5668]),
   .I5(level4_in[5669])
);

LUT6 #(
   .INIT(64'h38f0913d38f0913d)  
) LUT6_inst8721 (
   .O(to_level3[945]),
   .I0(level4_in[5670]),
   .I1(level4_in[5671]),
   .I2(level4_in[5672]),
   .I3(level4_in[5673]),
   .I4(level4_in[5674]),
   .I5(level4_in[5675])
);

LUT6 #(
   .INIT(64'h7e36cf9b7e36cf9b)  
) LUT6_inst8722 (
   .O(to_level3[946]),
   .I0(level4_in[5676]),
   .I1(level4_in[5677]),
   .I2(level4_in[5678]),
   .I3(level4_in[5679]),
   .I4(level4_in[5680]),
   .I5(level4_in[5681])
);

LUT6 #(
   .INIT(64'hb97408dab97408da)  
) LUT6_inst8723 (
   .O(to_level3[947]),
   .I0(level4_in[5682]),
   .I1(level4_in[5683]),
   .I2(level4_in[5684]),
   .I3(level4_in[5685]),
   .I4(level4_in[5686]),
   .I5(level4_in[5687])
);

LUT6 #(
   .INIT(64'h372697a4372697a4)  
) LUT6_inst8724 (
   .O(to_level3[948]),
   .I0(level4_in[5688]),
   .I1(level4_in[5689]),
   .I2(level4_in[5690]),
   .I3(level4_in[5691]),
   .I4(level4_in[5692]),
   .I5(level4_in[5693])
);

LUT6 #(
   .INIT(64'h983e47b9983e47b9)  
) LUT6_inst8725 (
   .O(to_level3[949]),
   .I0(level4_in[5694]),
   .I1(level4_in[5695]),
   .I2(level4_in[5696]),
   .I3(level4_in[5697]),
   .I4(level4_in[5698]),
   .I5(level4_in[5699])
);

LUT6 #(
   .INIT(64'h1d406f031d406f03)  
) LUT6_inst8726 (
   .O(to_level3[950]),
   .I0(level4_in[5700]),
   .I1(level4_in[5701]),
   .I2(level4_in[5702]),
   .I3(level4_in[5703]),
   .I4(level4_in[5704]),
   .I5(level4_in[5705])
);

LUT6 #(
   .INIT(64'hfd44f712fd44f712)  
) LUT6_inst8727 (
   .O(to_level3[951]),
   .I0(level4_in[5706]),
   .I1(level4_in[5707]),
   .I2(level4_in[5708]),
   .I3(level4_in[5709]),
   .I4(level4_in[5710]),
   .I5(level4_in[5711])
);

LUT6 #(
   .INIT(64'h06d7cb4106d7cb41)  
) LUT6_inst8728 (
   .O(to_level3[952]),
   .I0(level4_in[5712]),
   .I1(level4_in[5713]),
   .I2(level4_in[5714]),
   .I3(level4_in[5715]),
   .I4(level4_in[5716]),
   .I5(level4_in[5717])
);

LUT6 #(
   .INIT(64'hf5e0325df5e0325d)  
) LUT6_inst8729 (
   .O(to_level3[953]),
   .I0(level4_in[5718]),
   .I1(level4_in[5719]),
   .I2(level4_in[5720]),
   .I3(level4_in[5721]),
   .I4(level4_in[5722]),
   .I5(level4_in[5723])
);

LUT6 #(
   .INIT(64'h9da5a9ca9da5a9ca)  
) LUT6_inst8730 (
   .O(to_level3[954]),
   .I0(level4_in[5724]),
   .I1(level4_in[5725]),
   .I2(level4_in[5726]),
   .I3(level4_in[5727]),
   .I4(level4_in[5728]),
   .I5(level4_in[5729])
);

LUT6 #(
   .INIT(64'h6e462cde6e462cde)  
) LUT6_inst8731 (
   .O(to_level3[955]),
   .I0(level4_in[5730]),
   .I1(level4_in[5731]),
   .I2(level4_in[5732]),
   .I3(level4_in[5733]),
   .I4(level4_in[5734]),
   .I5(level4_in[5735])
);

LUT6 #(
   .INIT(64'ha734115ba734115b)  
) LUT6_inst8732 (
   .O(to_level3[956]),
   .I0(level4_in[5736]),
   .I1(level4_in[5737]),
   .I2(level4_in[5738]),
   .I3(level4_in[5739]),
   .I4(level4_in[5740]),
   .I5(level4_in[5741])
);

LUT6 #(
   .INIT(64'h7df19c6c7df19c6c)  
) LUT6_inst8733 (
   .O(to_level3[957]),
   .I0(level4_in[5742]),
   .I1(level4_in[5743]),
   .I2(level4_in[5744]),
   .I3(level4_in[5745]),
   .I4(level4_in[5746]),
   .I5(level4_in[5747])
);

LUT6 #(
   .INIT(64'h32ba0ac832ba0ac8)  
) LUT6_inst8734 (
   .O(to_level3[958]),
   .I0(level4_in[5748]),
   .I1(level4_in[5749]),
   .I2(level4_in[5750]),
   .I3(level4_in[5751]),
   .I4(level4_in[5752]),
   .I5(level4_in[5753])
);

LUT6 #(
   .INIT(64'h9d9c990e9d9c990e)  
) LUT6_inst8735 (
   .O(to_level3[959]),
   .I0(level4_in[5754]),
   .I1(level4_in[5755]),
   .I2(level4_in[5756]),
   .I3(level4_in[5757]),
   .I4(level4_in[5758]),
   .I5(level4_in[5759])
);

LUT6 #(
   .INIT(64'h8b4077cc8b4077cc)  
) LUT6_inst8736 (
   .O(to_level3[960]),
   .I0(level4_in[5760]),
   .I1(level4_in[5761]),
   .I2(level4_in[5762]),
   .I3(level4_in[5763]),
   .I4(level4_in[5764]),
   .I5(level4_in[5765])
);

LUT6 #(
   .INIT(64'h8699403286994032)  
) LUT6_inst8737 (
   .O(to_level3[961]),
   .I0(level4_in[5766]),
   .I1(level4_in[5767]),
   .I2(level4_in[5768]),
   .I3(level4_in[5769]),
   .I4(level4_in[5770]),
   .I5(level4_in[5771])
);

LUT6 #(
   .INIT(64'h7a2fafeb7a2fafeb)  
) LUT6_inst8738 (
   .O(to_level3[962]),
   .I0(level4_in[5772]),
   .I1(level4_in[5773]),
   .I2(level4_in[5774]),
   .I3(level4_in[5775]),
   .I4(level4_in[5776]),
   .I5(level4_in[5777])
);

LUT6 #(
   .INIT(64'h75a2012775a20127)  
) LUT6_inst8739 (
   .O(to_level3[963]),
   .I0(level4_in[5778]),
   .I1(level4_in[5779]),
   .I2(level4_in[5780]),
   .I3(level4_in[5781]),
   .I4(level4_in[5782]),
   .I5(level4_in[5783])
);

LUT6 #(
   .INIT(64'h3b994a333b994a33)  
) LUT6_inst8740 (
   .O(to_level3[964]),
   .I0(level4_in[5784]),
   .I1(level4_in[5785]),
   .I2(level4_in[5786]),
   .I3(level4_in[5787]),
   .I4(level4_in[5788]),
   .I5(level4_in[5789])
);

LUT6 #(
   .INIT(64'h7c7bc9da7c7bc9da)  
) LUT6_inst8741 (
   .O(to_level3[965]),
   .I0(level4_in[5790]),
   .I1(level4_in[5791]),
   .I2(level4_in[5792]),
   .I3(level4_in[5793]),
   .I4(level4_in[5794]),
   .I5(level4_in[5795])
);

LUT6 #(
   .INIT(64'hea2266d3ea2266d3)  
) LUT6_inst8742 (
   .O(to_level3[966]),
   .I0(level4_in[5796]),
   .I1(level4_in[5797]),
   .I2(level4_in[5798]),
   .I3(level4_in[5799]),
   .I4(level4_in[5800]),
   .I5(level4_in[5801])
);

LUT6 #(
   .INIT(64'h2753d8ff2753d8ff)  
) LUT6_inst8743 (
   .O(to_level3[967]),
   .I0(level4_in[5802]),
   .I1(level4_in[5803]),
   .I2(level4_in[5804]),
   .I3(level4_in[5805]),
   .I4(level4_in[5806]),
   .I5(level4_in[5807])
);

LUT6 #(
   .INIT(64'h6beab7746beab774)  
) LUT6_inst8744 (
   .O(to_level3[968]),
   .I0(level4_in[5808]),
   .I1(level4_in[5809]),
   .I2(level4_in[5810]),
   .I3(level4_in[5811]),
   .I4(level4_in[5812]),
   .I5(level4_in[5813])
);

LUT6 #(
   .INIT(64'h07a8325907a83259)  
) LUT6_inst8745 (
   .O(to_level3[969]),
   .I0(level4_in[5814]),
   .I1(level4_in[5815]),
   .I2(level4_in[5816]),
   .I3(level4_in[5817]),
   .I4(level4_in[5818]),
   .I5(level4_in[5819])
);

LUT6 #(
   .INIT(64'h624bac35624bac35)  
) LUT6_inst8746 (
   .O(to_level3[970]),
   .I0(level4_in[5820]),
   .I1(level4_in[5821]),
   .I2(level4_in[5822]),
   .I3(level4_in[5823]),
   .I4(level4_in[5824]),
   .I5(level4_in[5825])
);

LUT6 #(
   .INIT(64'hbde5e3d5bde5e3d5)  
) LUT6_inst8747 (
   .O(to_level3[971]),
   .I0(level4_in[5826]),
   .I1(level4_in[5827]),
   .I2(level4_in[5828]),
   .I3(level4_in[5829]),
   .I4(level4_in[5830]),
   .I5(level4_in[5831])
);

LUT6 #(
   .INIT(64'he37c7c06e37c7c06)  
) LUT6_inst8748 (
   .O(to_level3[972]),
   .I0(level4_in[5832]),
   .I1(level4_in[5833]),
   .I2(level4_in[5834]),
   .I3(level4_in[5835]),
   .I4(level4_in[5836]),
   .I5(level4_in[5837])
);

LUT6 #(
   .INIT(64'he4ac8995e4ac8995)  
) LUT6_inst8749 (
   .O(to_level3[973]),
   .I0(level4_in[5838]),
   .I1(level4_in[5839]),
   .I2(level4_in[5840]),
   .I3(level4_in[5841]),
   .I4(level4_in[5842]),
   .I5(level4_in[5843])
);

LUT6 #(
   .INIT(64'he7618f9de7618f9d)  
) LUT6_inst8750 (
   .O(to_level3[974]),
   .I0(level4_in[5844]),
   .I1(level4_in[5845]),
   .I2(level4_in[5846]),
   .I3(level4_in[5847]),
   .I4(level4_in[5848]),
   .I5(level4_in[5849])
);

LUT6 #(
   .INIT(64'h9a0de4299a0de429)  
) LUT6_inst8751 (
   .O(to_level3[975]),
   .I0(level4_in[5850]),
   .I1(level4_in[5851]),
   .I2(level4_in[5852]),
   .I3(level4_in[5853]),
   .I4(level4_in[5854]),
   .I5(level4_in[5855])
);

LUT6 #(
   .INIT(64'hc8f21976c8f21976)  
) LUT6_inst8752 (
   .O(to_level3[976]),
   .I0(level4_in[5856]),
   .I1(level4_in[5857]),
   .I2(level4_in[5858]),
   .I3(level4_in[5859]),
   .I4(level4_in[5860]),
   .I5(level4_in[5861])
);

LUT6 #(
   .INIT(64'h1c621a891c621a89)  
) LUT6_inst8753 (
   .O(to_level3[977]),
   .I0(level4_in[5862]),
   .I1(level4_in[5863]),
   .I2(level4_in[5864]),
   .I3(level4_in[5865]),
   .I4(level4_in[5866]),
   .I5(level4_in[5867])
);

LUT6 #(
   .INIT(64'h7af7d0587af7d058)  
) LUT6_inst8754 (
   .O(to_level3[978]),
   .I0(level4_in[5868]),
   .I1(level4_in[5869]),
   .I2(level4_in[5870]),
   .I3(level4_in[5871]),
   .I4(level4_in[5872]),
   .I5(level4_in[5873])
);

LUT6 #(
   .INIT(64'h3bd932413bd93241)  
) LUT6_inst8755 (
   .O(to_level3[979]),
   .I0(level4_in[5874]),
   .I1(level4_in[5875]),
   .I2(level4_in[5876]),
   .I3(level4_in[5877]),
   .I4(level4_in[5878]),
   .I5(level4_in[5879])
);

LUT6 #(
   .INIT(64'h367eac14367eac14)  
) LUT6_inst8756 (
   .O(to_level3[980]),
   .I0(level4_in[5880]),
   .I1(level4_in[5881]),
   .I2(level4_in[5882]),
   .I3(level4_in[5883]),
   .I4(level4_in[5884]),
   .I5(level4_in[5885])
);

LUT6 #(
   .INIT(64'h9d1e12d69d1e12d6)  
) LUT6_inst8757 (
   .O(to_level3[981]),
   .I0(level4_in[5886]),
   .I1(level4_in[5887]),
   .I2(level4_in[5888]),
   .I3(level4_in[5889]),
   .I4(level4_in[5890]),
   .I5(level4_in[5891])
);

LUT6 #(
   .INIT(64'h43cbfdea43cbfdea)  
) LUT6_inst8758 (
   .O(to_level3[982]),
   .I0(level4_in[5892]),
   .I1(level4_in[5893]),
   .I2(level4_in[5894]),
   .I3(level4_in[5895]),
   .I4(level4_in[5896]),
   .I5(level4_in[5897])
);

LUT6 #(
   .INIT(64'h53c6c35653c6c356)  
) LUT6_inst8759 (
   .O(to_level3[983]),
   .I0(level4_in[5898]),
   .I1(level4_in[5899]),
   .I2(level4_in[5900]),
   .I3(level4_in[5901]),
   .I4(level4_in[5902]),
   .I5(level4_in[5903])
);

LUT6 #(
   .INIT(64'h807dd556807dd556)  
) LUT6_inst8760 (
   .O(to_level3[984]),
   .I0(level4_in[5904]),
   .I1(level4_in[5905]),
   .I2(level4_in[5906]),
   .I3(level4_in[5907]),
   .I4(level4_in[5908]),
   .I5(level4_in[5909])
);

LUT6 #(
   .INIT(64'hb1854f20b1854f20)  
) LUT6_inst8761 (
   .O(to_level3[985]),
   .I0(level4_in[5910]),
   .I1(level4_in[5911]),
   .I2(level4_in[5912]),
   .I3(level4_in[5913]),
   .I4(level4_in[5914]),
   .I5(level4_in[5915])
);

LUT6 #(
   .INIT(64'he0e9168ae0e9168a)  
) LUT6_inst8762 (
   .O(to_level3[986]),
   .I0(level4_in[5916]),
   .I1(level4_in[5917]),
   .I2(level4_in[5918]),
   .I3(level4_in[5919]),
   .I4(level4_in[5920]),
   .I5(level4_in[5921])
);

LUT6 #(
   .INIT(64'hcedc3c89cedc3c89)  
) LUT6_inst8763 (
   .O(to_level3[987]),
   .I0(level4_in[5922]),
   .I1(level4_in[5923]),
   .I2(level4_in[5924]),
   .I3(level4_in[5925]),
   .I4(level4_in[5926]),
   .I5(level4_in[5927])
);

LUT6 #(
   .INIT(64'h33d8254633d82546)  
) LUT6_inst8764 (
   .O(to_level3[988]),
   .I0(level4_in[5928]),
   .I1(level4_in[5929]),
   .I2(level4_in[5930]),
   .I3(level4_in[5931]),
   .I4(level4_in[5932]),
   .I5(level4_in[5933])
);

LUT6 #(
   .INIT(64'hd8b3202fd8b3202f)  
) LUT6_inst8765 (
   .O(to_level3[989]),
   .I0(level4_in[5934]),
   .I1(level4_in[5935]),
   .I2(level4_in[5936]),
   .I3(level4_in[5937]),
   .I4(level4_in[5938]),
   .I5(level4_in[5939])
);

LUT6 #(
   .INIT(64'hbdfadc45bdfadc45)  
) LUT6_inst8766 (
   .O(to_level3[990]),
   .I0(level4_in[5940]),
   .I1(level4_in[5941]),
   .I2(level4_in[5942]),
   .I3(level4_in[5943]),
   .I4(level4_in[5944]),
   .I5(level4_in[5945])
);

LUT6 #(
   .INIT(64'h7241c3dc7241c3dc)  
) LUT6_inst8767 (
   .O(to_level3[991]),
   .I0(level4_in[5946]),
   .I1(level4_in[5947]),
   .I2(level4_in[5948]),
   .I3(level4_in[5949]),
   .I4(level4_in[5950]),
   .I5(level4_in[5951])
);

LUT6 #(
   .INIT(64'he4d5ac23e4d5ac23)  
) LUT6_inst8768 (
   .O(to_level3[992]),
   .I0(level4_in[5952]),
   .I1(level4_in[5953]),
   .I2(level4_in[5954]),
   .I3(level4_in[5955]),
   .I4(level4_in[5956]),
   .I5(level4_in[5957])
);

LUT6 #(
   .INIT(64'h8b36d3238b36d323)  
) LUT6_inst8769 (
   .O(to_level3[993]),
   .I0(level4_in[5958]),
   .I1(level4_in[5959]),
   .I2(level4_in[5960]),
   .I3(level4_in[5961]),
   .I4(level4_in[5962]),
   .I5(level4_in[5963])
);

LUT6 #(
   .INIT(64'h9901af6b9901af6b)  
) LUT6_inst8770 (
   .O(to_level3[994]),
   .I0(level4_in[5964]),
   .I1(level4_in[5965]),
   .I2(level4_in[5966]),
   .I3(level4_in[5967]),
   .I4(level4_in[5968]),
   .I5(level4_in[5969])
);

LUT6 #(
   .INIT(64'h8bc661278bc66127)  
) LUT6_inst8771 (
   .O(to_level3[995]),
   .I0(level4_in[5970]),
   .I1(level4_in[5971]),
   .I2(level4_in[5972]),
   .I3(level4_in[5973]),
   .I4(level4_in[5974]),
   .I5(level4_in[5975])
);

LUT6 #(
   .INIT(64'h61290bde61290bde)  
) LUT6_inst8772 (
   .O(to_level3[996]),
   .I0(level4_in[5976]),
   .I1(level4_in[5977]),
   .I2(level4_in[5978]),
   .I3(level4_in[5979]),
   .I4(level4_in[5980]),
   .I5(level4_in[5981])
);

LUT6 #(
   .INIT(64'h8cf408ab8cf408ab)  
) LUT6_inst8773 (
   .O(to_level3[997]),
   .I0(level4_in[5982]),
   .I1(level4_in[5983]),
   .I2(level4_in[5984]),
   .I3(level4_in[5985]),
   .I4(level4_in[5986]),
   .I5(level4_in[5987])
);

LUT6 #(
   .INIT(64'h6f5f91b06f5f91b0)  
) LUT6_inst8774 (
   .O(to_level3[998]),
   .I0(level4_in[5988]),
   .I1(level4_in[5989]),
   .I2(level4_in[5990]),
   .I3(level4_in[5991]),
   .I4(level4_in[5992]),
   .I5(level4_in[5993])
);

LUT6 #(
   .INIT(64'h5189cc565189cc56)  
) LUT6_inst8775 (
   .O(to_level3[999]),
   .I0(level4_in[5994]),
   .I1(level4_in[5995]),
   .I2(level4_in[5996]),
   .I3(level4_in[5997]),
   .I4(level4_in[5998]),
   .I5(level4_in[5999])
);

LUT6 #(
   .INIT(64'ha0f1a570a0f1a570)  
) LUT6_inst8776 (
   .O(to_level3[1000]),
   .I0(level4_in[6000]),
   .I1(level4_in[6001]),
   .I2(level4_in[6002]),
   .I3(level4_in[6003]),
   .I4(level4_in[6004]),
   .I5(level4_in[6005])
);

LUT6 #(
   .INIT(64'ha6323fd0a6323fd0)  
) LUT6_inst8777 (
   .O(to_level3[1001]),
   .I0(level4_in[6006]),
   .I1(level4_in[6007]),
   .I2(level4_in[6008]),
   .I3(level4_in[6009]),
   .I4(level4_in[6010]),
   .I5(level4_in[6011])
);

LUT6 #(
   .INIT(64'h11d3552011d35520)  
) LUT6_inst8778 (
   .O(to_level3[1002]),
   .I0(level4_in[6012]),
   .I1(level4_in[6013]),
   .I2(level4_in[6014]),
   .I3(level4_in[6015]),
   .I4(level4_in[6016]),
   .I5(level4_in[6017])
);

LUT6 #(
   .INIT(64'h42f60d1a42f60d1a)  
) LUT6_inst8779 (
   .O(to_level3[1003]),
   .I0(level4_in[6018]),
   .I1(level4_in[6019]),
   .I2(level4_in[6020]),
   .I3(level4_in[6021]),
   .I4(level4_in[6022]),
   .I5(level4_in[6023])
);

LUT6 #(
   .INIT(64'hbfaa9aa4bfaa9aa4)  
) LUT6_inst8780 (
   .O(to_level3[1004]),
   .I0(level4_in[6024]),
   .I1(level4_in[6025]),
   .I2(level4_in[6026]),
   .I3(level4_in[6027]),
   .I4(level4_in[6028]),
   .I5(level4_in[6029])
);

LUT6 #(
   .INIT(64'hfac2770bfac2770b)  
) LUT6_inst8781 (
   .O(to_level3[1005]),
   .I0(level4_in[6030]),
   .I1(level4_in[6031]),
   .I2(level4_in[6032]),
   .I3(level4_in[6033]),
   .I4(level4_in[6034]),
   .I5(level4_in[6035])
);

LUT6 #(
   .INIT(64'hdba65c87dba65c87)  
) LUT6_inst8782 (
   .O(to_level3[1006]),
   .I0(level4_in[6036]),
   .I1(level4_in[6037]),
   .I2(level4_in[6038]),
   .I3(level4_in[6039]),
   .I4(level4_in[6040]),
   .I5(level4_in[6041])
);

LUT6 #(
   .INIT(64'he4131c18e4131c18)  
) LUT6_inst8783 (
   .O(to_level3[1007]),
   .I0(level4_in[6042]),
   .I1(level4_in[6043]),
   .I2(level4_in[6044]),
   .I3(level4_in[6045]),
   .I4(level4_in[6046]),
   .I5(level4_in[6047])
);

LUT6 #(
   .INIT(64'hf63c9e5af63c9e5a)  
) LUT6_inst8784 (
   .O(to_level3[1008]),
   .I0(level4_in[6048]),
   .I1(level4_in[6049]),
   .I2(level4_in[6050]),
   .I3(level4_in[6051]),
   .I4(level4_in[6052]),
   .I5(level4_in[6053])
);

LUT6 #(
   .INIT(64'ha5c0722da5c0722d)  
) LUT6_inst8785 (
   .O(to_level3[1009]),
   .I0(level4_in[6054]),
   .I1(level4_in[6055]),
   .I2(level4_in[6056]),
   .I3(level4_in[6057]),
   .I4(level4_in[6058]),
   .I5(level4_in[6059])
);

LUT6 #(
   .INIT(64'h2e7f89892e7f8989)  
) LUT6_inst8786 (
   .O(to_level3[1010]),
   .I0(level4_in[6060]),
   .I1(level4_in[6061]),
   .I2(level4_in[6062]),
   .I3(level4_in[6063]),
   .I4(level4_in[6064]),
   .I5(level4_in[6065])
);

LUT6 #(
   .INIT(64'h184382da184382da)  
) LUT6_inst8787 (
   .O(to_level3[1011]),
   .I0(level4_in[6066]),
   .I1(level4_in[6067]),
   .I2(level4_in[6068]),
   .I3(level4_in[6069]),
   .I4(level4_in[6070]),
   .I5(level4_in[6071])
);

LUT6 #(
   .INIT(64'hd5ecd508d5ecd508)  
) LUT6_inst8788 (
   .O(to_level3[1012]),
   .I0(level4_in[6072]),
   .I1(level4_in[6073]),
   .I2(level4_in[6074]),
   .I3(level4_in[6075]),
   .I4(level4_in[6076]),
   .I5(level4_in[6077])
);

LUT6 #(
   .INIT(64'hfab6a159fab6a159)  
) LUT6_inst8789 (
   .O(to_level3[1013]),
   .I0(level4_in[6078]),
   .I1(level4_in[6079]),
   .I2(level4_in[6080]),
   .I3(level4_in[6081]),
   .I4(level4_in[6082]),
   .I5(level4_in[6083])
);

LUT6 #(
   .INIT(64'h593191cd593191cd)  
) LUT6_inst8790 (
   .O(to_level3[1014]),
   .I0(level4_in[6084]),
   .I1(level4_in[6085]),
   .I2(level4_in[6086]),
   .I3(level4_in[6087]),
   .I4(level4_in[6088]),
   .I5(level4_in[6089])
);

LUT6 #(
   .INIT(64'hb52899deb52899de)  
) LUT6_inst8791 (
   .O(to_level3[1015]),
   .I0(level4_in[6090]),
   .I1(level4_in[6091]),
   .I2(level4_in[6092]),
   .I3(level4_in[6093]),
   .I4(level4_in[6094]),
   .I5(level4_in[6095])
);

LUT6 #(
   .INIT(64'hc38b8157c38b8157)  
) LUT6_inst8792 (
   .O(to_level3[1016]),
   .I0(level4_in[6096]),
   .I1(level4_in[6097]),
   .I2(level4_in[6098]),
   .I3(level4_in[6099]),
   .I4(level4_in[6100]),
   .I5(level4_in[6101])
);

LUT6 #(
   .INIT(64'h869c0579869c0579)  
) LUT6_inst8793 (
   .O(to_level3[1017]),
   .I0(level4_in[6102]),
   .I1(level4_in[6103]),
   .I2(level4_in[6104]),
   .I3(level4_in[6105]),
   .I4(level4_in[6106]),
   .I5(level4_in[6107])
);

LUT6 #(
   .INIT(64'h2e6ce6bd2e6ce6bd)  
) LUT6_inst8794 (
   .O(to_level3[1018]),
   .I0(level4_in[6108]),
   .I1(level4_in[6109]),
   .I2(level4_in[6110]),
   .I3(level4_in[6111]),
   .I4(level4_in[6112]),
   .I5(level4_in[6113])
);

LUT6 #(
   .INIT(64'hcb0e2b66cb0e2b66)  
) LUT6_inst8795 (
   .O(to_level3[1019]),
   .I0(level4_in[6114]),
   .I1(level4_in[6115]),
   .I2(level4_in[6116]),
   .I3(level4_in[6117]),
   .I4(level4_in[6118]),
   .I5(level4_in[6119])
);

LUT6 #(
   .INIT(64'h911727b5911727b5)  
) LUT6_inst8796 (
   .O(to_level3[1020]),
   .I0(level4_in[6120]),
   .I1(level4_in[6121]),
   .I2(level4_in[6122]),
   .I3(level4_in[6123]),
   .I4(level4_in[6124]),
   .I5(level4_in[6125])
);

LUT6 #(
   .INIT(64'hecb34248ecb34248)  
) LUT6_inst8797 (
   .O(to_level3[1021]),
   .I0(level4_in[6126]),
   .I1(level4_in[6127]),
   .I2(level4_in[6128]),
   .I3(level4_in[6129]),
   .I4(level4_in[6130]),
   .I5(level4_in[6131])
);

LUT6 #(
   .INIT(64'h6bcb7ecc6bcb7ecc)  
) LUT6_inst8798 (
   .O(to_level3[1022]),
   .I0(level4_in[6132]),
   .I1(level4_in[6133]),
   .I2(level4_in[6134]),
   .I3(level4_in[6135]),
   .I4(level4_in[6136]),
   .I5(level4_in[6137])
);

LUT6 #(
   .INIT(64'h945db2db945db2db)  
) LUT6_inst8799 (
   .O(to_level3[1023]),
   .I0(level4_in[6138]),
   .I1(level4_in[6139]),
   .I2(level4_in[6140]),
   .I3(level4_in[6141]),
   .I4(level4_in[6142]),
   .I5(level4_in[6143])
);

LUT6 #(
   .INIT(64'h394a2d83394a2d83)  
) LUT6_inst8800 (
   .O(to_level3[1024]),
   .I0(level4_in[6144]),
   .I1(level4_in[6145]),
   .I2(level4_in[6146]),
   .I3(level4_in[6147]),
   .I4(level4_in[6148]),
   .I5(level4_in[6149])
);

LUT6 #(
   .INIT(64'hebebda88ebebda88)  
) LUT6_inst8801 (
   .O(to_level3[1025]),
   .I0(level4_in[6150]),
   .I1(level4_in[6151]),
   .I2(level4_in[6152]),
   .I3(level4_in[6153]),
   .I4(level4_in[6154]),
   .I5(level4_in[6155])
);

LUT6 #(
   .INIT(64'h14a7dd5c14a7dd5c)  
) LUT6_inst8802 (
   .O(to_level3[1026]),
   .I0(level4_in[6156]),
   .I1(level4_in[6157]),
   .I2(level4_in[6158]),
   .I3(level4_in[6159]),
   .I4(level4_in[6160]),
   .I5(level4_in[6161])
);

LUT6 #(
   .INIT(64'h821d7b58821d7b58)  
) LUT6_inst8803 (
   .O(to_level3[1027]),
   .I0(level4_in[6162]),
   .I1(level4_in[6163]),
   .I2(level4_in[6164]),
   .I3(level4_in[6165]),
   .I4(level4_in[6166]),
   .I5(level4_in[6167])
);

LUT6 #(
   .INIT(64'habfb760aabfb760a)  
) LUT6_inst8804 (
   .O(to_level3[1028]),
   .I0(level4_in[6168]),
   .I1(level4_in[6169]),
   .I2(level4_in[6170]),
   .I3(level4_in[6171]),
   .I4(level4_in[6172]),
   .I5(level4_in[6173])
);

LUT6 #(
   .INIT(64'h8931b1e08931b1e0)  
) LUT6_inst8805 (
   .O(to_level3[1029]),
   .I0(level4_in[6174]),
   .I1(level4_in[6175]),
   .I2(level4_in[6176]),
   .I3(level4_in[6177]),
   .I4(level4_in[6178]),
   .I5(level4_in[6179])
);

LUT6 #(
   .INIT(64'h4995789749957897)  
) LUT6_inst8806 (
   .O(to_level3[1030]),
   .I0(level4_in[6180]),
   .I1(level4_in[6181]),
   .I2(level4_in[6182]),
   .I3(level4_in[6183]),
   .I4(level4_in[6184]),
   .I5(level4_in[6185])
);

LUT6 #(
   .INIT(64'h1d9e3fec1d9e3fec)  
) LUT6_inst8807 (
   .O(to_level3[1031]),
   .I0(level4_in[6186]),
   .I1(level4_in[6187]),
   .I2(level4_in[6188]),
   .I3(level4_in[6189]),
   .I4(level4_in[6190]),
   .I5(level4_in[6191])
);

LUT6 #(
   .INIT(64'h137db874137db874)  
) LUT6_inst8808 (
   .O(to_level3[1032]),
   .I0(level4_in[6192]),
   .I1(level4_in[6193]),
   .I2(level4_in[6194]),
   .I3(level4_in[6195]),
   .I4(level4_in[6196]),
   .I5(level4_in[6197])
);

LUT6 #(
   .INIT(64'he25c79eae25c79ea)  
) LUT6_inst8809 (
   .O(to_level3[1033]),
   .I0(level4_in[6198]),
   .I1(level4_in[6199]),
   .I2(level4_in[6200]),
   .I3(level4_in[6201]),
   .I4(level4_in[6202]),
   .I5(level4_in[6203])
);

LUT6 #(
   .INIT(64'h4fc627aa4fc627aa)  
) LUT6_inst8810 (
   .O(to_level3[1034]),
   .I0(level4_in[6204]),
   .I1(level4_in[6205]),
   .I2(level4_in[6206]),
   .I3(level4_in[6207]),
   .I4(level4_in[6208]),
   .I5(level4_in[6209])
);

LUT6 #(
   .INIT(64'hfacf8c9efacf8c9e)  
) LUT6_inst8811 (
   .O(to_level3[1035]),
   .I0(level4_in[6210]),
   .I1(level4_in[6211]),
   .I2(level4_in[6212]),
   .I3(level4_in[6213]),
   .I4(level4_in[6214]),
   .I5(level4_in[6215])
);

LUT6 #(
   .INIT(64'hf2813be1f2813be1)  
) LUT6_inst8812 (
   .O(to_level3[1036]),
   .I0(level4_in[6216]),
   .I1(level4_in[6217]),
   .I2(level4_in[6218]),
   .I3(level4_in[6219]),
   .I4(level4_in[6220]),
   .I5(level4_in[6221])
);

LUT6 #(
   .INIT(64'h4f3288e44f3288e4)  
) LUT6_inst8813 (
   .O(to_level3[1037]),
   .I0(level4_in[6222]),
   .I1(level4_in[6223]),
   .I2(level4_in[6224]),
   .I3(level4_in[6225]),
   .I4(level4_in[6226]),
   .I5(level4_in[6227])
);

LUT6 #(
   .INIT(64'h868a9e99868a9e99)  
) LUT6_inst8814 (
   .O(to_level3[1038]),
   .I0(level4_in[6228]),
   .I1(level4_in[6229]),
   .I2(level4_in[6230]),
   .I3(level4_in[6231]),
   .I4(level4_in[6232]),
   .I5(level4_in[6233])
);

LUT6 #(
   .INIT(64'h12ad9d3512ad9d35)  
) LUT6_inst8815 (
   .O(to_level3[1039]),
   .I0(level4_in[6234]),
   .I1(level4_in[6235]),
   .I2(level4_in[6236]),
   .I3(level4_in[6237]),
   .I4(level4_in[6238]),
   .I5(level4_in[6239])
);

LUT6 #(
   .INIT(64'hb562e446b562e446)  
) LUT6_inst8816 (
   .O(to_level3[1040]),
   .I0(level4_in[6240]),
   .I1(level4_in[6241]),
   .I2(level4_in[6242]),
   .I3(level4_in[6243]),
   .I4(level4_in[6244]),
   .I5(level4_in[6245])
);

LUT6 #(
   .INIT(64'h1f43e2531f43e253)  
) LUT6_inst8817 (
   .O(to_level3[1041]),
   .I0(level4_in[6246]),
   .I1(level4_in[6247]),
   .I2(level4_in[6248]),
   .I3(level4_in[6249]),
   .I4(level4_in[6250]),
   .I5(level4_in[6251])
);

LUT6 #(
   .INIT(64'ha4ca0659a4ca0659)  
) LUT6_inst8818 (
   .O(to_level3[1042]),
   .I0(level4_in[6252]),
   .I1(level4_in[6253]),
   .I2(level4_in[6254]),
   .I3(level4_in[6255]),
   .I4(level4_in[6256]),
   .I5(level4_in[6257])
);

LUT6 #(
   .INIT(64'h6aed11a06aed11a0)  
) LUT6_inst8819 (
   .O(to_level3[1043]),
   .I0(level4_in[6258]),
   .I1(level4_in[6259]),
   .I2(level4_in[6260]),
   .I3(level4_in[6261]),
   .I4(level4_in[6262]),
   .I5(level4_in[6263])
);

LUT6 #(
   .INIT(64'h0e895b8b0e895b8b)  
) LUT6_inst8820 (
   .O(to_level3[1044]),
   .I0(level4_in[6264]),
   .I1(level4_in[6265]),
   .I2(level4_in[6266]),
   .I3(level4_in[6267]),
   .I4(level4_in[6268]),
   .I5(level4_in[6269])
);

LUT6 #(
   .INIT(64'he93f1d6ee93f1d6e)  
) LUT6_inst8821 (
   .O(to_level3[1045]),
   .I0(level4_in[6270]),
   .I1(level4_in[6271]),
   .I2(level4_in[6272]),
   .I3(level4_in[6273]),
   .I4(level4_in[6274]),
   .I5(level4_in[6275])
);

LUT6 #(
   .INIT(64'h5acd75b55acd75b5)  
) LUT6_inst8822 (
   .O(to_level3[1046]),
   .I0(level4_in[6276]),
   .I1(level4_in[6277]),
   .I2(level4_in[6278]),
   .I3(level4_in[6279]),
   .I4(level4_in[6280]),
   .I5(level4_in[6281])
);

LUT6 #(
   .INIT(64'h1d8583911d858391)  
) LUT6_inst8823 (
   .O(to_level3[1047]),
   .I0(level4_in[6282]),
   .I1(level4_in[6283]),
   .I2(level4_in[6284]),
   .I3(level4_in[6285]),
   .I4(level4_in[6286]),
   .I5(level4_in[6287])
);

LUT6 #(
   .INIT(64'hc90cc86dc90cc86d)  
) LUT6_inst8824 (
   .O(to_level3[1048]),
   .I0(level4_in[6288]),
   .I1(level4_in[6289]),
   .I2(level4_in[6290]),
   .I3(level4_in[6291]),
   .I4(level4_in[6292]),
   .I5(level4_in[6293])
);

LUT6 #(
   .INIT(64'h7d4f8f427d4f8f42)  
) LUT6_inst8825 (
   .O(to_level3[1049]),
   .I0(level4_in[6294]),
   .I1(level4_in[6295]),
   .I2(level4_in[6296]),
   .I3(level4_in[6297]),
   .I4(level4_in[6298]),
   .I5(level4_in[6299])
);

LUT6 #(
   .INIT(64'h9f36648e9f36648e)  
) LUT6_inst8826 (
   .O(to_level3[1050]),
   .I0(level4_in[6300]),
   .I1(level4_in[6301]),
   .I2(level4_in[6302]),
   .I3(level4_in[6303]),
   .I4(level4_in[6304]),
   .I5(level4_in[6305])
);

LUT6 #(
   .INIT(64'h80e6149f80e6149f)  
) LUT6_inst8827 (
   .O(to_level3[1051]),
   .I0(level4_in[6306]),
   .I1(level4_in[6307]),
   .I2(level4_in[6308]),
   .I3(level4_in[6309]),
   .I4(level4_in[6310]),
   .I5(level4_in[6311])
);

LUT6 #(
   .INIT(64'hfc2c32b0fc2c32b0)  
) LUT6_inst8828 (
   .O(to_level3[1052]),
   .I0(level4_in[6312]),
   .I1(level4_in[6313]),
   .I2(level4_in[6314]),
   .I3(level4_in[6315]),
   .I4(level4_in[6316]),
   .I5(level4_in[6317])
);

LUT6 #(
   .INIT(64'hb52a2dffb52a2dff)  
) LUT6_inst8829 (
   .O(to_level3[1053]),
   .I0(level4_in[6318]),
   .I1(level4_in[6319]),
   .I2(level4_in[6320]),
   .I3(level4_in[6321]),
   .I4(level4_in[6322]),
   .I5(level4_in[6323])
);

LUT6 #(
   .INIT(64'h56371b6656371b66)  
) LUT6_inst8830 (
   .O(to_level3[1054]),
   .I0(level4_in[6324]),
   .I1(level4_in[6325]),
   .I2(level4_in[6326]),
   .I3(level4_in[6327]),
   .I4(level4_in[6328]),
   .I5(level4_in[6329])
);

LUT6 #(
   .INIT(64'h10eb813510eb8135)  
) LUT6_inst8831 (
   .O(to_level3[1055]),
   .I0(level4_in[6330]),
   .I1(level4_in[6331]),
   .I2(level4_in[6332]),
   .I3(level4_in[6333]),
   .I4(level4_in[6334]),
   .I5(level4_in[6335])
);

LUT6 #(
   .INIT(64'ha3b81208a3b81208)  
) LUT6_inst8832 (
   .O(to_level3[1056]),
   .I0(level4_in[6336]),
   .I1(level4_in[6337]),
   .I2(level4_in[6338]),
   .I3(level4_in[6339]),
   .I4(level4_in[6340]),
   .I5(level4_in[6341])
);

LUT6 #(
   .INIT(64'hb1b47f8cb1b47f8c)  
) LUT6_inst8833 (
   .O(to_level3[1057]),
   .I0(level4_in[6342]),
   .I1(level4_in[6343]),
   .I2(level4_in[6344]),
   .I3(level4_in[6345]),
   .I4(level4_in[6346]),
   .I5(level4_in[6347])
);

LUT6 #(
   .INIT(64'hf62b72f8f62b72f8)  
) LUT6_inst8834 (
   .O(to_level3[1058]),
   .I0(level4_in[6348]),
   .I1(level4_in[6349]),
   .I2(level4_in[6350]),
   .I3(level4_in[6351]),
   .I4(level4_in[6352]),
   .I5(level4_in[6353])
);

LUT6 #(
   .INIT(64'h72a049d372a049d3)  
) LUT6_inst8835 (
   .O(to_level3[1059]),
   .I0(level4_in[6354]),
   .I1(level4_in[6355]),
   .I2(level4_in[6356]),
   .I3(level4_in[6357]),
   .I4(level4_in[6358]),
   .I5(level4_in[6359])
);

LUT6 #(
   .INIT(64'h25fac3e125fac3e1)  
) LUT6_inst8836 (
   .O(to_level3[1060]),
   .I0(level4_in[6360]),
   .I1(level4_in[6361]),
   .I2(level4_in[6362]),
   .I3(level4_in[6363]),
   .I4(level4_in[6364]),
   .I5(level4_in[6365])
);

LUT6 #(
   .INIT(64'hac7cccc2ac7cccc2)  
) LUT6_inst8837 (
   .O(to_level3[1061]),
   .I0(level4_in[6366]),
   .I1(level4_in[6367]),
   .I2(level4_in[6368]),
   .I3(level4_in[6369]),
   .I4(level4_in[6370]),
   .I5(level4_in[6371])
);

LUT6 #(
   .INIT(64'hb30c04afb30c04af)  
) LUT6_inst8838 (
   .O(to_level3[1062]),
   .I0(level4_in[6372]),
   .I1(level4_in[6373]),
   .I2(level4_in[6374]),
   .I3(level4_in[6375]),
   .I4(level4_in[6376]),
   .I5(level4_in[6377])
);

LUT6 #(
   .INIT(64'h74ca6cdc74ca6cdc)  
) LUT6_inst8839 (
   .O(to_level3[1063]),
   .I0(level4_in[6378]),
   .I1(level4_in[6379]),
   .I2(level4_in[6380]),
   .I3(level4_in[6381]),
   .I4(level4_in[6382]),
   .I5(level4_in[6383])
);

LUT6 #(
   .INIT(64'hff790caaff790caa)  
) LUT6_inst8840 (
   .O(to_level3[1064]),
   .I0(level4_in[6384]),
   .I1(level4_in[6385]),
   .I2(level4_in[6386]),
   .I3(level4_in[6387]),
   .I4(level4_in[6388]),
   .I5(level4_in[6389])
);

LUT6 #(
   .INIT(64'hd72f1b80d72f1b80)  
) LUT6_inst8841 (
   .O(to_level3[1065]),
   .I0(level4_in[6390]),
   .I1(level4_in[6391]),
   .I2(level4_in[6392]),
   .I3(level4_in[6393]),
   .I4(level4_in[6394]),
   .I5(level4_in[6395])
);

LUT6 #(
   .INIT(64'h271f1bde271f1bde)  
) LUT6_inst8842 (
   .O(to_level3[1066]),
   .I0(level4_in[6396]),
   .I1(level4_in[6397]),
   .I2(level4_in[6398]),
   .I3(level4_in[6399]),
   .I4(level4_in[6400]),
   .I5(level4_in[6401])
);

LUT6 #(
   .INIT(64'hfe5cb97afe5cb97a)  
) LUT6_inst8843 (
   .O(to_level3[1067]),
   .I0(level4_in[6402]),
   .I1(level4_in[6403]),
   .I2(level4_in[6404]),
   .I3(level4_in[6405]),
   .I4(level4_in[6406]),
   .I5(level4_in[6407])
);

LUT6 #(
   .INIT(64'hb73b79c8b73b79c8)  
) LUT6_inst8844 (
   .O(to_level3[1068]),
   .I0(level4_in[6408]),
   .I1(level4_in[6409]),
   .I2(level4_in[6410]),
   .I3(level4_in[6411]),
   .I4(level4_in[6412]),
   .I5(level4_in[6413])
);

LUT6 #(
   .INIT(64'hee26e679ee26e679)  
) LUT6_inst8845 (
   .O(to_level3[1069]),
   .I0(level4_in[6414]),
   .I1(level4_in[6415]),
   .I2(level4_in[6416]),
   .I3(level4_in[6417]),
   .I4(level4_in[6418]),
   .I5(level4_in[6419])
);

LUT6 #(
   .INIT(64'h030660db030660db)  
) LUT6_inst8846 (
   .O(to_level3[1070]),
   .I0(level4_in[6420]),
   .I1(level4_in[6421]),
   .I2(level4_in[6422]),
   .I3(level4_in[6423]),
   .I4(level4_in[6424]),
   .I5(level4_in[6425])
);

LUT6 #(
   .INIT(64'h2ec583ca2ec583ca)  
) LUT6_inst8847 (
   .O(to_level3[1071]),
   .I0(level4_in[6426]),
   .I1(level4_in[6427]),
   .I2(level4_in[6428]),
   .I3(level4_in[6429]),
   .I4(level4_in[6430]),
   .I5(level4_in[6431])
);

LUT6 #(
   .INIT(64'h1eae34621eae3462)  
) LUT6_inst8848 (
   .O(to_level3[1072]),
   .I0(level4_in[6432]),
   .I1(level4_in[6433]),
   .I2(level4_in[6434]),
   .I3(level4_in[6435]),
   .I4(level4_in[6436]),
   .I5(level4_in[6437])
);

LUT6 #(
   .INIT(64'h83f7752483f77524)  
) LUT6_inst8849 (
   .O(to_level3[1073]),
   .I0(level4_in[6438]),
   .I1(level4_in[6439]),
   .I2(level4_in[6440]),
   .I3(level4_in[6441]),
   .I4(level4_in[6442]),
   .I5(level4_in[6443])
);

LUT6 #(
   .INIT(64'h250f8fd0250f8fd0)  
) LUT6_inst8850 (
   .O(to_level3[1074]),
   .I0(level4_in[6444]),
   .I1(level4_in[6445]),
   .I2(level4_in[6446]),
   .I3(level4_in[6447]),
   .I4(level4_in[6448]),
   .I5(level4_in[6449])
);

LUT6 #(
   .INIT(64'h4be0f8ee4be0f8ee)  
) LUT6_inst8851 (
   .O(to_level3[1075]),
   .I0(level4_in[6450]),
   .I1(level4_in[6451]),
   .I2(level4_in[6452]),
   .I3(level4_in[6453]),
   .I4(level4_in[6454]),
   .I5(level4_in[6455])
);

LUT6 #(
   .INIT(64'h1b8039b51b8039b5)  
) LUT6_inst8852 (
   .O(to_level3[1076]),
   .I0(level4_in[6456]),
   .I1(level4_in[6457]),
   .I2(level4_in[6458]),
   .I3(level4_in[6459]),
   .I4(level4_in[6460]),
   .I5(level4_in[6461])
);

LUT6 #(
   .INIT(64'h73a3a21d73a3a21d)  
) LUT6_inst8853 (
   .O(to_level3[1077]),
   .I0(level4_in[6462]),
   .I1(level4_in[6463]),
   .I2(level4_in[6464]),
   .I3(level4_in[6465]),
   .I4(level4_in[6466]),
   .I5(level4_in[6467])
);

LUT6 #(
   .INIT(64'h7f97a3ed7f97a3ed)  
) LUT6_inst8854 (
   .O(to_level3[1078]),
   .I0(level4_in[6468]),
   .I1(level4_in[6469]),
   .I2(level4_in[6470]),
   .I3(level4_in[6471]),
   .I4(level4_in[6472]),
   .I5(level4_in[6473])
);

LUT6 #(
   .INIT(64'hb507bcbbb507bcbb)  
) LUT6_inst8855 (
   .O(to_level3[1079]),
   .I0(level4_in[6474]),
   .I1(level4_in[6475]),
   .I2(level4_in[6476]),
   .I3(level4_in[6477]),
   .I4(level4_in[6478]),
   .I5(level4_in[6479])
);

LUT6 #(
   .INIT(64'hcd29d3b2cd29d3b2)  
) LUT6_inst8856 (
   .O(to_level3[1080]),
   .I0(level4_in[6480]),
   .I1(level4_in[6481]),
   .I2(level4_in[6482]),
   .I3(level4_in[6483]),
   .I4(level4_in[6484]),
   .I5(level4_in[6485])
);

LUT6 #(
   .INIT(64'hb1c805b5b1c805b5)  
) LUT6_inst8857 (
   .O(to_level3[1081]),
   .I0(level4_in[6486]),
   .I1(level4_in[6487]),
   .I2(level4_in[6488]),
   .I3(level4_in[6489]),
   .I4(level4_in[6490]),
   .I5(level4_in[6491])
);

LUT6 #(
   .INIT(64'h3f9399143f939914)  
) LUT6_inst8858 (
   .O(to_level3[1082]),
   .I0(level4_in[6492]),
   .I1(level4_in[6493]),
   .I2(level4_in[6494]),
   .I3(level4_in[6495]),
   .I4(level4_in[6496]),
   .I5(level4_in[6497])
);

LUT6 #(
   .INIT(64'h16bd312e16bd312e)  
) LUT6_inst8859 (
   .O(to_level3[1083]),
   .I0(level4_in[6498]),
   .I1(level4_in[6499]),
   .I2(level4_in[6500]),
   .I3(level4_in[6501]),
   .I4(level4_in[6502]),
   .I5(level4_in[6503])
);

LUT6 #(
   .INIT(64'h5e016e715e016e71)  
) LUT6_inst8860 (
   .O(to_level3[1084]),
   .I0(level4_in[6504]),
   .I1(level4_in[6505]),
   .I2(level4_in[6506]),
   .I3(level4_in[6507]),
   .I4(level4_in[6508]),
   .I5(level4_in[6509])
);

LUT6 #(
   .INIT(64'h7b02ca507b02ca50)  
) LUT6_inst8861 (
   .O(to_level3[1085]),
   .I0(level4_in[6510]),
   .I1(level4_in[6511]),
   .I2(level4_in[6512]),
   .I3(level4_in[6513]),
   .I4(level4_in[6514]),
   .I5(level4_in[6515])
);

LUT6 #(
   .INIT(64'hb869dc4fb869dc4f)  
) LUT6_inst8862 (
   .O(to_level3[1086]),
   .I0(level4_in[6516]),
   .I1(level4_in[6517]),
   .I2(level4_in[6518]),
   .I3(level4_in[6519]),
   .I4(level4_in[6520]),
   .I5(level4_in[6521])
);

LUT6 #(
   .INIT(64'h0d1468f40d1468f4)  
) LUT6_inst8863 (
   .O(to_level3[1087]),
   .I0(level4_in[6522]),
   .I1(level4_in[6523]),
   .I2(level4_in[6524]),
   .I3(level4_in[6525]),
   .I4(level4_in[6526]),
   .I5(level4_in[6527])
);

LUT6 #(
   .INIT(64'h3e5897da3e5897da)  
) LUT6_inst8864 (
   .O(to_level3[1088]),
   .I0(level4_in[6528]),
   .I1(level4_in[6529]),
   .I2(level4_in[6530]),
   .I3(level4_in[6531]),
   .I4(level4_in[6532]),
   .I5(level4_in[6533])
);

LUT6 #(
   .INIT(64'h16c9cb3916c9cb39)  
) LUT6_inst8865 (
   .O(to_level3[1089]),
   .I0(level4_in[6534]),
   .I1(level4_in[6535]),
   .I2(level4_in[6536]),
   .I3(level4_in[6537]),
   .I4(level4_in[6538]),
   .I5(level4_in[6539])
);

LUT6 #(
   .INIT(64'h59b99a5959b99a59)  
) LUT6_inst8866 (
   .O(to_level3[1090]),
   .I0(level4_in[6540]),
   .I1(level4_in[6541]),
   .I2(level4_in[6542]),
   .I3(level4_in[6543]),
   .I4(level4_in[6544]),
   .I5(level4_in[6545])
);

LUT6 #(
   .INIT(64'h869a05d1869a05d1)  
) LUT6_inst8867 (
   .O(to_level3[1091]),
   .I0(level4_in[6546]),
   .I1(level4_in[6547]),
   .I2(level4_in[6548]),
   .I3(level4_in[6549]),
   .I4(level4_in[6550]),
   .I5(level4_in[6551])
);

LUT6 #(
   .INIT(64'hf87efc7df87efc7d)  
) LUT6_inst8868 (
   .O(to_level3[1092]),
   .I0(level4_in[6552]),
   .I1(level4_in[6553]),
   .I2(level4_in[6554]),
   .I3(level4_in[6555]),
   .I4(level4_in[6556]),
   .I5(level4_in[6557])
);

LUT6 #(
   .INIT(64'hefbf845defbf845d)  
) LUT6_inst8869 (
   .O(to_level3[1093]),
   .I0(level4_in[6558]),
   .I1(level4_in[6559]),
   .I2(level4_in[6560]),
   .I3(level4_in[6561]),
   .I4(level4_in[6562]),
   .I5(level4_in[6563])
);

LUT6 #(
   .INIT(64'hd7bf90f5d7bf90f5)  
) LUT6_inst8870 (
   .O(to_level3[1094]),
   .I0(level4_in[6564]),
   .I1(level4_in[6565]),
   .I2(level4_in[6566]),
   .I3(level4_in[6567]),
   .I4(level4_in[6568]),
   .I5(level4_in[6569])
);

LUT6 #(
   .INIT(64'h90186c4f90186c4f)  
) LUT6_inst8871 (
   .O(to_level3[1095]),
   .I0(level4_in[6570]),
   .I1(level4_in[6571]),
   .I2(level4_in[6572]),
   .I3(level4_in[6573]),
   .I4(level4_in[6574]),
   .I5(level4_in[6575])
);

LUT6 #(
   .INIT(64'h5d3fa92d5d3fa92d)  
) LUT6_inst8872 (
   .O(to_level3[1096]),
   .I0(level4_in[6576]),
   .I1(level4_in[6577]),
   .I2(level4_in[6578]),
   .I3(level4_in[6579]),
   .I4(level4_in[6580]),
   .I5(level4_in[6581])
);

LUT6 #(
   .INIT(64'hadc630eeadc630ee)  
) LUT6_inst8873 (
   .O(to_level3[1097]),
   .I0(level4_in[6582]),
   .I1(level4_in[6583]),
   .I2(level4_in[6584]),
   .I3(level4_in[6585]),
   .I4(level4_in[6586]),
   .I5(level4_in[6587])
);

LUT6 #(
   .INIT(64'he1f64bc7e1f64bc7)  
) LUT6_inst8874 (
   .O(to_level3[1098]),
   .I0(level4_in[6588]),
   .I1(level4_in[6589]),
   .I2(level4_in[6590]),
   .I3(level4_in[6591]),
   .I4(level4_in[6592]),
   .I5(level4_in[6593])
);

LUT6 #(
   .INIT(64'h68d580c968d580c9)  
) LUT6_inst8875 (
   .O(to_level3[1099]),
   .I0(level4_in[6594]),
   .I1(level4_in[6595]),
   .I2(level4_in[6596]),
   .I3(level4_in[6597]),
   .I4(level4_in[6598]),
   .I5(level4_in[6599])
);

LUT6 #(
   .INIT(64'h08d16e7208d16e72)  
) LUT6_inst8876 (
   .O(to_level3[1100]),
   .I0(level4_in[6600]),
   .I1(level4_in[6601]),
   .I2(level4_in[6602]),
   .I3(level4_in[6603]),
   .I4(level4_in[6604]),
   .I5(level4_in[6605])
);

LUT6 #(
   .INIT(64'h1f9aacb41f9aacb4)  
) LUT6_inst8877 (
   .O(to_level3[1101]),
   .I0(level4_in[6606]),
   .I1(level4_in[6607]),
   .I2(level4_in[6608]),
   .I3(level4_in[6609]),
   .I4(level4_in[6610]),
   .I5(level4_in[6611])
);

LUT6 #(
   .INIT(64'h7d64dc697d64dc69)  
) LUT6_inst8878 (
   .O(to_level3[1102]),
   .I0(level4_in[6612]),
   .I1(level4_in[6613]),
   .I2(level4_in[6614]),
   .I3(level4_in[6615]),
   .I4(level4_in[6616]),
   .I5(level4_in[6617])
);

LUT6 #(
   .INIT(64'h409506d1409506d1)  
) LUT6_inst8879 (
   .O(to_level3[1103]),
   .I0(level4_in[6618]),
   .I1(level4_in[6619]),
   .I2(level4_in[6620]),
   .I3(level4_in[6621]),
   .I4(level4_in[6622]),
   .I5(level4_in[6623])
);

LUT6 #(
   .INIT(64'h3c1aa9d83c1aa9d8)  
) LUT6_inst8880 (
   .O(to_level3[1104]),
   .I0(level4_in[6624]),
   .I1(level4_in[6625]),
   .I2(level4_in[6626]),
   .I3(level4_in[6627]),
   .I4(level4_in[6628]),
   .I5(level4_in[6629])
);

LUT6 #(
   .INIT(64'h1bf445ba1bf445ba)  
) LUT6_inst8881 (
   .O(to_level3[1105]),
   .I0(level4_in[6630]),
   .I1(level4_in[6631]),
   .I2(level4_in[6632]),
   .I3(level4_in[6633]),
   .I4(level4_in[6634]),
   .I5(level4_in[6635])
);

LUT6 #(
   .INIT(64'hbc6b0f2abc6b0f2a)  
) LUT6_inst8882 (
   .O(to_level3[1106]),
   .I0(level4_in[6636]),
   .I1(level4_in[6637]),
   .I2(level4_in[6638]),
   .I3(level4_in[6639]),
   .I4(level4_in[6640]),
   .I5(level4_in[6641])
);

LUT6 #(
   .INIT(64'hd46754add46754ad)  
) LUT6_inst8883 (
   .O(to_level3[1107]),
   .I0(level4_in[6642]),
   .I1(level4_in[6643]),
   .I2(level4_in[6644]),
   .I3(level4_in[6645]),
   .I4(level4_in[6646]),
   .I5(level4_in[6647])
);

LUT6 #(
   .INIT(64'h06f988b106f988b1)  
) LUT6_inst8884 (
   .O(to_level3[1108]),
   .I0(level4_in[6648]),
   .I1(level4_in[6649]),
   .I2(level4_in[6650]),
   .I3(level4_in[6651]),
   .I4(level4_in[6652]),
   .I5(level4_in[6653])
);

LUT6 #(
   .INIT(64'hc23c5891c23c5891)  
) LUT6_inst8885 (
   .O(to_level3[1109]),
   .I0(level4_in[6654]),
   .I1(level4_in[6655]),
   .I2(level4_in[6656]),
   .I3(level4_in[6657]),
   .I4(level4_in[6658]),
   .I5(level4_in[6659])
);

LUT6 #(
   .INIT(64'hd4ba466ed4ba466e)  
) LUT6_inst8886 (
   .O(to_level3[1110]),
   .I0(level4_in[6660]),
   .I1(level4_in[6661]),
   .I2(level4_in[6662]),
   .I3(level4_in[6663]),
   .I4(level4_in[6664]),
   .I5(level4_in[6665])
);

LUT6 #(
   .INIT(64'ha8b84e66a8b84e66)  
) LUT6_inst8887 (
   .O(to_level3[1111]),
   .I0(level4_in[6666]),
   .I1(level4_in[6667]),
   .I2(level4_in[6668]),
   .I3(level4_in[6669]),
   .I4(level4_in[6670]),
   .I5(level4_in[6671])
);

LUT6 #(
   .INIT(64'hc8fddd61c8fddd61)  
) LUT6_inst8888 (
   .O(to_level3[1112]),
   .I0(level4_in[6672]),
   .I1(level4_in[6673]),
   .I2(level4_in[6674]),
   .I3(level4_in[6675]),
   .I4(level4_in[6676]),
   .I5(level4_in[6677])
);

LUT6 #(
   .INIT(64'h5c12820c5c12820c)  
) LUT6_inst8889 (
   .O(to_level3[1113]),
   .I0(level4_in[6678]),
   .I1(level4_in[6679]),
   .I2(level4_in[6680]),
   .I3(level4_in[6681]),
   .I4(level4_in[6682]),
   .I5(level4_in[6683])
);

LUT6 #(
   .INIT(64'h468c9f8c468c9f8c)  
) LUT6_inst8890 (
   .O(to_level3[1114]),
   .I0(level4_in[6684]),
   .I1(level4_in[6685]),
   .I2(level4_in[6686]),
   .I3(level4_in[6687]),
   .I4(level4_in[6688]),
   .I5(level4_in[6689])
);

LUT6 #(
   .INIT(64'h978f8b5c978f8b5c)  
) LUT6_inst8891 (
   .O(to_level3[1115]),
   .I0(level4_in[6690]),
   .I1(level4_in[6691]),
   .I2(level4_in[6692]),
   .I3(level4_in[6693]),
   .I4(level4_in[6694]),
   .I5(level4_in[6695])
);

LUT6 #(
   .INIT(64'hf0ffd722f0ffd722)  
) LUT6_inst8892 (
   .O(to_level3[1116]),
   .I0(level4_in[6696]),
   .I1(level4_in[6697]),
   .I2(level4_in[6698]),
   .I3(level4_in[6699]),
   .I4(level4_in[6700]),
   .I5(level4_in[6701])
);

LUT6 #(
   .INIT(64'h4a9763844a976384)  
) LUT6_inst8893 (
   .O(to_level3[1117]),
   .I0(level4_in[6702]),
   .I1(level4_in[6703]),
   .I2(level4_in[6704]),
   .I3(level4_in[6705]),
   .I4(level4_in[6706]),
   .I5(level4_in[6707])
);

LUT6 #(
   .INIT(64'h8c7adc808c7adc80)  
) LUT6_inst8894 (
   .O(to_level3[1118]),
   .I0(level4_in[6708]),
   .I1(level4_in[6709]),
   .I2(level4_in[6710]),
   .I3(level4_in[6711]),
   .I4(level4_in[6712]),
   .I5(level4_in[6713])
);

LUT6 #(
   .INIT(64'h9813625198136251)  
) LUT6_inst8895 (
   .O(to_level3[1119]),
   .I0(level4_in[6714]),
   .I1(level4_in[6715]),
   .I2(level4_in[6716]),
   .I3(level4_in[6717]),
   .I4(level4_in[6718]),
   .I5(level4_in[6719])
);

LUT6 #(
   .INIT(64'h3336c6f43336c6f4)  
) LUT6_inst8896 (
   .O(to_level3[1120]),
   .I0(level4_in[6720]),
   .I1(level4_in[6721]),
   .I2(level4_in[6722]),
   .I3(level4_in[6723]),
   .I4(level4_in[6724]),
   .I5(level4_in[6725])
);

LUT6 #(
   .INIT(64'h1445f9b81445f9b8)  
) LUT6_inst8897 (
   .O(to_level3[1121]),
   .I0(level4_in[6726]),
   .I1(level4_in[6727]),
   .I2(level4_in[6728]),
   .I3(level4_in[6729]),
   .I4(level4_in[6730]),
   .I5(level4_in[6731])
);

LUT6 #(
   .INIT(64'h66694daa66694daa)  
) LUT6_inst8898 (
   .O(to_level3[1122]),
   .I0(level4_in[6732]),
   .I1(level4_in[6733]),
   .I2(level4_in[6734]),
   .I3(level4_in[6735]),
   .I4(level4_in[6736]),
   .I5(level4_in[6737])
);

LUT6 #(
   .INIT(64'hd714c95ed714c95e)  
) LUT6_inst8899 (
   .O(to_level3[1123]),
   .I0(level4_in[6738]),
   .I1(level4_in[6739]),
   .I2(level4_in[6740]),
   .I3(level4_in[6741]),
   .I4(level4_in[6742]),
   .I5(level4_in[6743])
);

LUT6 #(
   .INIT(64'h5e634cf85e634cf8)  
) LUT6_inst8900 (
   .O(to_level3[1124]),
   .I0(level4_in[6744]),
   .I1(level4_in[6745]),
   .I2(level4_in[6746]),
   .I3(level4_in[6747]),
   .I4(level4_in[6748]),
   .I5(level4_in[6749])
);

LUT6 #(
   .INIT(64'h8d14f3c88d14f3c8)  
) LUT6_inst8901 (
   .O(to_level3[1125]),
   .I0(level4_in[6750]),
   .I1(level4_in[6751]),
   .I2(level4_in[6752]),
   .I3(level4_in[6753]),
   .I4(level4_in[6754]),
   .I5(level4_in[6755])
);

LUT6 #(
   .INIT(64'hbfd914b1bfd914b1)  
) LUT6_inst8902 (
   .O(to_level3[1126]),
   .I0(level4_in[6756]),
   .I1(level4_in[6757]),
   .I2(level4_in[6758]),
   .I3(level4_in[6759]),
   .I4(level4_in[6760]),
   .I5(level4_in[6761])
);

LUT6 #(
   .INIT(64'h9cb1494f9cb1494f)  
) LUT6_inst8903 (
   .O(to_level3[1127]),
   .I0(level4_in[6762]),
   .I1(level4_in[6763]),
   .I2(level4_in[6764]),
   .I3(level4_in[6765]),
   .I4(level4_in[6766]),
   .I5(level4_in[6767])
);

LUT6 #(
   .INIT(64'h47b8bb0647b8bb06)  
) LUT6_inst8904 (
   .O(to_level3[1128]),
   .I0(level4_in[6768]),
   .I1(level4_in[6769]),
   .I2(level4_in[6770]),
   .I3(level4_in[6771]),
   .I4(level4_in[6772]),
   .I5(level4_in[6773])
);

LUT6 #(
   .INIT(64'h6f59f11d6f59f11d)  
) LUT6_inst8905 (
   .O(to_level3[1129]),
   .I0(level4_in[6774]),
   .I1(level4_in[6775]),
   .I2(level4_in[6776]),
   .I3(level4_in[6777]),
   .I4(level4_in[6778]),
   .I5(level4_in[6779])
);

LUT6 #(
   .INIT(64'h8897e2bc8897e2bc)  
) LUT6_inst8906 (
   .O(to_level3[1130]),
   .I0(level4_in[6780]),
   .I1(level4_in[6781]),
   .I2(level4_in[6782]),
   .I3(level4_in[6783]),
   .I4(level4_in[6784]),
   .I5(level4_in[6785])
);

LUT6 #(
   .INIT(64'h537629c5537629c5)  
) LUT6_inst8907 (
   .O(to_level3[1131]),
   .I0(level4_in[6786]),
   .I1(level4_in[6787]),
   .I2(level4_in[6788]),
   .I3(level4_in[6789]),
   .I4(level4_in[6790]),
   .I5(level4_in[6791])
);

LUT6 #(
   .INIT(64'h2e9e340a2e9e340a)  
) LUT6_inst8908 (
   .O(to_level3[1132]),
   .I0(level4_in[6792]),
   .I1(level4_in[6793]),
   .I2(level4_in[6794]),
   .I3(level4_in[6795]),
   .I4(level4_in[6796]),
   .I5(level4_in[6797])
);

LUT6 #(
   .INIT(64'hddc5e3e0ddc5e3e0)  
) LUT6_inst8909 (
   .O(to_level3[1133]),
   .I0(level4_in[6798]),
   .I1(level4_in[6799]),
   .I2(level4_in[6800]),
   .I3(level4_in[6801]),
   .I4(level4_in[6802]),
   .I5(level4_in[6803])
);

LUT6 #(
   .INIT(64'h0dbf2b5c0dbf2b5c)  
) LUT6_inst8910 (
   .O(to_level3[1134]),
   .I0(level4_in[6804]),
   .I1(level4_in[6805]),
   .I2(level4_in[6806]),
   .I3(level4_in[6807]),
   .I4(level4_in[6808]),
   .I5(level4_in[6809])
);

LUT6 #(
   .INIT(64'h9548417495484174)  
) LUT6_inst8911 (
   .O(to_level3[1135]),
   .I0(level4_in[6810]),
   .I1(level4_in[6811]),
   .I2(level4_in[6812]),
   .I3(level4_in[6813]),
   .I4(level4_in[6814]),
   .I5(level4_in[6815])
);

LUT6 #(
   .INIT(64'h4ae05cb44ae05cb4)  
) LUT6_inst8912 (
   .O(to_level3[1136]),
   .I0(level4_in[6816]),
   .I1(level4_in[6817]),
   .I2(level4_in[6818]),
   .I3(level4_in[6819]),
   .I4(level4_in[6820]),
   .I5(level4_in[6821])
);

LUT6 #(
   .INIT(64'hd2769b20d2769b20)  
) LUT6_inst8913 (
   .O(to_level3[1137]),
   .I0(level4_in[6822]),
   .I1(level4_in[6823]),
   .I2(level4_in[6824]),
   .I3(level4_in[6825]),
   .I4(level4_in[6826]),
   .I5(level4_in[6827])
);

LUT6 #(
   .INIT(64'h8206c1618206c161)  
) LUT6_inst8914 (
   .O(to_level3[1138]),
   .I0(level4_in[6828]),
   .I1(level4_in[6829]),
   .I2(level4_in[6830]),
   .I3(level4_in[6831]),
   .I4(level4_in[6832]),
   .I5(level4_in[6833])
);

LUT6 #(
   .INIT(64'h317b4c06317b4c06)  
) LUT6_inst8915 (
   .O(to_level3[1139]),
   .I0(level4_in[6834]),
   .I1(level4_in[6835]),
   .I2(level4_in[6836]),
   .I3(level4_in[6837]),
   .I4(level4_in[6838]),
   .I5(level4_in[6839])
);

LUT6 #(
   .INIT(64'h090083b9090083b9)  
) LUT6_inst8916 (
   .O(to_level3[1140]),
   .I0(level4_in[6840]),
   .I1(level4_in[6841]),
   .I2(level4_in[6842]),
   .I3(level4_in[6843]),
   .I4(level4_in[6844]),
   .I5(level4_in[6845])
);

LUT6 #(
   .INIT(64'hf1045af3f1045af3)  
) LUT6_inst8917 (
   .O(to_level3[1141]),
   .I0(level4_in[6846]),
   .I1(level4_in[6847]),
   .I2(level4_in[6848]),
   .I3(level4_in[6849]),
   .I4(level4_in[6850]),
   .I5(level4_in[6851])
);

LUT6 #(
   .INIT(64'h9150776391507763)  
) LUT6_inst8918 (
   .O(to_level3[1142]),
   .I0(level4_in[6852]),
   .I1(level4_in[6853]),
   .I2(level4_in[6854]),
   .I3(level4_in[6855]),
   .I4(level4_in[6856]),
   .I5(level4_in[6857])
);

LUT6 #(
   .INIT(64'h1ec142cb1ec142cb)  
) LUT6_inst8919 (
   .O(to_level3[1143]),
   .I0(level4_in[6858]),
   .I1(level4_in[6859]),
   .I2(level4_in[6860]),
   .I3(level4_in[6861]),
   .I4(level4_in[6862]),
   .I5(level4_in[6863])
);

LUT6 #(
   .INIT(64'hf5b2c093f5b2c093)  
) LUT6_inst8920 (
   .O(to_level3[1144]),
   .I0(level4_in[6864]),
   .I1(level4_in[6865]),
   .I2(level4_in[6866]),
   .I3(level4_in[6867]),
   .I4(level4_in[6868]),
   .I5(level4_in[6869])
);

LUT6 #(
   .INIT(64'h8866413188664131)  
) LUT6_inst8921 (
   .O(to_level3[1145]),
   .I0(level4_in[6870]),
   .I1(level4_in[6871]),
   .I2(level4_in[6872]),
   .I3(level4_in[6873]),
   .I4(level4_in[6874]),
   .I5(level4_in[6875])
);

LUT6 #(
   .INIT(64'hc04b91efc04b91ef)  
) LUT6_inst8922 (
   .O(to_level3[1146]),
   .I0(level4_in[6876]),
   .I1(level4_in[6877]),
   .I2(level4_in[6878]),
   .I3(level4_in[6879]),
   .I4(level4_in[6880]),
   .I5(level4_in[6881])
);

LUT6 #(
   .INIT(64'h3e753d233e753d23)  
) LUT6_inst8923 (
   .O(to_level3[1147]),
   .I0(level4_in[6882]),
   .I1(level4_in[6883]),
   .I2(level4_in[6884]),
   .I3(level4_in[6885]),
   .I4(level4_in[6886]),
   .I5(level4_in[6887])
);

LUT6 #(
   .INIT(64'hddf2c5cfddf2c5cf)  
) LUT6_inst8924 (
   .O(to_level3[1148]),
   .I0(level4_in[6888]),
   .I1(level4_in[6889]),
   .I2(level4_in[6890]),
   .I3(level4_in[6891]),
   .I4(level4_in[6892]),
   .I5(level4_in[6893])
);

LUT6 #(
   .INIT(64'h4ae113b54ae113b5)  
) LUT6_inst8925 (
   .O(to_level3[1149]),
   .I0(level4_in[6894]),
   .I1(level4_in[6895]),
   .I2(level4_in[6896]),
   .I3(level4_in[6897]),
   .I4(level4_in[6898]),
   .I5(level4_in[6899])
);

LUT6 #(
   .INIT(64'h0b8525430b852543)  
) LUT6_inst8926 (
   .O(to_level3[1150]),
   .I0(level4_in[6900]),
   .I1(level4_in[6901]),
   .I2(level4_in[6902]),
   .I3(level4_in[6903]),
   .I4(level4_in[6904]),
   .I5(level4_in[6905])
);

LUT6 #(
   .INIT(64'hf9f0a958f9f0a958)  
) LUT6_inst8927 (
   .O(to_level3[1151]),
   .I0(level4_in[6906]),
   .I1(level4_in[6907]),
   .I2(level4_in[6908]),
   .I3(level4_in[6909]),
   .I4(level4_in[6910]),
   .I5(level4_in[6911])
);

LUT6 #(
   .INIT(64'h9b7ac7af9b7ac7af)  
) LUT6_inst8928 (
   .O(to_level3[1152]),
   .I0(level4_in[6912]),
   .I1(level4_in[6913]),
   .I2(level4_in[6914]),
   .I3(level4_in[6915]),
   .I4(level4_in[6916]),
   .I5(level4_in[6917])
);

LUT6 #(
   .INIT(64'hf5421223f5421223)  
) LUT6_inst8929 (
   .O(to_level3[1153]),
   .I0(level4_in[6918]),
   .I1(level4_in[6919]),
   .I2(level4_in[6920]),
   .I3(level4_in[6921]),
   .I4(level4_in[6922]),
   .I5(level4_in[6923])
);

LUT6 #(
   .INIT(64'h3866c7e53866c7e5)  
) LUT6_inst8930 (
   .O(to_level3[1154]),
   .I0(level4_in[6924]),
   .I1(level4_in[6925]),
   .I2(level4_in[6926]),
   .I3(level4_in[6927]),
   .I4(level4_in[6928]),
   .I5(level4_in[6929])
);

LUT6 #(
   .INIT(64'h9149b0949149b094)  
) LUT6_inst8931 (
   .O(to_level3[1155]),
   .I0(level4_in[6930]),
   .I1(level4_in[6931]),
   .I2(level4_in[6932]),
   .I3(level4_in[6933]),
   .I4(level4_in[6934]),
   .I5(level4_in[6935])
);

LUT6 #(
   .INIT(64'h3113cc7b3113cc7b)  
) LUT6_inst8932 (
   .O(to_level3[1156]),
   .I0(level4_in[6936]),
   .I1(level4_in[6937]),
   .I2(level4_in[6938]),
   .I3(level4_in[6939]),
   .I4(level4_in[6940]),
   .I5(level4_in[6941])
);

LUT6 #(
   .INIT(64'h9fc642209fc64220)  
) LUT6_inst8933 (
   .O(to_level3[1157]),
   .I0(level4_in[6942]),
   .I1(level4_in[6943]),
   .I2(level4_in[6944]),
   .I3(level4_in[6945]),
   .I4(level4_in[6946]),
   .I5(level4_in[6947])
);

LUT6 #(
   .INIT(64'h8482ccfd8482ccfd)  
) LUT6_inst8934 (
   .O(to_level3[1158]),
   .I0(level4_in[6948]),
   .I1(level4_in[6949]),
   .I2(level4_in[6950]),
   .I3(level4_in[6951]),
   .I4(level4_in[6952]),
   .I5(level4_in[6953])
);

LUT6 #(
   .INIT(64'ha0c13ef7a0c13ef7)  
) LUT6_inst8935 (
   .O(to_level3[1159]),
   .I0(level4_in[6954]),
   .I1(level4_in[6955]),
   .I2(level4_in[6956]),
   .I3(level4_in[6957]),
   .I4(level4_in[6958]),
   .I5(level4_in[6959])
);

LUT6 #(
   .INIT(64'hf82e6a7ff82e6a7f)  
) LUT6_inst8936 (
   .O(to_level3[1160]),
   .I0(level4_in[6960]),
   .I1(level4_in[6961]),
   .I2(level4_in[6962]),
   .I3(level4_in[6963]),
   .I4(level4_in[6964]),
   .I5(level4_in[6965])
);

LUT6 #(
   .INIT(64'h47f5784647f57846)  
) LUT6_inst8937 (
   .O(to_level3[1161]),
   .I0(level4_in[6966]),
   .I1(level4_in[6967]),
   .I2(level4_in[6968]),
   .I3(level4_in[6969]),
   .I4(level4_in[6970]),
   .I5(level4_in[6971])
);

LUT6 #(
   .INIT(64'h37fb1aaa37fb1aaa)  
) LUT6_inst8938 (
   .O(to_level3[1162]),
   .I0(level4_in[6972]),
   .I1(level4_in[6973]),
   .I2(level4_in[6974]),
   .I3(level4_in[6975]),
   .I4(level4_in[6976]),
   .I5(level4_in[6977])
);

LUT6 #(
   .INIT(64'hf837bf77f837bf77)  
) LUT6_inst8939 (
   .O(to_level3[1163]),
   .I0(level4_in[6978]),
   .I1(level4_in[6979]),
   .I2(level4_in[6980]),
   .I3(level4_in[6981]),
   .I4(level4_in[6982]),
   .I5(level4_in[6983])
);

LUT6 #(
   .INIT(64'h247cf6b9247cf6b9)  
) LUT6_inst8940 (
   .O(to_level3[1164]),
   .I0(level4_in[6984]),
   .I1(level4_in[6985]),
   .I2(level4_in[6986]),
   .I3(level4_in[6987]),
   .I4(level4_in[6988]),
   .I5(level4_in[6989])
);

LUT6 #(
   .INIT(64'h42b4c60542b4c605)  
) LUT6_inst8941 (
   .O(to_level3[1165]),
   .I0(level4_in[6990]),
   .I1(level4_in[6991]),
   .I2(level4_in[6992]),
   .I3(level4_in[6993]),
   .I4(level4_in[6994]),
   .I5(level4_in[6995])
);

LUT6 #(
   .INIT(64'hce2058edce2058ed)  
) LUT6_inst8942 (
   .O(to_level3[1166]),
   .I0(level4_in[6996]),
   .I1(level4_in[6997]),
   .I2(level4_in[6998]),
   .I3(level4_in[6999]),
   .I4(level4_in[7000]),
   .I5(level4_in[7001])
);

LUT6 #(
   .INIT(64'h35e75fec35e75fec)  
) LUT6_inst8943 (
   .O(to_level3[1167]),
   .I0(level4_in[7002]),
   .I1(level4_in[7003]),
   .I2(level4_in[7004]),
   .I3(level4_in[7005]),
   .I4(level4_in[7006]),
   .I5(level4_in[7007])
);

LUT6 #(
   .INIT(64'h502a673e502a673e)  
) LUT6_inst8944 (
   .O(to_level3[1168]),
   .I0(level4_in[7008]),
   .I1(level4_in[7009]),
   .I2(level4_in[7010]),
   .I3(level4_in[7011]),
   .I4(level4_in[7012]),
   .I5(level4_in[7013])
);

LUT6 #(
   .INIT(64'h0085529000855290)  
) LUT6_inst8945 (
   .O(to_level3[1169]),
   .I0(level4_in[7014]),
   .I1(level4_in[7015]),
   .I2(level4_in[7016]),
   .I3(level4_in[7017]),
   .I4(level4_in[7018]),
   .I5(level4_in[7019])
);

LUT6 #(
   .INIT(64'ha1ebcdbda1ebcdbd)  
) LUT6_inst8946 (
   .O(to_level3[1170]),
   .I0(level4_in[7020]),
   .I1(level4_in[7021]),
   .I2(level4_in[7022]),
   .I3(level4_in[7023]),
   .I4(level4_in[7024]),
   .I5(level4_in[7025])
);

LUT6 #(
   .INIT(64'h8a47fc258a47fc25)  
) LUT6_inst8947 (
   .O(to_level3[1171]),
   .I0(level4_in[7026]),
   .I1(level4_in[7027]),
   .I2(level4_in[7028]),
   .I3(level4_in[7029]),
   .I4(level4_in[7030]),
   .I5(level4_in[7031])
);

LUT6 #(
   .INIT(64'h2edf54c72edf54c7)  
) LUT6_inst8948 (
   .O(to_level3[1172]),
   .I0(level4_in[7032]),
   .I1(level4_in[7033]),
   .I2(level4_in[7034]),
   .I3(level4_in[7035]),
   .I4(level4_in[7036]),
   .I5(level4_in[7037])
);

LUT6 #(
   .INIT(64'h2925c26f2925c26f)  
) LUT6_inst8949 (
   .O(to_level3[1173]),
   .I0(level4_in[7038]),
   .I1(level4_in[7039]),
   .I2(level4_in[7040]),
   .I3(level4_in[7041]),
   .I4(level4_in[7042]),
   .I5(level4_in[7043])
);

LUT6 #(
   .INIT(64'hc19260f6c19260f6)  
) LUT6_inst8950 (
   .O(to_level3[1174]),
   .I0(level4_in[7044]),
   .I1(level4_in[7045]),
   .I2(level4_in[7046]),
   .I3(level4_in[7047]),
   .I4(level4_in[7048]),
   .I5(level4_in[7049])
);

LUT6 #(
   .INIT(64'h035df2e4035df2e4)  
) LUT6_inst8951 (
   .O(to_level3[1175]),
   .I0(level4_in[7050]),
   .I1(level4_in[7051]),
   .I2(level4_in[7052]),
   .I3(level4_in[7053]),
   .I4(level4_in[7054]),
   .I5(level4_in[7055])
);

LUT6 #(
   .INIT(64'h7c61f6517c61f651)  
) LUT6_inst8952 (
   .O(to_level3[1176]),
   .I0(level4_in[7056]),
   .I1(level4_in[7057]),
   .I2(level4_in[7058]),
   .I3(level4_in[7059]),
   .I4(level4_in[7060]),
   .I5(level4_in[7061])
);

LUT6 #(
   .INIT(64'h5edf4a7e5edf4a7e)  
) LUT6_inst8953 (
   .O(to_level3[1177]),
   .I0(level4_in[7062]),
   .I1(level4_in[7063]),
   .I2(level4_in[7064]),
   .I3(level4_in[7065]),
   .I4(level4_in[7066]),
   .I5(level4_in[7067])
);

LUT6 #(
   .INIT(64'hf6dbb966f6dbb966)  
) LUT6_inst8954 (
   .O(to_level3[1178]),
   .I0(level4_in[7068]),
   .I1(level4_in[7069]),
   .I2(level4_in[7070]),
   .I3(level4_in[7071]),
   .I4(level4_in[7072]),
   .I5(level4_in[7073])
);

LUT6 #(
   .INIT(64'h149871bf149871bf)  
) LUT6_inst8955 (
   .O(to_level3[1179]),
   .I0(level4_in[7074]),
   .I1(level4_in[7075]),
   .I2(level4_in[7076]),
   .I3(level4_in[7077]),
   .I4(level4_in[7078]),
   .I5(level4_in[7079])
);

LUT6 #(
   .INIT(64'h3e42337f3e42337f)  
) LUT6_inst8956 (
   .O(to_level3[1180]),
   .I0(level4_in[7080]),
   .I1(level4_in[7081]),
   .I2(level4_in[7082]),
   .I3(level4_in[7083]),
   .I4(level4_in[7084]),
   .I5(level4_in[7085])
);

LUT6 #(
   .INIT(64'h861af3de861af3de)  
) LUT6_inst8957 (
   .O(to_level3[1181]),
   .I0(level4_in[7086]),
   .I1(level4_in[7087]),
   .I2(level4_in[7088]),
   .I3(level4_in[7089]),
   .I4(level4_in[7090]),
   .I5(level4_in[7091])
);

LUT6 #(
   .INIT(64'h4fc3f1a24fc3f1a2)  
) LUT6_inst8958 (
   .O(to_level3[1182]),
   .I0(level4_in[7092]),
   .I1(level4_in[7093]),
   .I2(level4_in[7094]),
   .I3(level4_in[7095]),
   .I4(level4_in[7096]),
   .I5(level4_in[7097])
);

LUT6 #(
   .INIT(64'h1bd757311bd75731)  
) LUT6_inst8959 (
   .O(to_level3[1183]),
   .I0(level4_in[7098]),
   .I1(level4_in[7099]),
   .I2(level4_in[7100]),
   .I3(level4_in[7101]),
   .I4(level4_in[7102]),
   .I5(level4_in[7103])
);

LUT6 #(
   .INIT(64'h9140a6e69140a6e6)  
) LUT6_inst8960 (
   .O(to_level3[1184]),
   .I0(level4_in[7104]),
   .I1(level4_in[7105]),
   .I2(level4_in[7106]),
   .I3(level4_in[7107]),
   .I4(level4_in[7108]),
   .I5(level4_in[7109])
);

LUT6 #(
   .INIT(64'hc4f941a5c4f941a5)  
) LUT6_inst8961 (
   .O(to_level3[1185]),
   .I0(level4_in[7110]),
   .I1(level4_in[7111]),
   .I2(level4_in[7112]),
   .I3(level4_in[7113]),
   .I4(level4_in[7114]),
   .I5(level4_in[7115])
);

LUT6 #(
   .INIT(64'hf8c92052f8c92052)  
) LUT6_inst8962 (
   .O(to_level3[1186]),
   .I0(level4_in[7116]),
   .I1(level4_in[7117]),
   .I2(level4_in[7118]),
   .I3(level4_in[7119]),
   .I4(level4_in[7120]),
   .I5(level4_in[7121])
);

LUT6 #(
   .INIT(64'hcc32e3bbcc32e3bb)  
) LUT6_inst8963 (
   .O(to_level3[1187]),
   .I0(level4_in[7122]),
   .I1(level4_in[7123]),
   .I2(level4_in[7124]),
   .I3(level4_in[7125]),
   .I4(level4_in[7126]),
   .I5(level4_in[7127])
);

LUT6 #(
   .INIT(64'heb879722eb879722)  
) LUT6_inst8964 (
   .O(to_level3[1188]),
   .I0(level4_in[7128]),
   .I1(level4_in[7129]),
   .I2(level4_in[7130]),
   .I3(level4_in[7131]),
   .I4(level4_in[7132]),
   .I5(level4_in[7133])
);

LUT6 #(
   .INIT(64'h30ed9dae30ed9dae)  
) LUT6_inst8965 (
   .O(to_level3[1189]),
   .I0(level4_in[7134]),
   .I1(level4_in[7135]),
   .I2(level4_in[7136]),
   .I3(level4_in[7137]),
   .I4(level4_in[7138]),
   .I5(level4_in[7139])
);

LUT6 #(
   .INIT(64'h61d5b0e461d5b0e4)  
) LUT6_inst8966 (
   .O(to_level3[1190]),
   .I0(level4_in[7140]),
   .I1(level4_in[7141]),
   .I2(level4_in[7142]),
   .I3(level4_in[7143]),
   .I4(level4_in[7144]),
   .I5(level4_in[7145])
);

LUT6 #(
   .INIT(64'hd7505480d7505480)  
) LUT6_inst8967 (
   .O(to_level3[1191]),
   .I0(level4_in[7146]),
   .I1(level4_in[7147]),
   .I2(level4_in[7148]),
   .I3(level4_in[7149]),
   .I4(level4_in[7150]),
   .I5(level4_in[7151])
);

LUT6 #(
   .INIT(64'h8aacc1928aacc192)  
) LUT6_inst8968 (
   .O(to_level3[1192]),
   .I0(level4_in[7152]),
   .I1(level4_in[7153]),
   .I2(level4_in[7154]),
   .I3(level4_in[7155]),
   .I4(level4_in[7156]),
   .I5(level4_in[7157])
);

LUT6 #(
   .INIT(64'h5eb1cf955eb1cf95)  
) LUT6_inst8969 (
   .O(to_level3[1193]),
   .I0(level4_in[7158]),
   .I1(level4_in[7159]),
   .I2(level4_in[7160]),
   .I3(level4_in[7161]),
   .I4(level4_in[7162]),
   .I5(level4_in[7163])
);

LUT6 #(
   .INIT(64'h264cecb9264cecb9)  
) LUT6_inst8970 (
   .O(to_level3[1194]),
   .I0(level4_in[7164]),
   .I1(level4_in[7165]),
   .I2(level4_in[7166]),
   .I3(level4_in[7167]),
   .I4(level4_in[7168]),
   .I5(level4_in[7169])
);

LUT6 #(
   .INIT(64'h52536b0a52536b0a)  
) LUT6_inst8971 (
   .O(to_level3[1195]),
   .I0(level4_in[7170]),
   .I1(level4_in[7171]),
   .I2(level4_in[7172]),
   .I3(level4_in[7173]),
   .I4(level4_in[7174]),
   .I5(level4_in[7175])
);

LUT6 #(
   .INIT(64'h24b5dc9924b5dc99)  
) LUT6_inst8972 (
   .O(to_level3[1196]),
   .I0(level4_in[7176]),
   .I1(level4_in[7177]),
   .I2(level4_in[7178]),
   .I3(level4_in[7179]),
   .I4(level4_in[7180]),
   .I5(level4_in[7181])
);

LUT6 #(
   .INIT(64'h98af7e4f98af7e4f)  
) LUT6_inst8973 (
   .O(to_level3[1197]),
   .I0(level4_in[7182]),
   .I1(level4_in[7183]),
   .I2(level4_in[7184]),
   .I3(level4_in[7185]),
   .I4(level4_in[7186]),
   .I5(level4_in[7187])
);

LUT6 #(
   .INIT(64'hd9b29c28d9b29c28)  
) LUT6_inst8974 (
   .O(to_level3[1198]),
   .I0(level4_in[7188]),
   .I1(level4_in[7189]),
   .I2(level4_in[7190]),
   .I3(level4_in[7191]),
   .I4(level4_in[7192]),
   .I5(level4_in[7193])
);

LUT6 #(
   .INIT(64'h4b9c68354b9c6835)  
) LUT6_inst8975 (
   .O(to_level3[1199]),
   .I0(level4_in[7194]),
   .I1(level4_in[7195]),
   .I2(level4_in[7196]),
   .I3(level4_in[7197]),
   .I4(level4_in[7198]),
   .I5(level4_in[7199])
);

LUT6 #(
   .INIT(64'h8901f4518901f451)  
) LUT6_inst8976 (
   .O(to_level3[1200]),
   .I0(level4_in[7200]),
   .I1(level4_in[7201]),
   .I2(level4_in[7202]),
   .I3(level4_in[7203]),
   .I4(level4_in[7204]),
   .I5(level4_in[7205])
);

LUT6 #(
   .INIT(64'hb15bc433b15bc433)  
) LUT6_inst8977 (
   .O(to_level3[1201]),
   .I0(level4_in[7206]),
   .I1(level4_in[7207]),
   .I2(level4_in[7208]),
   .I3(level4_in[7209]),
   .I4(level4_in[7210]),
   .I5(level4_in[7211])
);

LUT6 #(
   .INIT(64'h45434e4a45434e4a)  
) LUT6_inst8978 (
   .O(to_level3[1202]),
   .I0(level4_in[7212]),
   .I1(level4_in[7213]),
   .I2(level4_in[7214]),
   .I3(level4_in[7215]),
   .I4(level4_in[7216]),
   .I5(level4_in[7217])
);

LUT6 #(
   .INIT(64'heae47c33eae47c33)  
) LUT6_inst8979 (
   .O(to_level3[1203]),
   .I0(level4_in[7218]),
   .I1(level4_in[7219]),
   .I2(level4_in[7220]),
   .I3(level4_in[7221]),
   .I4(level4_in[7222]),
   .I5(level4_in[7223])
);

LUT6 #(
   .INIT(64'h907ef415907ef415)  
) LUT6_inst8980 (
   .O(to_level3[1204]),
   .I0(level4_in[7224]),
   .I1(level4_in[7225]),
   .I2(level4_in[7226]),
   .I3(level4_in[7227]),
   .I4(level4_in[7228]),
   .I5(level4_in[7229])
);

LUT6 #(
   .INIT(64'h75c9baed75c9baed)  
) LUT6_inst8981 (
   .O(to_level3[1205]),
   .I0(level4_in[7230]),
   .I1(level4_in[7231]),
   .I2(level4_in[7232]),
   .I3(level4_in[7233]),
   .I4(level4_in[7234]),
   .I5(level4_in[7235])
);

LUT6 #(
   .INIT(64'h9e9c1b409e9c1b40)  
) LUT6_inst8982 (
   .O(to_level3[1206]),
   .I0(level4_in[7236]),
   .I1(level4_in[7237]),
   .I2(level4_in[7238]),
   .I3(level4_in[7239]),
   .I4(level4_in[7240]),
   .I5(level4_in[7241])
);

LUT6 #(
   .INIT(64'hcf8559fbcf8559fb)  
) LUT6_inst8983 (
   .O(to_level3[1207]),
   .I0(level4_in[7242]),
   .I1(level4_in[7243]),
   .I2(level4_in[7244]),
   .I3(level4_in[7245]),
   .I4(level4_in[7246]),
   .I5(level4_in[7247])
);

LUT6 #(
   .INIT(64'h6a3458c76a3458c7)  
) LUT6_inst8984 (
   .O(to_level3[1208]),
   .I0(level4_in[7248]),
   .I1(level4_in[7249]),
   .I2(level4_in[7250]),
   .I3(level4_in[7251]),
   .I4(level4_in[7252]),
   .I5(level4_in[7253])
);

LUT6 #(
   .INIT(64'hf976c9ddf976c9dd)  
) LUT6_inst8985 (
   .O(to_level3[1209]),
   .I0(level4_in[7254]),
   .I1(level4_in[7255]),
   .I2(level4_in[7256]),
   .I3(level4_in[7257]),
   .I4(level4_in[7258]),
   .I5(level4_in[7259])
);

LUT6 #(
   .INIT(64'he174002ce174002c)  
) LUT6_inst8986 (
   .O(to_level3[1210]),
   .I0(level4_in[7260]),
   .I1(level4_in[7261]),
   .I2(level4_in[7262]),
   .I3(level4_in[7263]),
   .I4(level4_in[7264]),
   .I5(level4_in[7265])
);

LUT6 #(
   .INIT(64'h4324514843245148)  
) LUT6_inst8987 (
   .O(to_level3[1211]),
   .I0(level4_in[7266]),
   .I1(level4_in[7267]),
   .I2(level4_in[7268]),
   .I3(level4_in[7269]),
   .I4(level4_in[7270]),
   .I5(level4_in[7271])
);

LUT6 #(
   .INIT(64'h2ffa5c7e2ffa5c7e)  
) LUT6_inst8988 (
   .O(to_level3[1212]),
   .I0(level4_in[7272]),
   .I1(level4_in[7273]),
   .I2(level4_in[7274]),
   .I3(level4_in[7275]),
   .I4(level4_in[7276]),
   .I5(level4_in[7277])
);

LUT6 #(
   .INIT(64'h384d2d38384d2d38)  
) LUT6_inst8989 (
   .O(to_level3[1213]),
   .I0(level4_in[7278]),
   .I1(level4_in[7279]),
   .I2(level4_in[7280]),
   .I3(level4_in[7281]),
   .I4(level4_in[7282]),
   .I5(level4_in[7283])
);

LUT6 #(
   .INIT(64'h733f69c7733f69c7)  
) LUT6_inst8990 (
   .O(to_level3[1214]),
   .I0(level4_in[7284]),
   .I1(level4_in[7285]),
   .I2(level4_in[7286]),
   .I3(level4_in[7287]),
   .I4(level4_in[7288]),
   .I5(level4_in[7289])
);

LUT6 #(
   .INIT(64'h47d186f747d186f7)  
) LUT6_inst8991 (
   .O(to_level3[1215]),
   .I0(level4_in[7290]),
   .I1(level4_in[7291]),
   .I2(level4_in[7292]),
   .I3(level4_in[7293]),
   .I4(level4_in[7294]),
   .I5(level4_in[7295])
);

LUT6 #(
   .INIT(64'h40b1adf340b1adf3)  
) LUT6_inst8992 (
   .O(to_level3[1216]),
   .I0(level4_in[7296]),
   .I1(level4_in[7297]),
   .I2(level4_in[7298]),
   .I3(level4_in[7299]),
   .I4(level4_in[7300]),
   .I5(level4_in[7301])
);

LUT6 #(
   .INIT(64'h9966b0589966b058)  
) LUT6_inst8993 (
   .O(to_level3[1217]),
   .I0(level4_in[7302]),
   .I1(level4_in[7303]),
   .I2(level4_in[7304]),
   .I3(level4_in[7305]),
   .I4(level4_in[7306]),
   .I5(level4_in[7307])
);

LUT6 #(
   .INIT(64'hc1bd830dc1bd830d)  
) LUT6_inst8994 (
   .O(to_level3[1218]),
   .I0(level4_in[7308]),
   .I1(level4_in[7309]),
   .I2(level4_in[7310]),
   .I3(level4_in[7311]),
   .I4(level4_in[7312]),
   .I5(level4_in[7313])
);

LUT6 #(
   .INIT(64'ha4098cbea4098cbe)  
) LUT6_inst8995 (
   .O(to_level3[1219]),
   .I0(level4_in[7314]),
   .I1(level4_in[7315]),
   .I2(level4_in[7316]),
   .I3(level4_in[7317]),
   .I4(level4_in[7318]),
   .I5(level4_in[7319])
);

LUT6 #(
   .INIT(64'h67d8d71667d8d716)  
) LUT6_inst8996 (
   .O(to_level3[1220]),
   .I0(level4_in[7320]),
   .I1(level4_in[7321]),
   .I2(level4_in[7322]),
   .I3(level4_in[7323]),
   .I4(level4_in[7324]),
   .I5(level4_in[7325])
);

LUT6 #(
   .INIT(64'h9a940d4b9a940d4b)  
) LUT6_inst8997 (
   .O(to_level3[1221]),
   .I0(level4_in[7326]),
   .I1(level4_in[7327]),
   .I2(level4_in[7328]),
   .I3(level4_in[7329]),
   .I4(level4_in[7330]),
   .I5(level4_in[7331])
);

LUT6 #(
   .INIT(64'h700c0c90700c0c90)  
) LUT6_inst8998 (
   .O(to_level3[1222]),
   .I0(level4_in[7332]),
   .I1(level4_in[7333]),
   .I2(level4_in[7334]),
   .I3(level4_in[7335]),
   .I4(level4_in[7336]),
   .I5(level4_in[7337])
);

LUT6 #(
   .INIT(64'h5ca9c6155ca9c615)  
) LUT6_inst8999 (
   .O(to_level3[1223]),
   .I0(level4_in[7338]),
   .I1(level4_in[7339]),
   .I2(level4_in[7340]),
   .I3(level4_in[7341]),
   .I4(level4_in[7342]),
   .I5(level4_in[7343])
);

LUT6 #(
   .INIT(64'h165c0979165c0979)  
) LUT6_inst9000 (
   .O(to_level3[1224]),
   .I0(level4_in[7344]),
   .I1(level4_in[7345]),
   .I2(level4_in[7346]),
   .I3(level4_in[7347]),
   .I4(level4_in[7348]),
   .I5(level4_in[7349])
);

LUT6 #(
   .INIT(64'hcfd92023cfd92023)  
) LUT6_inst9001 (
   .O(to_level3[1225]),
   .I0(level4_in[7350]),
   .I1(level4_in[7351]),
   .I2(level4_in[7352]),
   .I3(level4_in[7353]),
   .I4(level4_in[7354]),
   .I5(level4_in[7355])
);

LUT6 #(
   .INIT(64'h50a5722550a57225)  
) LUT6_inst9002 (
   .O(to_level3[1226]),
   .I0(level4_in[7356]),
   .I1(level4_in[7357]),
   .I2(level4_in[7358]),
   .I3(level4_in[7359]),
   .I4(level4_in[7360]),
   .I5(level4_in[7361])
);

LUT6 #(
   .INIT(64'ha9d53997a9d53997)  
) LUT6_inst9003 (
   .O(to_level3[1227]),
   .I0(level4_in[7362]),
   .I1(level4_in[7363]),
   .I2(level4_in[7364]),
   .I3(level4_in[7365]),
   .I4(level4_in[7366]),
   .I5(level4_in[7367])
);

LUT6 #(
   .INIT(64'h4753f1b54753f1b5)  
) LUT6_inst9004 (
   .O(to_level3[1228]),
   .I0(level4_in[7368]),
   .I1(level4_in[7369]),
   .I2(level4_in[7370]),
   .I3(level4_in[7371]),
   .I4(level4_in[7372]),
   .I5(level4_in[7373])
);

LUT6 #(
   .INIT(64'he9a0f5c7e9a0f5c7)  
) LUT6_inst9005 (
   .O(to_level3[1229]),
   .I0(level4_in[7374]),
   .I1(level4_in[7375]),
   .I2(level4_in[7376]),
   .I3(level4_in[7377]),
   .I4(level4_in[7378]),
   .I5(level4_in[7379])
);

LUT6 #(
   .INIT(64'h57aef32657aef326)  
) LUT6_inst9006 (
   .O(to_level3[1230]),
   .I0(level4_in[7380]),
   .I1(level4_in[7381]),
   .I2(level4_in[7382]),
   .I3(level4_in[7383]),
   .I4(level4_in[7384]),
   .I5(level4_in[7385])
);

LUT6 #(
   .INIT(64'hd0718887d0718887)  
) LUT6_inst9007 (
   .O(to_level3[1231]),
   .I0(level4_in[7386]),
   .I1(level4_in[7387]),
   .I2(level4_in[7388]),
   .I3(level4_in[7389]),
   .I4(level4_in[7390]),
   .I5(level4_in[7391])
);

LUT6 #(
   .INIT(64'h0f922e560f922e56)  
) LUT6_inst9008 (
   .O(to_level3[1232]),
   .I0(level4_in[7392]),
   .I1(level4_in[7393]),
   .I2(level4_in[7394]),
   .I3(level4_in[7395]),
   .I4(level4_in[7396]),
   .I5(level4_in[7397])
);

LUT6 #(
   .INIT(64'h0ef40a140ef40a14)  
) LUT6_inst9009 (
   .O(to_level3[1233]),
   .I0(level4_in[7398]),
   .I1(level4_in[7399]),
   .I2(level4_in[7400]),
   .I3(level4_in[7401]),
   .I4(level4_in[7402]),
   .I5(level4_in[7403])
);

LUT6 #(
   .INIT(64'h85494e2285494e22)  
) LUT6_inst9010 (
   .O(to_level3[1234]),
   .I0(level4_in[7404]),
   .I1(level4_in[7405]),
   .I2(level4_in[7406]),
   .I3(level4_in[7407]),
   .I4(level4_in[7408]),
   .I5(level4_in[7409])
);

LUT6 #(
   .INIT(64'h8b7df84b8b7df84b)  
) LUT6_inst9011 (
   .O(to_level3[1235]),
   .I0(level4_in[7410]),
   .I1(level4_in[7411]),
   .I2(level4_in[7412]),
   .I3(level4_in[7413]),
   .I4(level4_in[7414]),
   .I5(level4_in[7415])
);

LUT6 #(
   .INIT(64'h68099ebd68099ebd)  
) LUT6_inst9012 (
   .O(to_level3[1236]),
   .I0(level4_in[7416]),
   .I1(level4_in[7417]),
   .I2(level4_in[7418]),
   .I3(level4_in[7419]),
   .I4(level4_in[7420]),
   .I5(level4_in[7421])
);

LUT6 #(
   .INIT(64'h1f0a5bc71f0a5bc7)  
) LUT6_inst9013 (
   .O(to_level3[1237]),
   .I0(level4_in[7422]),
   .I1(level4_in[7423]),
   .I2(level4_in[7424]),
   .I3(level4_in[7425]),
   .I4(level4_in[7426]),
   .I5(level4_in[7427])
);

LUT6 #(
   .INIT(64'h2267d26c2267d26c)  
) LUT6_inst9014 (
   .O(to_level3[1238]),
   .I0(level4_in[7428]),
   .I1(level4_in[7429]),
   .I2(level4_in[7430]),
   .I3(level4_in[7431]),
   .I4(level4_in[7432]),
   .I5(level4_in[7433])
);

LUT6 #(
   .INIT(64'h4e65910b4e65910b)  
) LUT6_inst9015 (
   .O(to_level3[1239]),
   .I0(level4_in[7434]),
   .I1(level4_in[7435]),
   .I2(level4_in[7436]),
   .I3(level4_in[7437]),
   .I4(level4_in[7438]),
   .I5(level4_in[7439])
);

LUT6 #(
   .INIT(64'hd646211fd646211f)  
) LUT6_inst9016 (
   .O(to_level3[1240]),
   .I0(level4_in[7440]),
   .I1(level4_in[7441]),
   .I2(level4_in[7442]),
   .I3(level4_in[7443]),
   .I4(level4_in[7444]),
   .I5(level4_in[7445])
);

LUT6 #(
   .INIT(64'h6285c7886285c788)  
) LUT6_inst9017 (
   .O(to_level3[1241]),
   .I0(level4_in[7446]),
   .I1(level4_in[7447]),
   .I2(level4_in[7448]),
   .I3(level4_in[7449]),
   .I4(level4_in[7450]),
   .I5(level4_in[7451])
);

LUT6 #(
   .INIT(64'had22a03bad22a03b)  
) LUT6_inst9018 (
   .O(to_level3[1242]),
   .I0(level4_in[7452]),
   .I1(level4_in[7453]),
   .I2(level4_in[7454]),
   .I3(level4_in[7455]),
   .I4(level4_in[7456]),
   .I5(level4_in[7457])
);

LUT6 #(
   .INIT(64'hf631f7e8f631f7e8)  
) LUT6_inst9019 (
   .O(to_level3[1243]),
   .I0(level4_in[7458]),
   .I1(level4_in[7459]),
   .I2(level4_in[7460]),
   .I3(level4_in[7461]),
   .I4(level4_in[7462]),
   .I5(level4_in[7463])
);

LUT6 #(
   .INIT(64'hc72339d5c72339d5)  
) LUT6_inst9020 (
   .O(to_level3[1244]),
   .I0(level4_in[7464]),
   .I1(level4_in[7465]),
   .I2(level4_in[7466]),
   .I3(level4_in[7467]),
   .I4(level4_in[7468]),
   .I5(level4_in[7469])
);

LUT6 #(
   .INIT(64'h6b94dced6b94dced)  
) LUT6_inst9021 (
   .O(to_level3[1245]),
   .I0(level4_in[7470]),
   .I1(level4_in[7471]),
   .I2(level4_in[7472]),
   .I3(level4_in[7473]),
   .I4(level4_in[7474]),
   .I5(level4_in[7475])
);

LUT6 #(
   .INIT(64'h901298cc901298cc)  
) LUT6_inst9022 (
   .O(to_level3[1246]),
   .I0(level4_in[7476]),
   .I1(level4_in[7477]),
   .I2(level4_in[7478]),
   .I3(level4_in[7479]),
   .I4(level4_in[7480]),
   .I5(level4_in[7481])
);

LUT6 #(
   .INIT(64'h972851d4972851d4)  
) LUT6_inst9023 (
   .O(to_level3[1247]),
   .I0(level4_in[7482]),
   .I1(level4_in[7483]),
   .I2(level4_in[7484]),
   .I3(level4_in[7485]),
   .I4(level4_in[7486]),
   .I5(level4_in[7487])
);

LUT6 #(
   .INIT(64'hd0e7c4e0d0e7c4e0)  
) LUT6_inst9024 (
   .O(to_level3[1248]),
   .I0(level4_in[7488]),
   .I1(level4_in[7489]),
   .I2(level4_in[7490]),
   .I3(level4_in[7491]),
   .I4(level4_in[7492]),
   .I5(level4_in[7493])
);

LUT6 #(
   .INIT(64'h90c1886590c18865)  
) LUT6_inst9025 (
   .O(to_level3[1249]),
   .I0(level4_in[7494]),
   .I1(level4_in[7495]),
   .I2(level4_in[7496]),
   .I3(level4_in[7497]),
   .I4(level4_in[7498]),
   .I5(level4_in[7499])
);

LUT6 #(
   .INIT(64'hbc4cfa1fbc4cfa1f)  
) LUT6_inst9026 (
   .O(to_level3[1250]),
   .I0(level4_in[7500]),
   .I1(level4_in[7501]),
   .I2(level4_in[7502]),
   .I3(level4_in[7503]),
   .I4(level4_in[7504]),
   .I5(level4_in[7505])
);

LUT6 #(
   .INIT(64'h31eab6d831eab6d8)  
) LUT6_inst9027 (
   .O(to_level3[1251]),
   .I0(level4_in[7506]),
   .I1(level4_in[7507]),
   .I2(level4_in[7508]),
   .I3(level4_in[7509]),
   .I4(level4_in[7510]),
   .I5(level4_in[7511])
);

LUT6 #(
   .INIT(64'hdd43a560dd43a560)  
) LUT6_inst9028 (
   .O(to_level3[1252]),
   .I0(level4_in[7512]),
   .I1(level4_in[7513]),
   .I2(level4_in[7514]),
   .I3(level4_in[7515]),
   .I4(level4_in[7516]),
   .I5(level4_in[7517])
);

LUT6 #(
   .INIT(64'hb5e6ab52b5e6ab52)  
) LUT6_inst9029 (
   .O(to_level3[1253]),
   .I0(level4_in[7518]),
   .I1(level4_in[7519]),
   .I2(level4_in[7520]),
   .I3(level4_in[7521]),
   .I4(level4_in[7522]),
   .I5(level4_in[7523])
);

LUT6 #(
   .INIT(64'hcb01e93acb01e93a)  
) LUT6_inst9030 (
   .O(to_level3[1254]),
   .I0(level4_in[7524]),
   .I1(level4_in[7525]),
   .I2(level4_in[7526]),
   .I3(level4_in[7527]),
   .I4(level4_in[7528]),
   .I5(level4_in[7529])
);

LUT6 #(
   .INIT(64'h37b5aebf37b5aebf)  
) LUT6_inst9031 (
   .O(to_level3[1255]),
   .I0(level4_in[7530]),
   .I1(level4_in[7531]),
   .I2(level4_in[7532]),
   .I3(level4_in[7533]),
   .I4(level4_in[7534]),
   .I5(level4_in[7535])
);

LUT6 #(
   .INIT(64'hc6573e4fc6573e4f)  
) LUT6_inst9032 (
   .O(to_level3[1256]),
   .I0(level4_in[7536]),
   .I1(level4_in[7537]),
   .I2(level4_in[7538]),
   .I3(level4_in[7539]),
   .I4(level4_in[7540]),
   .I5(level4_in[7541])
);

LUT6 #(
   .INIT(64'h9456a50a9456a50a)  
) LUT6_inst9033 (
   .O(to_level3[1257]),
   .I0(level4_in[7542]),
   .I1(level4_in[7543]),
   .I2(level4_in[7544]),
   .I3(level4_in[7545]),
   .I4(level4_in[7546]),
   .I5(level4_in[7547])
);

LUT6 #(
   .INIT(64'hf03ef7f6f03ef7f6)  
) LUT6_inst9034 (
   .O(to_level3[1258]),
   .I0(level4_in[7548]),
   .I1(level4_in[7549]),
   .I2(level4_in[7550]),
   .I3(level4_in[7551]),
   .I4(level4_in[7552]),
   .I5(level4_in[7553])
);

LUT6 #(
   .INIT(64'hf9f56139f9f56139)  
) LUT6_inst9035 (
   .O(to_level3[1259]),
   .I0(level4_in[7554]),
   .I1(level4_in[7555]),
   .I2(level4_in[7556]),
   .I3(level4_in[7557]),
   .I4(level4_in[7558]),
   .I5(level4_in[7559])
);

LUT6 #(
   .INIT(64'hb89f6f46b89f6f46)  
) LUT6_inst9036 (
   .O(to_level3[1260]),
   .I0(level4_in[7560]),
   .I1(level4_in[7561]),
   .I2(level4_in[7562]),
   .I3(level4_in[7563]),
   .I4(level4_in[7564]),
   .I5(level4_in[7565])
);

LUT6 #(
   .INIT(64'h5fd386a85fd386a8)  
) LUT6_inst9037 (
   .O(to_level3[1261]),
   .I0(level4_in[7566]),
   .I1(level4_in[7567]),
   .I2(level4_in[7568]),
   .I3(level4_in[7569]),
   .I4(level4_in[7570]),
   .I5(level4_in[7571])
);

LUT6 #(
   .INIT(64'h65feb52165feb521)  
) LUT6_inst9038 (
   .O(to_level3[1262]),
   .I0(level4_in[7572]),
   .I1(level4_in[7573]),
   .I2(level4_in[7574]),
   .I3(level4_in[7575]),
   .I4(level4_in[7576]),
   .I5(level4_in[7577])
);

LUT6 #(
   .INIT(64'h1fa0d7fe1fa0d7fe)  
) LUT6_inst9039 (
   .O(to_level3[1263]),
   .I0(level4_in[7578]),
   .I1(level4_in[7579]),
   .I2(level4_in[7580]),
   .I3(level4_in[7581]),
   .I4(level4_in[7582]),
   .I5(level4_in[7583])
);

LUT6 #(
   .INIT(64'hecf40e48ecf40e48)  
) LUT6_inst9040 (
   .O(to_level3[1264]),
   .I0(level4_in[7584]),
   .I1(level4_in[7585]),
   .I2(level4_in[7586]),
   .I3(level4_in[7587]),
   .I4(level4_in[7588]),
   .I5(level4_in[7589])
);

LUT6 #(
   .INIT(64'h01892f4c01892f4c)  
) LUT6_inst9041 (
   .O(to_level3[1265]),
   .I0(level4_in[7590]),
   .I1(level4_in[7591]),
   .I2(level4_in[7592]),
   .I3(level4_in[7593]),
   .I4(level4_in[7594]),
   .I5(level4_in[7595])
);

LUT6 #(
   .INIT(64'h7df7067d7df7067d)  
) LUT6_inst9042 (
   .O(to_level3[1266]),
   .I0(level4_in[7596]),
   .I1(level4_in[7597]),
   .I2(level4_in[7598]),
   .I3(level4_in[7599]),
   .I4(level4_in[7600]),
   .I5(level4_in[7601])
);

LUT6 #(
   .INIT(64'h662b9a75662b9a75)  
) LUT6_inst9043 (
   .O(to_level3[1267]),
   .I0(level4_in[7602]),
   .I1(level4_in[7603]),
   .I2(level4_in[7604]),
   .I3(level4_in[7605]),
   .I4(level4_in[7606]),
   .I5(level4_in[7607])
);

LUT6 #(
   .INIT(64'hd0c96bc8d0c96bc8)  
) LUT6_inst9044 (
   .O(to_level3[1268]),
   .I0(level4_in[7608]),
   .I1(level4_in[7609]),
   .I2(level4_in[7610]),
   .I3(level4_in[7611]),
   .I4(level4_in[7612]),
   .I5(level4_in[7613])
);

LUT6 #(
   .INIT(64'h1ff3c1091ff3c109)  
) LUT6_inst9045 (
   .O(to_level3[1269]),
   .I0(level4_in[7614]),
   .I1(level4_in[7615]),
   .I2(level4_in[7616]),
   .I3(level4_in[7617]),
   .I4(level4_in[7618]),
   .I5(level4_in[7619])
);

LUT6 #(
   .INIT(64'h963c9f83963c9f83)  
) LUT6_inst9046 (
   .O(to_level3[1270]),
   .I0(level4_in[7620]),
   .I1(level4_in[7621]),
   .I2(level4_in[7622]),
   .I3(level4_in[7623]),
   .I4(level4_in[7624]),
   .I5(level4_in[7625])
);

LUT6 #(
   .INIT(64'hc935d34ec935d34e)  
) LUT6_inst9047 (
   .O(to_level3[1271]),
   .I0(level4_in[7626]),
   .I1(level4_in[7627]),
   .I2(level4_in[7628]),
   .I3(level4_in[7629]),
   .I4(level4_in[7630]),
   .I5(level4_in[7631])
);

LUT6 #(
   .INIT(64'h0cb18b610cb18b61)  
) LUT6_inst9048 (
   .O(to_level3[1272]),
   .I0(level4_in[7632]),
   .I1(level4_in[7633]),
   .I2(level4_in[7634]),
   .I3(level4_in[7635]),
   .I4(level4_in[7636]),
   .I5(level4_in[7637])
);

LUT6 #(
   .INIT(64'hf5178ea9f5178ea9)  
) LUT6_inst9049 (
   .O(to_level3[1273]),
   .I0(level4_in[7638]),
   .I1(level4_in[7639]),
   .I2(level4_in[7640]),
   .I3(level4_in[7641]),
   .I4(level4_in[7642]),
   .I5(level4_in[7643])
);

LUT6 #(
   .INIT(64'h721dd3cd721dd3cd)  
) LUT6_inst9050 (
   .O(to_level3[1274]),
   .I0(level4_in[7644]),
   .I1(level4_in[7645]),
   .I2(level4_in[7646]),
   .I3(level4_in[7647]),
   .I4(level4_in[7648]),
   .I5(level4_in[7649])
);

LUT6 #(
   .INIT(64'h36eb6caa36eb6caa)  
) LUT6_inst9051 (
   .O(to_level3[1275]),
   .I0(level4_in[7650]),
   .I1(level4_in[7651]),
   .I2(level4_in[7652]),
   .I3(level4_in[7653]),
   .I4(level4_in[7654]),
   .I5(level4_in[7655])
);

LUT6 #(
   .INIT(64'h33f903af33f903af)  
) LUT6_inst9052 (
   .O(to_level3[1276]),
   .I0(level4_in[7656]),
   .I1(level4_in[7657]),
   .I2(level4_in[7658]),
   .I3(level4_in[7659]),
   .I4(level4_in[7660]),
   .I5(level4_in[7661])
);

LUT6 #(
   .INIT(64'h4738090747380907)  
) LUT6_inst9053 (
   .O(to_level3[1277]),
   .I0(level4_in[7662]),
   .I1(level4_in[7663]),
   .I2(level4_in[7664]),
   .I3(level4_in[7665]),
   .I4(level4_in[7666]),
   .I5(level4_in[7667])
);

LUT6 #(
   .INIT(64'he086a7cbe086a7cb)  
) LUT6_inst9054 (
   .O(to_level3[1278]),
   .I0(level4_in[7668]),
   .I1(level4_in[7669]),
   .I2(level4_in[7670]),
   .I3(level4_in[7671]),
   .I4(level4_in[7672]),
   .I5(level4_in[7673])
);

LUT6 #(
   .INIT(64'h17d6e0e217d6e0e2)  
) LUT6_inst9055 (
   .O(to_level3[1279]),
   .I0(level4_in[7674]),
   .I1(level4_in[7675]),
   .I2(level4_in[7676]),
   .I3(level4_in[7677]),
   .I4(level4_in[7678]),
   .I5(level4_in[7679])
);

LUT6 #(
   .INIT(64'h5cfb47d65cfb47d6)  
) LUT6_inst9056 (
   .O(to_level3[1280]),
   .I0(level4_in[7680]),
   .I1(level4_in[7681]),
   .I2(level4_in[7682]),
   .I3(level4_in[7683]),
   .I4(level4_in[7684]),
   .I5(level4_in[7685])
);

LUT6 #(
   .INIT(64'hf216c4d7f216c4d7)  
) LUT6_inst9057 (
   .O(to_level3[1281]),
   .I0(level4_in[7686]),
   .I1(level4_in[7687]),
   .I2(level4_in[7688]),
   .I3(level4_in[7689]),
   .I4(level4_in[7690]),
   .I5(level4_in[7691])
);

LUT6 #(
   .INIT(64'he3afbfb3e3afbfb3)  
) LUT6_inst9058 (
   .O(to_level3[1282]),
   .I0(level4_in[7692]),
   .I1(level4_in[7693]),
   .I2(level4_in[7694]),
   .I3(level4_in[7695]),
   .I4(level4_in[7696]),
   .I5(level4_in[7697])
);

LUT6 #(
   .INIT(64'hbdfc8921bdfc8921)  
) LUT6_inst9059 (
   .O(to_level3[1283]),
   .I0(level4_in[7698]),
   .I1(level4_in[7699]),
   .I2(level4_in[7700]),
   .I3(level4_in[7701]),
   .I4(level4_in[7702]),
   .I5(level4_in[7703])
);

LUT6 #(
   .INIT(64'h79cf3c4c79cf3c4c)  
) LUT6_inst9060 (
   .O(to_level3[1284]),
   .I0(level4_in[7704]),
   .I1(level4_in[7705]),
   .I2(level4_in[7706]),
   .I3(level4_in[7707]),
   .I4(level4_in[7708]),
   .I5(level4_in[7709])
);

LUT6 #(
   .INIT(64'hde0ca2cdde0ca2cd)  
) LUT6_inst9061 (
   .O(to_level3[1285]),
   .I0(level4_in[7710]),
   .I1(level4_in[7711]),
   .I2(level4_in[7712]),
   .I3(level4_in[7713]),
   .I4(level4_in[7714]),
   .I5(level4_in[7715])
);

LUT6 #(
   .INIT(64'h9b2d52dd9b2d52dd)  
) LUT6_inst9062 (
   .O(to_level3[1286]),
   .I0(level4_in[7716]),
   .I1(level4_in[7717]),
   .I2(level4_in[7718]),
   .I3(level4_in[7719]),
   .I4(level4_in[7720]),
   .I5(level4_in[7721])
);

LUT6 #(
   .INIT(64'h94af059894af0598)  
) LUT6_inst9063 (
   .O(to_level3[1287]),
   .I0(level4_in[7722]),
   .I1(level4_in[7723]),
   .I2(level4_in[7724]),
   .I3(level4_in[7725]),
   .I4(level4_in[7726]),
   .I5(level4_in[7727])
);

LUT6 #(
   .INIT(64'hb4b8781cb4b8781c)  
) LUT6_inst9064 (
   .O(to_level3[1288]),
   .I0(level4_in[7728]),
   .I1(level4_in[7729]),
   .I2(level4_in[7730]),
   .I3(level4_in[7731]),
   .I4(level4_in[7732]),
   .I5(level4_in[7733])
);

LUT6 #(
   .INIT(64'h1663586416635864)  
) LUT6_inst9065 (
   .O(to_level3[1289]),
   .I0(level4_in[7734]),
   .I1(level4_in[7735]),
   .I2(level4_in[7736]),
   .I3(level4_in[7737]),
   .I4(level4_in[7738]),
   .I5(level4_in[7739])
);

LUT6 #(
   .INIT(64'h3e1384573e138457)  
) LUT6_inst9066 (
   .O(to_level3[1290]),
   .I0(level4_in[7740]),
   .I1(level4_in[7741]),
   .I2(level4_in[7742]),
   .I3(level4_in[7743]),
   .I4(level4_in[7744]),
   .I5(level4_in[7745])
);

LUT6 #(
   .INIT(64'h7ccefd1a7ccefd1a)  
) LUT6_inst9067 (
   .O(to_level3[1291]),
   .I0(level4_in[7746]),
   .I1(level4_in[7747]),
   .I2(level4_in[7748]),
   .I3(level4_in[7749]),
   .I4(level4_in[7750]),
   .I5(level4_in[7751])
);

LUT6 #(
   .INIT(64'h7174516771745167)  
) LUT6_inst9068 (
   .O(to_level3[1292]),
   .I0(level4_in[7752]),
   .I1(level4_in[7753]),
   .I2(level4_in[7754]),
   .I3(level4_in[7755]),
   .I4(level4_in[7756]),
   .I5(level4_in[7757])
);

LUT6 #(
   .INIT(64'hf45f3a0bf45f3a0b)  
) LUT6_inst9069 (
   .O(to_level3[1293]),
   .I0(level4_in[7758]),
   .I1(level4_in[7759]),
   .I2(level4_in[7760]),
   .I3(level4_in[7761]),
   .I4(level4_in[7762]),
   .I5(level4_in[7763])
);

LUT6 #(
   .INIT(64'h3aeddc233aeddc23)  
) LUT6_inst9070 (
   .O(to_level3[1294]),
   .I0(level4_in[7764]),
   .I1(level4_in[7765]),
   .I2(level4_in[7766]),
   .I3(level4_in[7767]),
   .I4(level4_in[7768]),
   .I5(level4_in[7769])
);

LUT6 #(
   .INIT(64'h215480a2215480a2)  
) LUT6_inst9071 (
   .O(to_level3[1295]),
   .I0(level4_in[7770]),
   .I1(level4_in[7771]),
   .I2(level4_in[7772]),
   .I3(level4_in[7773]),
   .I4(level4_in[7774]),
   .I5(level4_in[7775])
);
////////////// level 3 starts below:/n
LUT6 #(
   .INIT(64'h5942de315942de31)  
) LUT6_inst9072 (
   .O(to_level2[0]),
   .I0(level3_in[0]),
   .I1(level3_in[1]),
   .I2(level3_in[2]),
   .I3(level3_in[3]),
   .I4(level3_in[4]),
   .I5(level3_in[5])
);

LUT6 #(
   .INIT(64'hf5334c15f5334c15)  
) LUT6_inst9073 (
   .O(to_level2[1]),
   .I0(level3_in[6]),
   .I1(level3_in[7]),
   .I2(level3_in[8]),
   .I3(level3_in[9]),
   .I4(level3_in[10]),
   .I5(level3_in[11])
);

LUT6 #(
   .INIT(64'h3787825737878257)  
) LUT6_inst9074 (
   .O(to_level2[2]),
   .I0(level3_in[12]),
   .I1(level3_in[13]),
   .I2(level3_in[14]),
   .I3(level3_in[15]),
   .I4(level3_in[16]),
   .I5(level3_in[17])
);

LUT6 #(
   .INIT(64'hb7186afcb7186afc)  
) LUT6_inst9075 (
   .O(to_level2[3]),
   .I0(level3_in[18]),
   .I1(level3_in[19]),
   .I2(level3_in[20]),
   .I3(level3_in[21]),
   .I4(level3_in[22]),
   .I5(level3_in[23])
);

LUT6 #(
   .INIT(64'hd2a87662d2a87662)  
) LUT6_inst9076 (
   .O(to_level2[4]),
   .I0(level3_in[24]),
   .I1(level3_in[25]),
   .I2(level3_in[26]),
   .I3(level3_in[27]),
   .I4(level3_in[28]),
   .I5(level3_in[29])
);

LUT6 #(
   .INIT(64'h91cc14cb91cc14cb)  
) LUT6_inst9077 (
   .O(to_level2[5]),
   .I0(level3_in[30]),
   .I1(level3_in[31]),
   .I2(level3_in[32]),
   .I3(level3_in[33]),
   .I4(level3_in[34]),
   .I5(level3_in[35])
);

LUT6 #(
   .INIT(64'hf5279db0f5279db0)  
) LUT6_inst9078 (
   .O(to_level2[6]),
   .I0(level3_in[36]),
   .I1(level3_in[37]),
   .I2(level3_in[38]),
   .I3(level3_in[39]),
   .I4(level3_in[40]),
   .I5(level3_in[41])
);

LUT6 #(
   .INIT(64'h59e029cc59e029cc)  
) LUT6_inst9079 (
   .O(to_level2[7]),
   .I0(level3_in[42]),
   .I1(level3_in[43]),
   .I2(level3_in[44]),
   .I3(level3_in[45]),
   .I4(level3_in[46]),
   .I5(level3_in[47])
);

LUT6 #(
   .INIT(64'hf69e70d8f69e70d8)  
) LUT6_inst9080 (
   .O(to_level2[8]),
   .I0(level3_in[48]),
   .I1(level3_in[49]),
   .I2(level3_in[50]),
   .I3(level3_in[51]),
   .I4(level3_in[52]),
   .I5(level3_in[53])
);

LUT6 #(
   .INIT(64'haa35084aaa35084a)  
) LUT6_inst9081 (
   .O(to_level2[9]),
   .I0(level3_in[54]),
   .I1(level3_in[55]),
   .I2(level3_in[56]),
   .I3(level3_in[57]),
   .I4(level3_in[58]),
   .I5(level3_in[59])
);

LUT6 #(
   .INIT(64'h5c6185fb5c6185fb)  
) LUT6_inst9082 (
   .O(to_level2[10]),
   .I0(level3_in[60]),
   .I1(level3_in[61]),
   .I2(level3_in[62]),
   .I3(level3_in[63]),
   .I4(level3_in[64]),
   .I5(level3_in[65])
);

LUT6 #(
   .INIT(64'h3d5aebb83d5aebb8)  
) LUT6_inst9083 (
   .O(to_level2[11]),
   .I0(level3_in[66]),
   .I1(level3_in[67]),
   .I2(level3_in[68]),
   .I3(level3_in[69]),
   .I4(level3_in[70]),
   .I5(level3_in[71])
);

LUT6 #(
   .INIT(64'h9b84e6169b84e616)  
) LUT6_inst9084 (
   .O(to_level2[12]),
   .I0(level3_in[72]),
   .I1(level3_in[73]),
   .I2(level3_in[74]),
   .I3(level3_in[75]),
   .I4(level3_in[76]),
   .I5(level3_in[77])
);

LUT6 #(
   .INIT(64'hf724fea1f724fea1)  
) LUT6_inst9085 (
   .O(to_level2[13]),
   .I0(level3_in[78]),
   .I1(level3_in[79]),
   .I2(level3_in[80]),
   .I3(level3_in[81]),
   .I4(level3_in[82]),
   .I5(level3_in[83])
);

LUT6 #(
   .INIT(64'h7d86a1ee7d86a1ee)  
) LUT6_inst9086 (
   .O(to_level2[14]),
   .I0(level3_in[84]),
   .I1(level3_in[85]),
   .I2(level3_in[86]),
   .I3(level3_in[87]),
   .I4(level3_in[88]),
   .I5(level3_in[89])
);

LUT6 #(
   .INIT(64'hff066e3bff066e3b)  
) LUT6_inst9087 (
   .O(to_level2[15]),
   .I0(level3_in[90]),
   .I1(level3_in[91]),
   .I2(level3_in[92]),
   .I3(level3_in[93]),
   .I4(level3_in[94]),
   .I5(level3_in[95])
);

LUT6 #(
   .INIT(64'hfe192fe0fe192fe0)  
) LUT6_inst9088 (
   .O(to_level2[16]),
   .I0(level3_in[96]),
   .I1(level3_in[97]),
   .I2(level3_in[98]),
   .I3(level3_in[99]),
   .I4(level3_in[100]),
   .I5(level3_in[101])
);

LUT6 #(
   .INIT(64'hbaad9de7baad9de7)  
) LUT6_inst9089 (
   .O(to_level2[17]),
   .I0(level3_in[102]),
   .I1(level3_in[103]),
   .I2(level3_in[104]),
   .I3(level3_in[105]),
   .I4(level3_in[106]),
   .I5(level3_in[107])
);

LUT6 #(
   .INIT(64'h82e1dce282e1dce2)  
) LUT6_inst9090 (
   .O(to_level2[18]),
   .I0(level3_in[108]),
   .I1(level3_in[109]),
   .I2(level3_in[110]),
   .I3(level3_in[111]),
   .I4(level3_in[112]),
   .I5(level3_in[113])
);

LUT6 #(
   .INIT(64'h244b21d5244b21d5)  
) LUT6_inst9091 (
   .O(to_level2[19]),
   .I0(level3_in[114]),
   .I1(level3_in[115]),
   .I2(level3_in[116]),
   .I3(level3_in[117]),
   .I4(level3_in[118]),
   .I5(level3_in[119])
);

LUT6 #(
   .INIT(64'h34a885c234a885c2)  
) LUT6_inst9092 (
   .O(to_level2[20]),
   .I0(level3_in[120]),
   .I1(level3_in[121]),
   .I2(level3_in[122]),
   .I3(level3_in[123]),
   .I4(level3_in[124]),
   .I5(level3_in[125])
);

LUT6 #(
   .INIT(64'h0c001ce50c001ce5)  
) LUT6_inst9093 (
   .O(to_level2[21]),
   .I0(level3_in[126]),
   .I1(level3_in[127]),
   .I2(level3_in[128]),
   .I3(level3_in[129]),
   .I4(level3_in[130]),
   .I5(level3_in[131])
);

LUT6 #(
   .INIT(64'hec6c9fa2ec6c9fa2)  
) LUT6_inst9094 (
   .O(to_level2[22]),
   .I0(level3_in[132]),
   .I1(level3_in[133]),
   .I2(level3_in[134]),
   .I3(level3_in[135]),
   .I4(level3_in[136]),
   .I5(level3_in[137])
);

LUT6 #(
   .INIT(64'h9bb125ca9bb125ca)  
) LUT6_inst9095 (
   .O(to_level2[23]),
   .I0(level3_in[138]),
   .I1(level3_in[139]),
   .I2(level3_in[140]),
   .I3(level3_in[141]),
   .I4(level3_in[142]),
   .I5(level3_in[143])
);

LUT6 #(
   .INIT(64'hfba8f21cfba8f21c)  
) LUT6_inst9096 (
   .O(to_level2[24]),
   .I0(level3_in[144]),
   .I1(level3_in[145]),
   .I2(level3_in[146]),
   .I3(level3_in[147]),
   .I4(level3_in[148]),
   .I5(level3_in[149])
);

LUT6 #(
   .INIT(64'h4029735a4029735a)  
) LUT6_inst9097 (
   .O(to_level2[25]),
   .I0(level3_in[150]),
   .I1(level3_in[151]),
   .I2(level3_in[152]),
   .I3(level3_in[153]),
   .I4(level3_in[154]),
   .I5(level3_in[155])
);

LUT6 #(
   .INIT(64'h156c3351156c3351)  
) LUT6_inst9098 (
   .O(to_level2[26]),
   .I0(level3_in[156]),
   .I1(level3_in[157]),
   .I2(level3_in[158]),
   .I3(level3_in[159]),
   .I4(level3_in[160]),
   .I5(level3_in[161])
);

LUT6 #(
   .INIT(64'h3b5a29643b5a2964)  
) LUT6_inst9099 (
   .O(to_level2[27]),
   .I0(level3_in[162]),
   .I1(level3_in[163]),
   .I2(level3_in[164]),
   .I3(level3_in[165]),
   .I4(level3_in[166]),
   .I5(level3_in[167])
);

LUT6 #(
   .INIT(64'hcb3cef32cb3cef32)  
) LUT6_inst9100 (
   .O(to_level2[28]),
   .I0(level3_in[168]),
   .I1(level3_in[169]),
   .I2(level3_in[170]),
   .I3(level3_in[171]),
   .I4(level3_in[172]),
   .I5(level3_in[173])
);

LUT6 #(
   .INIT(64'hf1513b0af1513b0a)  
) LUT6_inst9101 (
   .O(to_level2[29]),
   .I0(level3_in[174]),
   .I1(level3_in[175]),
   .I2(level3_in[176]),
   .I3(level3_in[177]),
   .I4(level3_in[178]),
   .I5(level3_in[179])
);

LUT6 #(
   .INIT(64'hd2948466d2948466)  
) LUT6_inst9102 (
   .O(to_level2[30]),
   .I0(level3_in[180]),
   .I1(level3_in[181]),
   .I2(level3_in[182]),
   .I3(level3_in[183]),
   .I4(level3_in[184]),
   .I5(level3_in[185])
);

LUT6 #(
   .INIT(64'h21969ebe21969ebe)  
) LUT6_inst9103 (
   .O(to_level2[31]),
   .I0(level3_in[186]),
   .I1(level3_in[187]),
   .I2(level3_in[188]),
   .I3(level3_in[189]),
   .I4(level3_in[190]),
   .I5(level3_in[191])
);

LUT6 #(
   .INIT(64'h52b6986a52b6986a)  
) LUT6_inst9104 (
   .O(to_level2[32]),
   .I0(level3_in[192]),
   .I1(level3_in[193]),
   .I2(level3_in[194]),
   .I3(level3_in[195]),
   .I4(level3_in[196]),
   .I5(level3_in[197])
);

LUT6 #(
   .INIT(64'hd21e9c7ad21e9c7a)  
) LUT6_inst9105 (
   .O(to_level2[33]),
   .I0(level3_in[198]),
   .I1(level3_in[199]),
   .I2(level3_in[200]),
   .I3(level3_in[201]),
   .I4(level3_in[202]),
   .I5(level3_in[203])
);

LUT6 #(
   .INIT(64'hfc020bfafc020bfa)  
) LUT6_inst9106 (
   .O(to_level2[34]),
   .I0(level3_in[204]),
   .I1(level3_in[205]),
   .I2(level3_in[206]),
   .I3(level3_in[207]),
   .I4(level3_in[208]),
   .I5(level3_in[209])
);

LUT6 #(
   .INIT(64'ha65f94dba65f94db)  
) LUT6_inst9107 (
   .O(to_level2[35]),
   .I0(level3_in[210]),
   .I1(level3_in[211]),
   .I2(level3_in[212]),
   .I3(level3_in[213]),
   .I4(level3_in[214]),
   .I5(level3_in[215])
);

LUT6 #(
   .INIT(64'hb8f1e8c4b8f1e8c4)  
) LUT6_inst9108 (
   .O(to_level2[36]),
   .I0(level3_in[216]),
   .I1(level3_in[217]),
   .I2(level3_in[218]),
   .I3(level3_in[219]),
   .I4(level3_in[220]),
   .I5(level3_in[221])
);

LUT6 #(
   .INIT(64'hbf818f29bf818f29)  
) LUT6_inst9109 (
   .O(to_level2[37]),
   .I0(level3_in[222]),
   .I1(level3_in[223]),
   .I2(level3_in[224]),
   .I3(level3_in[225]),
   .I4(level3_in[226]),
   .I5(level3_in[227])
);

LUT6 #(
   .INIT(64'h7940e51c7940e51c)  
) LUT6_inst9110 (
   .O(to_level2[38]),
   .I0(level3_in[228]),
   .I1(level3_in[229]),
   .I2(level3_in[230]),
   .I3(level3_in[231]),
   .I4(level3_in[232]),
   .I5(level3_in[233])
);

LUT6 #(
   .INIT(64'h1acfceb11acfceb1)  
) LUT6_inst9111 (
   .O(to_level2[39]),
   .I0(level3_in[234]),
   .I1(level3_in[235]),
   .I2(level3_in[236]),
   .I3(level3_in[237]),
   .I4(level3_in[238]),
   .I5(level3_in[239])
);

LUT6 #(
   .INIT(64'hdd284a7fdd284a7f)  
) LUT6_inst9112 (
   .O(to_level2[40]),
   .I0(level3_in[240]),
   .I1(level3_in[241]),
   .I2(level3_in[242]),
   .I3(level3_in[243]),
   .I4(level3_in[244]),
   .I5(level3_in[245])
);

LUT6 #(
   .INIT(64'h9c197f959c197f95)  
) LUT6_inst9113 (
   .O(to_level2[41]),
   .I0(level3_in[246]),
   .I1(level3_in[247]),
   .I2(level3_in[248]),
   .I3(level3_in[249]),
   .I4(level3_in[250]),
   .I5(level3_in[251])
);

LUT6 #(
   .INIT(64'h8447fde18447fde1)  
) LUT6_inst9114 (
   .O(to_level2[42]),
   .I0(level3_in[252]),
   .I1(level3_in[253]),
   .I2(level3_in[254]),
   .I3(level3_in[255]),
   .I4(level3_in[256]),
   .I5(level3_in[257])
);

LUT6 #(
   .INIT(64'h169a8d2c169a8d2c)  
) LUT6_inst9115 (
   .O(to_level2[43]),
   .I0(level3_in[258]),
   .I1(level3_in[259]),
   .I2(level3_in[260]),
   .I3(level3_in[261]),
   .I4(level3_in[262]),
   .I5(level3_in[263])
);

LUT6 #(
   .INIT(64'h1affeb421affeb42)  
) LUT6_inst9116 (
   .O(to_level2[44]),
   .I0(level3_in[264]),
   .I1(level3_in[265]),
   .I2(level3_in[266]),
   .I3(level3_in[267]),
   .I4(level3_in[268]),
   .I5(level3_in[269])
);

LUT6 #(
   .INIT(64'h95a1c60495a1c604)  
) LUT6_inst9117 (
   .O(to_level2[45]),
   .I0(level3_in[270]),
   .I1(level3_in[271]),
   .I2(level3_in[272]),
   .I3(level3_in[273]),
   .I4(level3_in[274]),
   .I5(level3_in[275])
);

LUT6 #(
   .INIT(64'h624bc030624bc030)  
) LUT6_inst9118 (
   .O(to_level2[46]),
   .I0(level3_in[276]),
   .I1(level3_in[277]),
   .I2(level3_in[278]),
   .I3(level3_in[279]),
   .I4(level3_in[280]),
   .I5(level3_in[281])
);

LUT6 #(
   .INIT(64'h59d0f50959d0f509)  
) LUT6_inst9119 (
   .O(to_level2[47]),
   .I0(level3_in[282]),
   .I1(level3_in[283]),
   .I2(level3_in[284]),
   .I3(level3_in[285]),
   .I4(level3_in[286]),
   .I5(level3_in[287])
);

LUT6 #(
   .INIT(64'hbf5a9748bf5a9748)  
) LUT6_inst9120 (
   .O(to_level2[48]),
   .I0(level3_in[288]),
   .I1(level3_in[289]),
   .I2(level3_in[290]),
   .I3(level3_in[291]),
   .I4(level3_in[292]),
   .I5(level3_in[293])
);

LUT6 #(
   .INIT(64'h00612eaf00612eaf)  
) LUT6_inst9121 (
   .O(to_level2[49]),
   .I0(level3_in[294]),
   .I1(level3_in[295]),
   .I2(level3_in[296]),
   .I3(level3_in[297]),
   .I4(level3_in[298]),
   .I5(level3_in[299])
);

LUT6 #(
   .INIT(64'ha02c7be6a02c7be6)  
) LUT6_inst9122 (
   .O(to_level2[50]),
   .I0(level3_in[300]),
   .I1(level3_in[301]),
   .I2(level3_in[302]),
   .I3(level3_in[303]),
   .I4(level3_in[304]),
   .I5(level3_in[305])
);

LUT6 #(
   .INIT(64'hcf01a8fdcf01a8fd)  
) LUT6_inst9123 (
   .O(to_level2[51]),
   .I0(level3_in[306]),
   .I1(level3_in[307]),
   .I2(level3_in[308]),
   .I3(level3_in[309]),
   .I4(level3_in[310]),
   .I5(level3_in[311])
);

LUT6 #(
   .INIT(64'h68e7db0e68e7db0e)  
) LUT6_inst9124 (
   .O(to_level2[52]),
   .I0(level3_in[312]),
   .I1(level3_in[313]),
   .I2(level3_in[314]),
   .I3(level3_in[315]),
   .I4(level3_in[316]),
   .I5(level3_in[317])
);

LUT6 #(
   .INIT(64'h6b1c33a56b1c33a5)  
) LUT6_inst9125 (
   .O(to_level2[53]),
   .I0(level3_in[318]),
   .I1(level3_in[319]),
   .I2(level3_in[320]),
   .I3(level3_in[321]),
   .I4(level3_in[322]),
   .I5(level3_in[323])
);

LUT6 #(
   .INIT(64'hd6f7ccb4d6f7ccb4)  
) LUT6_inst9126 (
   .O(to_level2[54]),
   .I0(level3_in[324]),
   .I1(level3_in[325]),
   .I2(level3_in[326]),
   .I3(level3_in[327]),
   .I4(level3_in[328]),
   .I5(level3_in[329])
);

LUT6 #(
   .INIT(64'h68e5097068e50970)  
) LUT6_inst9127 (
   .O(to_level2[55]),
   .I0(level3_in[330]),
   .I1(level3_in[331]),
   .I2(level3_in[332]),
   .I3(level3_in[333]),
   .I4(level3_in[334]),
   .I5(level3_in[335])
);

LUT6 #(
   .INIT(64'hc441c668c441c668)  
) LUT6_inst9128 (
   .O(to_level2[56]),
   .I0(level3_in[336]),
   .I1(level3_in[337]),
   .I2(level3_in[338]),
   .I3(level3_in[339]),
   .I4(level3_in[340]),
   .I5(level3_in[341])
);

LUT6 #(
   .INIT(64'h4cb201084cb20108)  
) LUT6_inst9129 (
   .O(to_level2[57]),
   .I0(level3_in[342]),
   .I1(level3_in[343]),
   .I2(level3_in[344]),
   .I3(level3_in[345]),
   .I4(level3_in[346]),
   .I5(level3_in[347])
);

LUT6 #(
   .INIT(64'hc0453f30c0453f30)  
) LUT6_inst9130 (
   .O(to_level2[58]),
   .I0(level3_in[348]),
   .I1(level3_in[349]),
   .I2(level3_in[350]),
   .I3(level3_in[351]),
   .I4(level3_in[352]),
   .I5(level3_in[353])
);

LUT6 #(
   .INIT(64'h60e40d2060e40d20)  
) LUT6_inst9131 (
   .O(to_level2[59]),
   .I0(level3_in[354]),
   .I1(level3_in[355]),
   .I2(level3_in[356]),
   .I3(level3_in[357]),
   .I4(level3_in[358]),
   .I5(level3_in[359])
);

LUT6 #(
   .INIT(64'hb1e135dfb1e135df)  
) LUT6_inst9132 (
   .O(to_level2[60]),
   .I0(level3_in[360]),
   .I1(level3_in[361]),
   .I2(level3_in[362]),
   .I3(level3_in[363]),
   .I4(level3_in[364]),
   .I5(level3_in[365])
);

LUT6 #(
   .INIT(64'h72d184bf72d184bf)  
) LUT6_inst9133 (
   .O(to_level2[61]),
   .I0(level3_in[366]),
   .I1(level3_in[367]),
   .I2(level3_in[368]),
   .I3(level3_in[369]),
   .I4(level3_in[370]),
   .I5(level3_in[371])
);

LUT6 #(
   .INIT(64'h660ee5e4660ee5e4)  
) LUT6_inst9134 (
   .O(to_level2[62]),
   .I0(level3_in[372]),
   .I1(level3_in[373]),
   .I2(level3_in[374]),
   .I3(level3_in[375]),
   .I4(level3_in[376]),
   .I5(level3_in[377])
);

LUT6 #(
   .INIT(64'h3990594c3990594c)  
) LUT6_inst9135 (
   .O(to_level2[63]),
   .I0(level3_in[378]),
   .I1(level3_in[379]),
   .I2(level3_in[380]),
   .I3(level3_in[381]),
   .I4(level3_in[382]),
   .I5(level3_in[383])
);

LUT6 #(
   .INIT(64'h3f5a87ef3f5a87ef)  
) LUT6_inst9136 (
   .O(to_level2[64]),
   .I0(level3_in[384]),
   .I1(level3_in[385]),
   .I2(level3_in[386]),
   .I3(level3_in[387]),
   .I4(level3_in[388]),
   .I5(level3_in[389])
);

LUT6 #(
   .INIT(64'he4522995e4522995)  
) LUT6_inst9137 (
   .O(to_level2[65]),
   .I0(level3_in[390]),
   .I1(level3_in[391]),
   .I2(level3_in[392]),
   .I3(level3_in[393]),
   .I4(level3_in[394]),
   .I5(level3_in[395])
);

LUT6 #(
   .INIT(64'hc7928b6ec7928b6e)  
) LUT6_inst9138 (
   .O(to_level2[66]),
   .I0(level3_in[396]),
   .I1(level3_in[397]),
   .I2(level3_in[398]),
   .I3(level3_in[399]),
   .I4(level3_in[400]),
   .I5(level3_in[401])
);

LUT6 #(
   .INIT(64'h3f1a313b3f1a313b)  
) LUT6_inst9139 (
   .O(to_level2[67]),
   .I0(level3_in[402]),
   .I1(level3_in[403]),
   .I2(level3_in[404]),
   .I3(level3_in[405]),
   .I4(level3_in[406]),
   .I5(level3_in[407])
);

LUT6 #(
   .INIT(64'h7cbddc087cbddc08)  
) LUT6_inst9140 (
   .O(to_level2[68]),
   .I0(level3_in[408]),
   .I1(level3_in[409]),
   .I2(level3_in[410]),
   .I3(level3_in[411]),
   .I4(level3_in[412]),
   .I5(level3_in[413])
);

LUT6 #(
   .INIT(64'h926b1d5a926b1d5a)  
) LUT6_inst9141 (
   .O(to_level2[69]),
   .I0(level3_in[414]),
   .I1(level3_in[415]),
   .I2(level3_in[416]),
   .I3(level3_in[417]),
   .I4(level3_in[418]),
   .I5(level3_in[419])
);

LUT6 #(
   .INIT(64'h3bc2a1e23bc2a1e2)  
) LUT6_inst9142 (
   .O(to_level2[70]),
   .I0(level3_in[420]),
   .I1(level3_in[421]),
   .I2(level3_in[422]),
   .I3(level3_in[423]),
   .I4(level3_in[424]),
   .I5(level3_in[425])
);

LUT6 #(
   .INIT(64'h35edbb2735edbb27)  
) LUT6_inst9143 (
   .O(to_level2[71]),
   .I0(level3_in[426]),
   .I1(level3_in[427]),
   .I2(level3_in[428]),
   .I3(level3_in[429]),
   .I4(level3_in[430]),
   .I5(level3_in[431])
);

LUT6 #(
   .INIT(64'hdb68e26fdb68e26f)  
) LUT6_inst9144 (
   .O(to_level2[72]),
   .I0(level3_in[432]),
   .I1(level3_in[433]),
   .I2(level3_in[434]),
   .I3(level3_in[435]),
   .I4(level3_in[436]),
   .I5(level3_in[437])
);

LUT6 #(
   .INIT(64'hf4de0eb4f4de0eb4)  
) LUT6_inst9145 (
   .O(to_level2[73]),
   .I0(level3_in[438]),
   .I1(level3_in[439]),
   .I2(level3_in[440]),
   .I3(level3_in[441]),
   .I4(level3_in[442]),
   .I5(level3_in[443])
);

LUT6 #(
   .INIT(64'h03ba47b703ba47b7)  
) LUT6_inst9146 (
   .O(to_level2[74]),
   .I0(level3_in[444]),
   .I1(level3_in[445]),
   .I2(level3_in[446]),
   .I3(level3_in[447]),
   .I4(level3_in[448]),
   .I5(level3_in[449])
);

LUT6 #(
   .INIT(64'heae36e3feae36e3f)  
) LUT6_inst9147 (
   .O(to_level2[75]),
   .I0(level3_in[450]),
   .I1(level3_in[451]),
   .I2(level3_in[452]),
   .I3(level3_in[453]),
   .I4(level3_in[454]),
   .I5(level3_in[455])
);

LUT6 #(
   .INIT(64'hb9643b50b9643b50)  
) LUT6_inst9148 (
   .O(to_level2[76]),
   .I0(level3_in[456]),
   .I1(level3_in[457]),
   .I2(level3_in[458]),
   .I3(level3_in[459]),
   .I4(level3_in[460]),
   .I5(level3_in[461])
);

LUT6 #(
   .INIT(64'h3bca7a2a3bca7a2a)  
) LUT6_inst9149 (
   .O(to_level2[77]),
   .I0(level3_in[462]),
   .I1(level3_in[463]),
   .I2(level3_in[464]),
   .I3(level3_in[465]),
   .I4(level3_in[466]),
   .I5(level3_in[467])
);

LUT6 #(
   .INIT(64'he8f02ef9e8f02ef9)  
) LUT6_inst9150 (
   .O(to_level2[78]),
   .I0(level3_in[468]),
   .I1(level3_in[469]),
   .I2(level3_in[470]),
   .I3(level3_in[471]),
   .I4(level3_in[472]),
   .I5(level3_in[473])
);

LUT6 #(
   .INIT(64'h50709f6650709f66)  
) LUT6_inst9151 (
   .O(to_level2[79]),
   .I0(level3_in[474]),
   .I1(level3_in[475]),
   .I2(level3_in[476]),
   .I3(level3_in[477]),
   .I4(level3_in[478]),
   .I5(level3_in[479])
);

LUT6 #(
   .INIT(64'hebe8b7f7ebe8b7f7)  
) LUT6_inst9152 (
   .O(to_level2[80]),
   .I0(level3_in[480]),
   .I1(level3_in[481]),
   .I2(level3_in[482]),
   .I3(level3_in[483]),
   .I4(level3_in[484]),
   .I5(level3_in[485])
);

LUT6 #(
   .INIT(64'h009c813a009c813a)  
) LUT6_inst9153 (
   .O(to_level2[81]),
   .I0(level3_in[486]),
   .I1(level3_in[487]),
   .I2(level3_in[488]),
   .I3(level3_in[489]),
   .I4(level3_in[490]),
   .I5(level3_in[491])
);

LUT6 #(
   .INIT(64'h7a99b6d97a99b6d9)  
) LUT6_inst9154 (
   .O(to_level2[82]),
   .I0(level3_in[492]),
   .I1(level3_in[493]),
   .I2(level3_in[494]),
   .I3(level3_in[495]),
   .I4(level3_in[496]),
   .I5(level3_in[497])
);

LUT6 #(
   .INIT(64'ha74736a3a74736a3)  
) LUT6_inst9155 (
   .O(to_level2[83]),
   .I0(level3_in[498]),
   .I1(level3_in[499]),
   .I2(level3_in[500]),
   .I3(level3_in[501]),
   .I4(level3_in[502]),
   .I5(level3_in[503])
);

LUT6 #(
   .INIT(64'h0fa637380fa63738)  
) LUT6_inst9156 (
   .O(to_level2[84]),
   .I0(level3_in[504]),
   .I1(level3_in[505]),
   .I2(level3_in[506]),
   .I3(level3_in[507]),
   .I4(level3_in[508]),
   .I5(level3_in[509])
);

LUT6 #(
   .INIT(64'h155a0147155a0147)  
) LUT6_inst9157 (
   .O(to_level2[85]),
   .I0(level3_in[510]),
   .I1(level3_in[511]),
   .I2(level3_in[512]),
   .I3(level3_in[513]),
   .I4(level3_in[514]),
   .I5(level3_in[515])
);

LUT6 #(
   .INIT(64'ha3f7e12da3f7e12d)  
) LUT6_inst9158 (
   .O(to_level2[86]),
   .I0(level3_in[516]),
   .I1(level3_in[517]),
   .I2(level3_in[518]),
   .I3(level3_in[519]),
   .I4(level3_in[520]),
   .I5(level3_in[521])
);

LUT6 #(
   .INIT(64'h1464dac41464dac4)  
) LUT6_inst9159 (
   .O(to_level2[87]),
   .I0(level3_in[522]),
   .I1(level3_in[523]),
   .I2(level3_in[524]),
   .I3(level3_in[525]),
   .I4(level3_in[526]),
   .I5(level3_in[527])
);

LUT6 #(
   .INIT(64'h2abf1d1b2abf1d1b)  
) LUT6_inst9160 (
   .O(to_level2[88]),
   .I0(level3_in[528]),
   .I1(level3_in[529]),
   .I2(level3_in[530]),
   .I3(level3_in[531]),
   .I4(level3_in[532]),
   .I5(level3_in[533])
);

LUT6 #(
   .INIT(64'h34384b9734384b97)  
) LUT6_inst9161 (
   .O(to_level2[89]),
   .I0(level3_in[534]),
   .I1(level3_in[535]),
   .I2(level3_in[536]),
   .I3(level3_in[537]),
   .I4(level3_in[538]),
   .I5(level3_in[539])
);

LUT6 #(
   .INIT(64'h67d792fc67d792fc)  
) LUT6_inst9162 (
   .O(to_level2[90]),
   .I0(level3_in[540]),
   .I1(level3_in[541]),
   .I2(level3_in[542]),
   .I3(level3_in[543]),
   .I4(level3_in[544]),
   .I5(level3_in[545])
);

LUT6 #(
   .INIT(64'h2574b4782574b478)  
) LUT6_inst9163 (
   .O(to_level2[91]),
   .I0(level3_in[546]),
   .I1(level3_in[547]),
   .I2(level3_in[548]),
   .I3(level3_in[549]),
   .I4(level3_in[550]),
   .I5(level3_in[551])
);

LUT6 #(
   .INIT(64'h5cac5b6a5cac5b6a)  
) LUT6_inst9164 (
   .O(to_level2[92]),
   .I0(level3_in[552]),
   .I1(level3_in[553]),
   .I2(level3_in[554]),
   .I3(level3_in[555]),
   .I4(level3_in[556]),
   .I5(level3_in[557])
);

LUT6 #(
   .INIT(64'h80196e5480196e54)  
) LUT6_inst9165 (
   .O(to_level2[93]),
   .I0(level3_in[558]),
   .I1(level3_in[559]),
   .I2(level3_in[560]),
   .I3(level3_in[561]),
   .I4(level3_in[562]),
   .I5(level3_in[563])
);

LUT6 #(
   .INIT(64'h007409e7007409e7)  
) LUT6_inst9166 (
   .O(to_level2[94]),
   .I0(level3_in[564]),
   .I1(level3_in[565]),
   .I2(level3_in[566]),
   .I3(level3_in[567]),
   .I4(level3_in[568]),
   .I5(level3_in[569])
);

LUT6 #(
   .INIT(64'h625cbc76625cbc76)  
) LUT6_inst9167 (
   .O(to_level2[95]),
   .I0(level3_in[570]),
   .I1(level3_in[571]),
   .I2(level3_in[572]),
   .I3(level3_in[573]),
   .I4(level3_in[574]),
   .I5(level3_in[575])
);

LUT6 #(
   .INIT(64'hec48a4d8ec48a4d8)  
) LUT6_inst9168 (
   .O(to_level2[96]),
   .I0(level3_in[576]),
   .I1(level3_in[577]),
   .I2(level3_in[578]),
   .I3(level3_in[579]),
   .I4(level3_in[580]),
   .I5(level3_in[581])
);

LUT6 #(
   .INIT(64'h240a2caf240a2caf)  
) LUT6_inst9169 (
   .O(to_level2[97]),
   .I0(level3_in[582]),
   .I1(level3_in[583]),
   .I2(level3_in[584]),
   .I3(level3_in[585]),
   .I4(level3_in[586]),
   .I5(level3_in[587])
);

LUT6 #(
   .INIT(64'hd1634bcfd1634bcf)  
) LUT6_inst9170 (
   .O(to_level2[98]),
   .I0(level3_in[588]),
   .I1(level3_in[589]),
   .I2(level3_in[590]),
   .I3(level3_in[591]),
   .I4(level3_in[592]),
   .I5(level3_in[593])
);

LUT6 #(
   .INIT(64'haa627b36aa627b36)  
) LUT6_inst9171 (
   .O(to_level2[99]),
   .I0(level3_in[594]),
   .I1(level3_in[595]),
   .I2(level3_in[596]),
   .I3(level3_in[597]),
   .I4(level3_in[598]),
   .I5(level3_in[599])
);

LUT6 #(
   .INIT(64'h49066b2749066b27)  
) LUT6_inst9172 (
   .O(to_level2[100]),
   .I0(level3_in[600]),
   .I1(level3_in[601]),
   .I2(level3_in[602]),
   .I3(level3_in[603]),
   .I4(level3_in[604]),
   .I5(level3_in[605])
);

LUT6 #(
   .INIT(64'h6583e67b6583e67b)  
) LUT6_inst9173 (
   .O(to_level2[101]),
   .I0(level3_in[606]),
   .I1(level3_in[607]),
   .I2(level3_in[608]),
   .I3(level3_in[609]),
   .I4(level3_in[610]),
   .I5(level3_in[611])
);

LUT6 #(
   .INIT(64'h47c80b1b47c80b1b)  
) LUT6_inst9174 (
   .O(to_level2[102]),
   .I0(level3_in[612]),
   .I1(level3_in[613]),
   .I2(level3_in[614]),
   .I3(level3_in[615]),
   .I4(level3_in[616]),
   .I5(level3_in[617])
);

LUT6 #(
   .INIT(64'hb4543b47b4543b47)  
) LUT6_inst9175 (
   .O(to_level2[103]),
   .I0(level3_in[618]),
   .I1(level3_in[619]),
   .I2(level3_in[620]),
   .I3(level3_in[621]),
   .I4(level3_in[622]),
   .I5(level3_in[623])
);

LUT6 #(
   .INIT(64'hfb8994e2fb8994e2)  
) LUT6_inst9176 (
   .O(to_level2[104]),
   .I0(level3_in[624]),
   .I1(level3_in[625]),
   .I2(level3_in[626]),
   .I3(level3_in[627]),
   .I4(level3_in[628]),
   .I5(level3_in[629])
);

LUT6 #(
   .INIT(64'hdd9dbdb1dd9dbdb1)  
) LUT6_inst9177 (
   .O(to_level2[105]),
   .I0(level3_in[630]),
   .I1(level3_in[631]),
   .I2(level3_in[632]),
   .I3(level3_in[633]),
   .I4(level3_in[634]),
   .I5(level3_in[635])
);

LUT6 #(
   .INIT(64'h15e28c7815e28c78)  
) LUT6_inst9178 (
   .O(to_level2[106]),
   .I0(level3_in[636]),
   .I1(level3_in[637]),
   .I2(level3_in[638]),
   .I3(level3_in[639]),
   .I4(level3_in[640]),
   .I5(level3_in[641])
);

LUT6 #(
   .INIT(64'hc351b6ebc351b6eb)  
) LUT6_inst9179 (
   .O(to_level2[107]),
   .I0(level3_in[642]),
   .I1(level3_in[643]),
   .I2(level3_in[644]),
   .I3(level3_in[645]),
   .I4(level3_in[646]),
   .I5(level3_in[647])
);

LUT6 #(
   .INIT(64'hb3fde267b3fde267)  
) LUT6_inst9180 (
   .O(to_level2[108]),
   .I0(level3_in[648]),
   .I1(level3_in[649]),
   .I2(level3_in[650]),
   .I3(level3_in[651]),
   .I4(level3_in[652]),
   .I5(level3_in[653])
);

LUT6 #(
   .INIT(64'h03a9454d03a9454d)  
) LUT6_inst9181 (
   .O(to_level2[109]),
   .I0(level3_in[654]),
   .I1(level3_in[655]),
   .I2(level3_in[656]),
   .I3(level3_in[657]),
   .I4(level3_in[658]),
   .I5(level3_in[659])
);

LUT6 #(
   .INIT(64'h09ade43509ade435)  
) LUT6_inst9182 (
   .O(to_level2[110]),
   .I0(level3_in[660]),
   .I1(level3_in[661]),
   .I2(level3_in[662]),
   .I3(level3_in[663]),
   .I4(level3_in[664]),
   .I5(level3_in[665])
);

LUT6 #(
   .INIT(64'h0ef0867b0ef0867b)  
) LUT6_inst9183 (
   .O(to_level2[111]),
   .I0(level3_in[666]),
   .I1(level3_in[667]),
   .I2(level3_in[668]),
   .I3(level3_in[669]),
   .I4(level3_in[670]),
   .I5(level3_in[671])
);

LUT6 #(
   .INIT(64'h7bddab287bddab28)  
) LUT6_inst9184 (
   .O(to_level2[112]),
   .I0(level3_in[672]),
   .I1(level3_in[673]),
   .I2(level3_in[674]),
   .I3(level3_in[675]),
   .I4(level3_in[676]),
   .I5(level3_in[677])
);

LUT6 #(
   .INIT(64'hd347efc2d347efc2)  
) LUT6_inst9185 (
   .O(to_level2[113]),
   .I0(level3_in[678]),
   .I1(level3_in[679]),
   .I2(level3_in[680]),
   .I3(level3_in[681]),
   .I4(level3_in[682]),
   .I5(level3_in[683])
);

LUT6 #(
   .INIT(64'h0743a7b60743a7b6)  
) LUT6_inst9186 (
   .O(to_level2[114]),
   .I0(level3_in[684]),
   .I1(level3_in[685]),
   .I2(level3_in[686]),
   .I3(level3_in[687]),
   .I4(level3_in[688]),
   .I5(level3_in[689])
);

LUT6 #(
   .INIT(64'hd727f701d727f701)  
) LUT6_inst9187 (
   .O(to_level2[115]),
   .I0(level3_in[690]),
   .I1(level3_in[691]),
   .I2(level3_in[692]),
   .I3(level3_in[693]),
   .I4(level3_in[694]),
   .I5(level3_in[695])
);

LUT6 #(
   .INIT(64'h4310c46b4310c46b)  
) LUT6_inst9188 (
   .O(to_level2[116]),
   .I0(level3_in[696]),
   .I1(level3_in[697]),
   .I2(level3_in[698]),
   .I3(level3_in[699]),
   .I4(level3_in[700]),
   .I5(level3_in[701])
);

LUT6 #(
   .INIT(64'h33d4a0e533d4a0e5)  
) LUT6_inst9189 (
   .O(to_level2[117]),
   .I0(level3_in[702]),
   .I1(level3_in[703]),
   .I2(level3_in[704]),
   .I3(level3_in[705]),
   .I4(level3_in[706]),
   .I5(level3_in[707])
);

LUT6 #(
   .INIT(64'h5f773a265f773a26)  
) LUT6_inst9190 (
   .O(to_level2[118]),
   .I0(level3_in[708]),
   .I1(level3_in[709]),
   .I2(level3_in[710]),
   .I3(level3_in[711]),
   .I4(level3_in[712]),
   .I5(level3_in[713])
);

LUT6 #(
   .INIT(64'hc959b3cfc959b3cf)  
) LUT6_inst9191 (
   .O(to_level2[119]),
   .I0(level3_in[714]),
   .I1(level3_in[715]),
   .I2(level3_in[716]),
   .I3(level3_in[717]),
   .I4(level3_in[718]),
   .I5(level3_in[719])
);

LUT6 #(
   .INIT(64'h4619f35d4619f35d)  
) LUT6_inst9192 (
   .O(to_level2[120]),
   .I0(level3_in[720]),
   .I1(level3_in[721]),
   .I2(level3_in[722]),
   .I3(level3_in[723]),
   .I4(level3_in[724]),
   .I5(level3_in[725])
);

LUT6 #(
   .INIT(64'h41c63a1141c63a11)  
) LUT6_inst9193 (
   .O(to_level2[121]),
   .I0(level3_in[726]),
   .I1(level3_in[727]),
   .I2(level3_in[728]),
   .I3(level3_in[729]),
   .I4(level3_in[730]),
   .I5(level3_in[731])
);

LUT6 #(
   .INIT(64'h262d84b1262d84b1)  
) LUT6_inst9194 (
   .O(to_level2[122]),
   .I0(level3_in[732]),
   .I1(level3_in[733]),
   .I2(level3_in[734]),
   .I3(level3_in[735]),
   .I4(level3_in[736]),
   .I5(level3_in[737])
);

LUT6 #(
   .INIT(64'h8545589785455897)  
) LUT6_inst9195 (
   .O(to_level2[123]),
   .I0(level3_in[738]),
   .I1(level3_in[739]),
   .I2(level3_in[740]),
   .I3(level3_in[741]),
   .I4(level3_in[742]),
   .I5(level3_in[743])
);

LUT6 #(
   .INIT(64'he7996dfde7996dfd)  
) LUT6_inst9196 (
   .O(to_level2[124]),
   .I0(level3_in[744]),
   .I1(level3_in[745]),
   .I2(level3_in[746]),
   .I3(level3_in[747]),
   .I4(level3_in[748]),
   .I5(level3_in[749])
);

LUT6 #(
   .INIT(64'h5525e3f45525e3f4)  
) LUT6_inst9197 (
   .O(to_level2[125]),
   .I0(level3_in[750]),
   .I1(level3_in[751]),
   .I2(level3_in[752]),
   .I3(level3_in[753]),
   .I4(level3_in[754]),
   .I5(level3_in[755])
);

LUT6 #(
   .INIT(64'hebe01b69ebe01b69)  
) LUT6_inst9198 (
   .O(to_level2[126]),
   .I0(level3_in[756]),
   .I1(level3_in[757]),
   .I2(level3_in[758]),
   .I3(level3_in[759]),
   .I4(level3_in[760]),
   .I5(level3_in[761])
);

LUT6 #(
   .INIT(64'he615f265e615f265)  
) LUT6_inst9199 (
   .O(to_level2[127]),
   .I0(level3_in[762]),
   .I1(level3_in[763]),
   .I2(level3_in[764]),
   .I3(level3_in[765]),
   .I4(level3_in[766]),
   .I5(level3_in[767])
);

LUT6 #(
   .INIT(64'ha1ba2a6fa1ba2a6f)  
) LUT6_inst9200 (
   .O(to_level2[128]),
   .I0(level3_in[768]),
   .I1(level3_in[769]),
   .I2(level3_in[770]),
   .I3(level3_in[771]),
   .I4(level3_in[772]),
   .I5(level3_in[773])
);

LUT6 #(
   .INIT(64'hcd40a0a3cd40a0a3)  
) LUT6_inst9201 (
   .O(to_level2[129]),
   .I0(level3_in[774]),
   .I1(level3_in[775]),
   .I2(level3_in[776]),
   .I3(level3_in[777]),
   .I4(level3_in[778]),
   .I5(level3_in[779])
);

LUT6 #(
   .INIT(64'h358d5736358d5736)  
) LUT6_inst9202 (
   .O(to_level2[130]),
   .I0(level3_in[780]),
   .I1(level3_in[781]),
   .I2(level3_in[782]),
   .I3(level3_in[783]),
   .I4(level3_in[784]),
   .I5(level3_in[785])
);

LUT6 #(
   .INIT(64'hf1617d06f1617d06)  
) LUT6_inst9203 (
   .O(to_level2[131]),
   .I0(level3_in[786]),
   .I1(level3_in[787]),
   .I2(level3_in[788]),
   .I3(level3_in[789]),
   .I4(level3_in[790]),
   .I5(level3_in[791])
);

LUT6 #(
   .INIT(64'h3717b06d3717b06d)  
) LUT6_inst9204 (
   .O(to_level2[132]),
   .I0(level3_in[792]),
   .I1(level3_in[793]),
   .I2(level3_in[794]),
   .I3(level3_in[795]),
   .I4(level3_in[796]),
   .I5(level3_in[797])
);

LUT6 #(
   .INIT(64'h31f5349431f53494)  
) LUT6_inst9205 (
   .O(to_level2[133]),
   .I0(level3_in[798]),
   .I1(level3_in[799]),
   .I2(level3_in[800]),
   .I3(level3_in[801]),
   .I4(level3_in[802]),
   .I5(level3_in[803])
);

LUT6 #(
   .INIT(64'he55a0de2e55a0de2)  
) LUT6_inst9206 (
   .O(to_level2[134]),
   .I0(level3_in[804]),
   .I1(level3_in[805]),
   .I2(level3_in[806]),
   .I3(level3_in[807]),
   .I4(level3_in[808]),
   .I5(level3_in[809])
);

LUT6 #(
   .INIT(64'he24e482be24e482b)  
) LUT6_inst9207 (
   .O(to_level2[135]),
   .I0(level3_in[810]),
   .I1(level3_in[811]),
   .I2(level3_in[812]),
   .I3(level3_in[813]),
   .I4(level3_in[814]),
   .I5(level3_in[815])
);

LUT6 #(
   .INIT(64'h56a478e356a478e3)  
) LUT6_inst9208 (
   .O(to_level2[136]),
   .I0(level3_in[816]),
   .I1(level3_in[817]),
   .I2(level3_in[818]),
   .I3(level3_in[819]),
   .I4(level3_in[820]),
   .I5(level3_in[821])
);

LUT6 #(
   .INIT(64'h5170b8c65170b8c6)  
) LUT6_inst9209 (
   .O(to_level2[137]),
   .I0(level3_in[822]),
   .I1(level3_in[823]),
   .I2(level3_in[824]),
   .I3(level3_in[825]),
   .I4(level3_in[826]),
   .I5(level3_in[827])
);

LUT6 #(
   .INIT(64'hb3fae75eb3fae75e)  
) LUT6_inst9210 (
   .O(to_level2[138]),
   .I0(level3_in[828]),
   .I1(level3_in[829]),
   .I2(level3_in[830]),
   .I3(level3_in[831]),
   .I4(level3_in[832]),
   .I5(level3_in[833])
);

LUT6 #(
   .INIT(64'hfc0c707cfc0c707c)  
) LUT6_inst9211 (
   .O(to_level2[139]),
   .I0(level3_in[834]),
   .I1(level3_in[835]),
   .I2(level3_in[836]),
   .I3(level3_in[837]),
   .I4(level3_in[838]),
   .I5(level3_in[839])
);

LUT6 #(
   .INIT(64'h22c3399322c33993)  
) LUT6_inst9212 (
   .O(to_level2[140]),
   .I0(level3_in[840]),
   .I1(level3_in[841]),
   .I2(level3_in[842]),
   .I3(level3_in[843]),
   .I4(level3_in[844]),
   .I5(level3_in[845])
);

LUT6 #(
   .INIT(64'h27674f6827674f68)  
) LUT6_inst9213 (
   .O(to_level2[141]),
   .I0(level3_in[846]),
   .I1(level3_in[847]),
   .I2(level3_in[848]),
   .I3(level3_in[849]),
   .I4(level3_in[850]),
   .I5(level3_in[851])
);

LUT6 #(
   .INIT(64'hef7f1d1cef7f1d1c)  
) LUT6_inst9214 (
   .O(to_level2[142]),
   .I0(level3_in[852]),
   .I1(level3_in[853]),
   .I2(level3_in[854]),
   .I3(level3_in[855]),
   .I4(level3_in[856]),
   .I5(level3_in[857])
);

LUT6 #(
   .INIT(64'hac78e453ac78e453)  
) LUT6_inst9215 (
   .O(to_level2[143]),
   .I0(level3_in[858]),
   .I1(level3_in[859]),
   .I2(level3_in[860]),
   .I3(level3_in[861]),
   .I4(level3_in[862]),
   .I5(level3_in[863])
);

LUT6 #(
   .INIT(64'ha8438d05a8438d05)  
) LUT6_inst9216 (
   .O(to_level2[144]),
   .I0(level3_in[864]),
   .I1(level3_in[865]),
   .I2(level3_in[866]),
   .I3(level3_in[867]),
   .I4(level3_in[868]),
   .I5(level3_in[869])
);

LUT6 #(
   .INIT(64'h93ae535093ae5350)  
) LUT6_inst9217 (
   .O(to_level2[145]),
   .I0(level3_in[870]),
   .I1(level3_in[871]),
   .I2(level3_in[872]),
   .I3(level3_in[873]),
   .I4(level3_in[874]),
   .I5(level3_in[875])
);

LUT6 #(
   .INIT(64'h846488c6846488c6)  
) LUT6_inst9218 (
   .O(to_level2[146]),
   .I0(level3_in[876]),
   .I1(level3_in[877]),
   .I2(level3_in[878]),
   .I3(level3_in[879]),
   .I4(level3_in[880]),
   .I5(level3_in[881])
);

LUT6 #(
   .INIT(64'h99ecf34299ecf342)  
) LUT6_inst9219 (
   .O(to_level2[147]),
   .I0(level3_in[882]),
   .I1(level3_in[883]),
   .I2(level3_in[884]),
   .I3(level3_in[885]),
   .I4(level3_in[886]),
   .I5(level3_in[887])
);

LUT6 #(
   .INIT(64'h3e5eacc23e5eacc2)  
) LUT6_inst9220 (
   .O(to_level2[148]),
   .I0(level3_in[888]),
   .I1(level3_in[889]),
   .I2(level3_in[890]),
   .I3(level3_in[891]),
   .I4(level3_in[892]),
   .I5(level3_in[893])
);

LUT6 #(
   .INIT(64'hffc45988ffc45988)  
) LUT6_inst9221 (
   .O(to_level2[149]),
   .I0(level3_in[894]),
   .I1(level3_in[895]),
   .I2(level3_in[896]),
   .I3(level3_in[897]),
   .I4(level3_in[898]),
   .I5(level3_in[899])
);

LUT6 #(
   .INIT(64'h12a2d0d912a2d0d9)  
) LUT6_inst9222 (
   .O(to_level2[150]),
   .I0(level3_in[900]),
   .I1(level3_in[901]),
   .I2(level3_in[902]),
   .I3(level3_in[903]),
   .I4(level3_in[904]),
   .I5(level3_in[905])
);

LUT6 #(
   .INIT(64'ha1debe9ba1debe9b)  
) LUT6_inst9223 (
   .O(to_level2[151]),
   .I0(level3_in[906]),
   .I1(level3_in[907]),
   .I2(level3_in[908]),
   .I3(level3_in[909]),
   .I4(level3_in[910]),
   .I5(level3_in[911])
);

LUT6 #(
   .INIT(64'h438c803a438c803a)  
) LUT6_inst9224 (
   .O(to_level2[152]),
   .I0(level3_in[912]),
   .I1(level3_in[913]),
   .I2(level3_in[914]),
   .I3(level3_in[915]),
   .I4(level3_in[916]),
   .I5(level3_in[917])
);

LUT6 #(
   .INIT(64'h9e861acf9e861acf)  
) LUT6_inst9225 (
   .O(to_level2[153]),
   .I0(level3_in[918]),
   .I1(level3_in[919]),
   .I2(level3_in[920]),
   .I3(level3_in[921]),
   .I4(level3_in[922]),
   .I5(level3_in[923])
);

LUT6 #(
   .INIT(64'h057f12b7057f12b7)  
) LUT6_inst9226 (
   .O(to_level2[154]),
   .I0(level3_in[924]),
   .I1(level3_in[925]),
   .I2(level3_in[926]),
   .I3(level3_in[927]),
   .I4(level3_in[928]),
   .I5(level3_in[929])
);

LUT6 #(
   .INIT(64'hb9510287b9510287)  
) LUT6_inst9227 (
   .O(to_level2[155]),
   .I0(level3_in[930]),
   .I1(level3_in[931]),
   .I2(level3_in[932]),
   .I3(level3_in[933]),
   .I4(level3_in[934]),
   .I5(level3_in[935])
);

LUT6 #(
   .INIT(64'h7cd094c17cd094c1)  
) LUT6_inst9228 (
   .O(to_level2[156]),
   .I0(level3_in[936]),
   .I1(level3_in[937]),
   .I2(level3_in[938]),
   .I3(level3_in[939]),
   .I4(level3_in[940]),
   .I5(level3_in[941])
);

LUT6 #(
   .INIT(64'h0a2c2ea80a2c2ea8)  
) LUT6_inst9229 (
   .O(to_level2[157]),
   .I0(level3_in[942]),
   .I1(level3_in[943]),
   .I2(level3_in[944]),
   .I3(level3_in[945]),
   .I4(level3_in[946]),
   .I5(level3_in[947])
);

LUT6 #(
   .INIT(64'h1f9d35a41f9d35a4)  
) LUT6_inst9230 (
   .O(to_level2[158]),
   .I0(level3_in[948]),
   .I1(level3_in[949]),
   .I2(level3_in[950]),
   .I3(level3_in[951]),
   .I4(level3_in[952]),
   .I5(level3_in[953])
);

LUT6 #(
   .INIT(64'hd1e42335d1e42335)  
) LUT6_inst9231 (
   .O(to_level2[159]),
   .I0(level3_in[954]),
   .I1(level3_in[955]),
   .I2(level3_in[956]),
   .I3(level3_in[957]),
   .I4(level3_in[958]),
   .I5(level3_in[959])
);

LUT6 #(
   .INIT(64'h99ba219f99ba219f)  
) LUT6_inst9232 (
   .O(to_level2[160]),
   .I0(level3_in[960]),
   .I1(level3_in[961]),
   .I2(level3_in[962]),
   .I3(level3_in[963]),
   .I4(level3_in[964]),
   .I5(level3_in[965])
);

LUT6 #(
   .INIT(64'he74ddedae74ddeda)  
) LUT6_inst9233 (
   .O(to_level2[161]),
   .I0(level3_in[966]),
   .I1(level3_in[967]),
   .I2(level3_in[968]),
   .I3(level3_in[969]),
   .I4(level3_in[970]),
   .I5(level3_in[971])
);

LUT6 #(
   .INIT(64'h1c2bc7de1c2bc7de)  
) LUT6_inst9234 (
   .O(to_level2[162]),
   .I0(level3_in[972]),
   .I1(level3_in[973]),
   .I2(level3_in[974]),
   .I3(level3_in[975]),
   .I4(level3_in[976]),
   .I5(level3_in[977])
);

LUT6 #(
   .INIT(64'h605240b5605240b5)  
) LUT6_inst9235 (
   .O(to_level2[163]),
   .I0(level3_in[978]),
   .I1(level3_in[979]),
   .I2(level3_in[980]),
   .I3(level3_in[981]),
   .I4(level3_in[982]),
   .I5(level3_in[983])
);

LUT6 #(
   .INIT(64'h7209f5e27209f5e2)  
) LUT6_inst9236 (
   .O(to_level2[164]),
   .I0(level3_in[984]),
   .I1(level3_in[985]),
   .I2(level3_in[986]),
   .I3(level3_in[987]),
   .I4(level3_in[988]),
   .I5(level3_in[989])
);

LUT6 #(
   .INIT(64'h20ea03d020ea03d0)  
) LUT6_inst9237 (
   .O(to_level2[165]),
   .I0(level3_in[990]),
   .I1(level3_in[991]),
   .I2(level3_in[992]),
   .I3(level3_in[993]),
   .I4(level3_in[994]),
   .I5(level3_in[995])
);

LUT6 #(
   .INIT(64'h10a3e27110a3e271)  
) LUT6_inst9238 (
   .O(to_level2[166]),
   .I0(level3_in[996]),
   .I1(level3_in[997]),
   .I2(level3_in[998]),
   .I3(level3_in[999]),
   .I4(level3_in[1000]),
   .I5(level3_in[1001])
);

LUT6 #(
   .INIT(64'hb7d50afdb7d50afd)  
) LUT6_inst9239 (
   .O(to_level2[167]),
   .I0(level3_in[1002]),
   .I1(level3_in[1003]),
   .I2(level3_in[1004]),
   .I3(level3_in[1005]),
   .I4(level3_in[1006]),
   .I5(level3_in[1007])
);

LUT6 #(
   .INIT(64'h36e499ba36e499ba)  
) LUT6_inst9240 (
   .O(to_level2[168]),
   .I0(level3_in[1008]),
   .I1(level3_in[1009]),
   .I2(level3_in[1010]),
   .I3(level3_in[1011]),
   .I4(level3_in[1012]),
   .I5(level3_in[1013])
);

LUT6 #(
   .INIT(64'haa92270daa92270d)  
) LUT6_inst9241 (
   .O(to_level2[169]),
   .I0(level3_in[1014]),
   .I1(level3_in[1015]),
   .I2(level3_in[1016]),
   .I3(level3_in[1017]),
   .I4(level3_in[1018]),
   .I5(level3_in[1019])
);

LUT6 #(
   .INIT(64'h260d7162260d7162)  
) LUT6_inst9242 (
   .O(to_level2[170]),
   .I0(level3_in[1020]),
   .I1(level3_in[1021]),
   .I2(level3_in[1022]),
   .I3(level3_in[1023]),
   .I4(level3_in[1024]),
   .I5(level3_in[1025])
);

LUT6 #(
   .INIT(64'h6d1fd5da6d1fd5da)  
) LUT6_inst9243 (
   .O(to_level2[171]),
   .I0(level3_in[1026]),
   .I1(level3_in[1027]),
   .I2(level3_in[1028]),
   .I3(level3_in[1029]),
   .I4(level3_in[1030]),
   .I5(level3_in[1031])
);

LUT6 #(
   .INIT(64'h2ff11afe2ff11afe)  
) LUT6_inst9244 (
   .O(to_level2[172]),
   .I0(level3_in[1032]),
   .I1(level3_in[1033]),
   .I2(level3_in[1034]),
   .I3(level3_in[1035]),
   .I4(level3_in[1036]),
   .I5(level3_in[1037])
);

LUT6 #(
   .INIT(64'ha12f95b4a12f95b4)  
) LUT6_inst9245 (
   .O(to_level2[173]),
   .I0(level3_in[1038]),
   .I1(level3_in[1039]),
   .I2(level3_in[1040]),
   .I3(level3_in[1041]),
   .I4(level3_in[1042]),
   .I5(level3_in[1043])
);

LUT6 #(
   .INIT(64'ha59ee2aaa59ee2aa)  
) LUT6_inst9246 (
   .O(to_level2[174]),
   .I0(level3_in[1044]),
   .I1(level3_in[1045]),
   .I2(level3_in[1046]),
   .I3(level3_in[1047]),
   .I4(level3_in[1048]),
   .I5(level3_in[1049])
);

LUT6 #(
   .INIT(64'h3524b3293524b329)  
) LUT6_inst9247 (
   .O(to_level2[175]),
   .I0(level3_in[1050]),
   .I1(level3_in[1051]),
   .I2(level3_in[1052]),
   .I3(level3_in[1053]),
   .I4(level3_in[1054]),
   .I5(level3_in[1055])
);

LUT6 #(
   .INIT(64'h8d5475a78d5475a7)  
) LUT6_inst9248 (
   .O(to_level2[176]),
   .I0(level3_in[1056]),
   .I1(level3_in[1057]),
   .I2(level3_in[1058]),
   .I3(level3_in[1059]),
   .I4(level3_in[1060]),
   .I5(level3_in[1061])
);

LUT6 #(
   .INIT(64'h6ac9062f6ac9062f)  
) LUT6_inst9249 (
   .O(to_level2[177]),
   .I0(level3_in[1062]),
   .I1(level3_in[1063]),
   .I2(level3_in[1064]),
   .I3(level3_in[1065]),
   .I4(level3_in[1066]),
   .I5(level3_in[1067])
);

LUT6 #(
   .INIT(64'h1905620419056204)  
) LUT6_inst9250 (
   .O(to_level2[178]),
   .I0(level3_in[1068]),
   .I1(level3_in[1069]),
   .I2(level3_in[1070]),
   .I3(level3_in[1071]),
   .I4(level3_in[1072]),
   .I5(level3_in[1073])
);

LUT6 #(
   .INIT(64'hf77f577ef77f577e)  
) LUT6_inst9251 (
   .O(to_level2[179]),
   .I0(level3_in[1074]),
   .I1(level3_in[1075]),
   .I2(level3_in[1076]),
   .I3(level3_in[1077]),
   .I4(level3_in[1078]),
   .I5(level3_in[1079])
);

LUT6 #(
   .INIT(64'h0b7a08550b7a0855)  
) LUT6_inst9252 (
   .O(to_level2[180]),
   .I0(level3_in[1080]),
   .I1(level3_in[1081]),
   .I2(level3_in[1082]),
   .I3(level3_in[1083]),
   .I4(level3_in[1084]),
   .I5(level3_in[1085])
);

LUT6 #(
   .INIT(64'h6434187c6434187c)  
) LUT6_inst9253 (
   .O(to_level2[181]),
   .I0(level3_in[1086]),
   .I1(level3_in[1087]),
   .I2(level3_in[1088]),
   .I3(level3_in[1089]),
   .I4(level3_in[1090]),
   .I5(level3_in[1091])
);

LUT6 #(
   .INIT(64'hf7a0ce41f7a0ce41)  
) LUT6_inst9254 (
   .O(to_level2[182]),
   .I0(level3_in[1092]),
   .I1(level3_in[1093]),
   .I2(level3_in[1094]),
   .I3(level3_in[1095]),
   .I4(level3_in[1096]),
   .I5(level3_in[1097])
);

LUT6 #(
   .INIT(64'hc6fd1362c6fd1362)  
) LUT6_inst9255 (
   .O(to_level2[183]),
   .I0(level3_in[1098]),
   .I1(level3_in[1099]),
   .I2(level3_in[1100]),
   .I3(level3_in[1101]),
   .I4(level3_in[1102]),
   .I5(level3_in[1103])
);

LUT6 #(
   .INIT(64'h4a1fffeb4a1fffeb)  
) LUT6_inst9256 (
   .O(to_level2[184]),
   .I0(level3_in[1104]),
   .I1(level3_in[1105]),
   .I2(level3_in[1106]),
   .I3(level3_in[1107]),
   .I4(level3_in[1108]),
   .I5(level3_in[1109])
);

LUT6 #(
   .INIT(64'h3580e49d3580e49d)  
) LUT6_inst9257 (
   .O(to_level2[185]),
   .I0(level3_in[1110]),
   .I1(level3_in[1111]),
   .I2(level3_in[1112]),
   .I3(level3_in[1113]),
   .I4(level3_in[1114]),
   .I5(level3_in[1115])
);

LUT6 #(
   .INIT(64'h30d873f830d873f8)  
) LUT6_inst9258 (
   .O(to_level2[186]),
   .I0(level3_in[1116]),
   .I1(level3_in[1117]),
   .I2(level3_in[1118]),
   .I3(level3_in[1119]),
   .I4(level3_in[1120]),
   .I5(level3_in[1121])
);

LUT6 #(
   .INIT(64'hcbe2ee72cbe2ee72)  
) LUT6_inst9259 (
   .O(to_level2[187]),
   .I0(level3_in[1122]),
   .I1(level3_in[1123]),
   .I2(level3_in[1124]),
   .I3(level3_in[1125]),
   .I4(level3_in[1126]),
   .I5(level3_in[1127])
);

LUT6 #(
   .INIT(64'h348c09d0348c09d0)  
) LUT6_inst9260 (
   .O(to_level2[188]),
   .I0(level3_in[1128]),
   .I1(level3_in[1129]),
   .I2(level3_in[1130]),
   .I3(level3_in[1131]),
   .I4(level3_in[1132]),
   .I5(level3_in[1133])
);

LUT6 #(
   .INIT(64'hab3b589aab3b589a)  
) LUT6_inst9261 (
   .O(to_level2[189]),
   .I0(level3_in[1134]),
   .I1(level3_in[1135]),
   .I2(level3_in[1136]),
   .I3(level3_in[1137]),
   .I4(level3_in[1138]),
   .I5(level3_in[1139])
);

LUT6 #(
   .INIT(64'hb99481a3b99481a3)  
) LUT6_inst9262 (
   .O(to_level2[190]),
   .I0(level3_in[1140]),
   .I1(level3_in[1141]),
   .I2(level3_in[1142]),
   .I3(level3_in[1143]),
   .I4(level3_in[1144]),
   .I5(level3_in[1145])
);

LUT6 #(
   .INIT(64'h5be37a0e5be37a0e)  
) LUT6_inst9263 (
   .O(to_level2[191]),
   .I0(level3_in[1146]),
   .I1(level3_in[1147]),
   .I2(level3_in[1148]),
   .I3(level3_in[1149]),
   .I4(level3_in[1150]),
   .I5(level3_in[1151])
);

LUT6 #(
   .INIT(64'hbe73c5a2be73c5a2)  
) LUT6_inst9264 (
   .O(to_level2[192]),
   .I0(level3_in[1152]),
   .I1(level3_in[1153]),
   .I2(level3_in[1154]),
   .I3(level3_in[1155]),
   .I4(level3_in[1156]),
   .I5(level3_in[1157])
);

LUT6 #(
   .INIT(64'hae1dc14eae1dc14e)  
) LUT6_inst9265 (
   .O(to_level2[193]),
   .I0(level3_in[1158]),
   .I1(level3_in[1159]),
   .I2(level3_in[1160]),
   .I3(level3_in[1161]),
   .I4(level3_in[1162]),
   .I5(level3_in[1163])
);

LUT6 #(
   .INIT(64'h8156d6df8156d6df)  
) LUT6_inst9266 (
   .O(to_level2[194]),
   .I0(level3_in[1164]),
   .I1(level3_in[1165]),
   .I2(level3_in[1166]),
   .I3(level3_in[1167]),
   .I4(level3_in[1168]),
   .I5(level3_in[1169])
);

LUT6 #(
   .INIT(64'h002f1e7d002f1e7d)  
) LUT6_inst9267 (
   .O(to_level2[195]),
   .I0(level3_in[1170]),
   .I1(level3_in[1171]),
   .I2(level3_in[1172]),
   .I3(level3_in[1173]),
   .I4(level3_in[1174]),
   .I5(level3_in[1175])
);

LUT6 #(
   .INIT(64'h13e633b113e633b1)  
) LUT6_inst9268 (
   .O(to_level2[196]),
   .I0(level3_in[1176]),
   .I1(level3_in[1177]),
   .I2(level3_in[1178]),
   .I3(level3_in[1179]),
   .I4(level3_in[1180]),
   .I5(level3_in[1181])
);

LUT6 #(
   .INIT(64'h5d7c7c695d7c7c69)  
) LUT6_inst9269 (
   .O(to_level2[197]),
   .I0(level3_in[1182]),
   .I1(level3_in[1183]),
   .I2(level3_in[1184]),
   .I3(level3_in[1185]),
   .I4(level3_in[1186]),
   .I5(level3_in[1187])
);

LUT6 #(
   .INIT(64'hf2ddc2d1f2ddc2d1)  
) LUT6_inst9270 (
   .O(to_level2[198]),
   .I0(level3_in[1188]),
   .I1(level3_in[1189]),
   .I2(level3_in[1190]),
   .I3(level3_in[1191]),
   .I4(level3_in[1192]),
   .I5(level3_in[1193])
);

LUT6 #(
   .INIT(64'h6e12bed86e12bed8)  
) LUT6_inst9271 (
   .O(to_level2[199]),
   .I0(level3_in[1194]),
   .I1(level3_in[1195]),
   .I2(level3_in[1196]),
   .I3(level3_in[1197]),
   .I4(level3_in[1198]),
   .I5(level3_in[1199])
);

LUT6 #(
   .INIT(64'ha6521053a6521053)  
) LUT6_inst9272 (
   .O(to_level2[200]),
   .I0(level3_in[1200]),
   .I1(level3_in[1201]),
   .I2(level3_in[1202]),
   .I3(level3_in[1203]),
   .I4(level3_in[1204]),
   .I5(level3_in[1205])
);

LUT6 #(
   .INIT(64'he11c2680e11c2680)  
) LUT6_inst9273 (
   .O(to_level2[201]),
   .I0(level3_in[1206]),
   .I1(level3_in[1207]),
   .I2(level3_in[1208]),
   .I3(level3_in[1209]),
   .I4(level3_in[1210]),
   .I5(level3_in[1211])
);

LUT6 #(
   .INIT(64'h6a3465e06a3465e0)  
) LUT6_inst9274 (
   .O(to_level2[202]),
   .I0(level3_in[1212]),
   .I1(level3_in[1213]),
   .I2(level3_in[1214]),
   .I3(level3_in[1215]),
   .I4(level3_in[1216]),
   .I5(level3_in[1217])
);

LUT6 #(
   .INIT(64'h6395015f6395015f)  
) LUT6_inst9275 (
   .O(to_level2[203]),
   .I0(level3_in[1218]),
   .I1(level3_in[1219]),
   .I2(level3_in[1220]),
   .I3(level3_in[1221]),
   .I4(level3_in[1222]),
   .I5(level3_in[1223])
);

LUT6 #(
   .INIT(64'hd5b1dfc1d5b1dfc1)  
) LUT6_inst9276 (
   .O(to_level2[204]),
   .I0(level3_in[1224]),
   .I1(level3_in[1225]),
   .I2(level3_in[1226]),
   .I3(level3_in[1227]),
   .I4(level3_in[1228]),
   .I5(level3_in[1229])
);

LUT6 #(
   .INIT(64'hba0b5e5bba0b5e5b)  
) LUT6_inst9277 (
   .O(to_level2[205]),
   .I0(level3_in[1230]),
   .I1(level3_in[1231]),
   .I2(level3_in[1232]),
   .I3(level3_in[1233]),
   .I4(level3_in[1234]),
   .I5(level3_in[1235])
);

LUT6 #(
   .INIT(64'h74047f2774047f27)  
) LUT6_inst9278 (
   .O(to_level2[206]),
   .I0(level3_in[1236]),
   .I1(level3_in[1237]),
   .I2(level3_in[1238]),
   .I3(level3_in[1239]),
   .I4(level3_in[1240]),
   .I5(level3_in[1241])
);

LUT6 #(
   .INIT(64'he20d3d05e20d3d05)  
) LUT6_inst9279 (
   .O(to_level2[207]),
   .I0(level3_in[1242]),
   .I1(level3_in[1243]),
   .I2(level3_in[1244]),
   .I3(level3_in[1245]),
   .I4(level3_in[1246]),
   .I5(level3_in[1247])
);

LUT6 #(
   .INIT(64'h453a8f19453a8f19)  
) LUT6_inst9280 (
   .O(to_level2[208]),
   .I0(level3_in[1248]),
   .I1(level3_in[1249]),
   .I2(level3_in[1250]),
   .I3(level3_in[1251]),
   .I4(level3_in[1252]),
   .I5(level3_in[1253])
);

LUT6 #(
   .INIT(64'h63d3034863d30348)  
) LUT6_inst9281 (
   .O(to_level2[209]),
   .I0(level3_in[1254]),
   .I1(level3_in[1255]),
   .I2(level3_in[1256]),
   .I3(level3_in[1257]),
   .I4(level3_in[1258]),
   .I5(level3_in[1259])
);

LUT6 #(
   .INIT(64'hb05161b8b05161b8)  
) LUT6_inst9282 (
   .O(to_level2[210]),
   .I0(level3_in[1260]),
   .I1(level3_in[1261]),
   .I2(level3_in[1262]),
   .I3(level3_in[1263]),
   .I4(level3_in[1264]),
   .I5(level3_in[1265])
);

LUT6 #(
   .INIT(64'h1b1b5ab11b1b5ab1)  
) LUT6_inst9283 (
   .O(to_level2[211]),
   .I0(level3_in[1266]),
   .I1(level3_in[1267]),
   .I2(level3_in[1268]),
   .I3(level3_in[1269]),
   .I4(level3_in[1270]),
   .I5(level3_in[1271])
);

LUT6 #(
   .INIT(64'hd39fe26fd39fe26f)  
) LUT6_inst9284 (
   .O(to_level2[212]),
   .I0(level3_in[1272]),
   .I1(level3_in[1273]),
   .I2(level3_in[1274]),
   .I3(level3_in[1275]),
   .I4(level3_in[1276]),
   .I5(level3_in[1277])
);

LUT6 #(
   .INIT(64'hac6f15a9ac6f15a9)  
) LUT6_inst9285 (
   .O(to_level2[213]),
   .I0(level3_in[1278]),
   .I1(level3_in[1279]),
   .I2(level3_in[1280]),
   .I3(level3_in[1281]),
   .I4(level3_in[1282]),
   .I5(level3_in[1283])
);

LUT6 #(
   .INIT(64'h388c4c98388c4c98)  
) LUT6_inst9286 (
   .O(to_level2[214]),
   .I0(level3_in[1284]),
   .I1(level3_in[1285]),
   .I2(level3_in[1286]),
   .I3(level3_in[1287]),
   .I4(level3_in[1288]),
   .I5(level3_in[1289])
);

LUT6 #(
   .INIT(64'h42efdf5f42efdf5f)  
) LUT6_inst9287 (
   .O(to_level2[215]),
   .I0(level3_in[1290]),
   .I1(level3_in[1291]),
   .I2(level3_in[1292]),
   .I3(level3_in[1293]),
   .I4(level3_in[1294]),
   .I5(level3_in[1295])
);
////////////// level 2 starts below:/n
LUT6 #(
   .INIT(64'h65ff5a8a65ff5a8a)  
) LUT6_inst9288 (
   .O(to_level1[0]),
   .I0(level2_in[0]),
   .I1(level2_in[1]),
   .I2(level2_in[2]),
   .I3(level2_in[3]),
   .I4(level2_in[4]),
   .I5(level2_in[5])
);

LUT6 #(
   .INIT(64'h4f00d2d44f00d2d4)  
) LUT6_inst9289 (
   .O(to_level1[1]),
   .I0(level2_in[6]),
   .I1(level2_in[7]),
   .I2(level2_in[8]),
   .I3(level2_in[9]),
   .I4(level2_in[10]),
   .I5(level2_in[11])
);

LUT6 #(
   .INIT(64'hef53b3a0ef53b3a0)  
) LUT6_inst9290 (
   .O(to_level1[2]),
   .I0(level2_in[12]),
   .I1(level2_in[13]),
   .I2(level2_in[14]),
   .I3(level2_in[15]),
   .I4(level2_in[16]),
   .I5(level2_in[17])
);

LUT6 #(
   .INIT(64'he6021481e6021481)  
) LUT6_inst9291 (
   .O(to_level1[3]),
   .I0(level2_in[18]),
   .I1(level2_in[19]),
   .I2(level2_in[20]),
   .I3(level2_in[21]),
   .I4(level2_in[22]),
   .I5(level2_in[23])
);

LUT6 #(
   .INIT(64'h2ac6d8552ac6d855)  
) LUT6_inst9292 (
   .O(to_level1[4]),
   .I0(level2_in[24]),
   .I1(level2_in[25]),
   .I2(level2_in[26]),
   .I3(level2_in[27]),
   .I4(level2_in[28]),
   .I5(level2_in[29])
);

LUT6 #(
   .INIT(64'h617a7cf5617a7cf5)  
) LUT6_inst9293 (
   .O(to_level1[5]),
   .I0(level2_in[30]),
   .I1(level2_in[31]),
   .I2(level2_in[32]),
   .I3(level2_in[33]),
   .I4(level2_in[34]),
   .I5(level2_in[35])
);

LUT6 #(
   .INIT(64'hf01028aef01028ae)  
) LUT6_inst9294 (
   .O(to_level1[6]),
   .I0(level2_in[36]),
   .I1(level2_in[37]),
   .I2(level2_in[38]),
   .I3(level2_in[39]),
   .I4(level2_in[40]),
   .I5(level2_in[41])
);

LUT6 #(
   .INIT(64'h8e4cf10b8e4cf10b)  
) LUT6_inst9295 (
   .O(to_level1[7]),
   .I0(level2_in[42]),
   .I1(level2_in[43]),
   .I2(level2_in[44]),
   .I3(level2_in[45]),
   .I4(level2_in[46]),
   .I5(level2_in[47])
);

LUT6 #(
   .INIT(64'h4afd20924afd2092)  
) LUT6_inst9296 (
   .O(to_level1[8]),
   .I0(level2_in[48]),
   .I1(level2_in[49]),
   .I2(level2_in[50]),
   .I3(level2_in[51]),
   .I4(level2_in[52]),
   .I5(level2_in[53])
);

LUT6 #(
   .INIT(64'h2bd8a31a2bd8a31a)  
) LUT6_inst9297 (
   .O(to_level1[9]),
   .I0(level2_in[54]),
   .I1(level2_in[55]),
   .I2(level2_in[56]),
   .I3(level2_in[57]),
   .I4(level2_in[58]),
   .I5(level2_in[59])
);

LUT6 #(
   .INIT(64'hbe499f46be499f46)  
) LUT6_inst9298 (
   .O(to_level1[10]),
   .I0(level2_in[60]),
   .I1(level2_in[61]),
   .I2(level2_in[62]),
   .I3(level2_in[63]),
   .I4(level2_in[64]),
   .I5(level2_in[65])
);

LUT6 #(
   .INIT(64'hea11f148ea11f148)  
) LUT6_inst9299 (
   .O(to_level1[11]),
   .I0(level2_in[66]),
   .I1(level2_in[67]),
   .I2(level2_in[68]),
   .I3(level2_in[69]),
   .I4(level2_in[70]),
   .I5(level2_in[71])
);

LUT6 #(
   .INIT(64'h44e884f544e884f5)  
) LUT6_inst9300 (
   .O(to_level1[12]),
   .I0(level2_in[72]),
   .I1(level2_in[73]),
   .I2(level2_in[74]),
   .I3(level2_in[75]),
   .I4(level2_in[76]),
   .I5(level2_in[77])
);

LUT6 #(
   .INIT(64'he1b6c859e1b6c859)  
) LUT6_inst9301 (
   .O(to_level1[13]),
   .I0(level2_in[78]),
   .I1(level2_in[79]),
   .I2(level2_in[80]),
   .I3(level2_in[81]),
   .I4(level2_in[82]),
   .I5(level2_in[83])
);

LUT6 #(
   .INIT(64'hc4f2a92dc4f2a92d)  
) LUT6_inst9302 (
   .O(to_level1[14]),
   .I0(level2_in[84]),
   .I1(level2_in[85]),
   .I2(level2_in[86]),
   .I3(level2_in[87]),
   .I4(level2_in[88]),
   .I5(level2_in[89])
);

LUT6 #(
   .INIT(64'h02306cd602306cd6)  
) LUT6_inst9303 (
   .O(to_level1[15]),
   .I0(level2_in[90]),
   .I1(level2_in[91]),
   .I2(level2_in[92]),
   .I3(level2_in[93]),
   .I4(level2_in[94]),
   .I5(level2_in[95])
);

LUT6 #(
   .INIT(64'hbf3919f7bf3919f7)  
) LUT6_inst9304 (
   .O(to_level1[16]),
   .I0(level2_in[96]),
   .I1(level2_in[97]),
   .I2(level2_in[98]),
   .I3(level2_in[99]),
   .I4(level2_in[100]),
   .I5(level2_in[101])
);

LUT6 #(
   .INIT(64'h1118ee791118ee79)  
) LUT6_inst9305 (
   .O(to_level1[17]),
   .I0(level2_in[102]),
   .I1(level2_in[103]),
   .I2(level2_in[104]),
   .I3(level2_in[105]),
   .I4(level2_in[106]),
   .I5(level2_in[107])
);

LUT6 #(
   .INIT(64'hb899ccd0b899ccd0)  
) LUT6_inst9306 (
   .O(to_level1[18]),
   .I0(level2_in[108]),
   .I1(level2_in[109]),
   .I2(level2_in[110]),
   .I3(level2_in[111]),
   .I4(level2_in[112]),
   .I5(level2_in[113])
);

LUT6 #(
   .INIT(64'he5c60c06e5c60c06)  
) LUT6_inst9307 (
   .O(to_level1[19]),
   .I0(level2_in[114]),
   .I1(level2_in[115]),
   .I2(level2_in[116]),
   .I3(level2_in[117]),
   .I4(level2_in[118]),
   .I5(level2_in[119])
);

LUT6 #(
   .INIT(64'h5e0d72065e0d7206)  
) LUT6_inst9308 (
   .O(to_level1[20]),
   .I0(level2_in[120]),
   .I1(level2_in[121]),
   .I2(level2_in[122]),
   .I3(level2_in[123]),
   .I4(level2_in[124]),
   .I5(level2_in[125])
);

LUT6 #(
   .INIT(64'h7e34a6677e34a667)  
) LUT6_inst9309 (
   .O(to_level1[21]),
   .I0(level2_in[126]),
   .I1(level2_in[127]),
   .I2(level2_in[128]),
   .I3(level2_in[129]),
   .I4(level2_in[130]),
   .I5(level2_in[131])
);

LUT6 #(
   .INIT(64'h560becaf560becaf)  
) LUT6_inst9310 (
   .O(to_level1[22]),
   .I0(level2_in[132]),
   .I1(level2_in[133]),
   .I2(level2_in[134]),
   .I3(level2_in[135]),
   .I4(level2_in[136]),
   .I5(level2_in[137])
);

LUT6 #(
   .INIT(64'hde5d8c12de5d8c12)  
) LUT6_inst9311 (
   .O(to_level1[23]),
   .I0(level2_in[138]),
   .I1(level2_in[139]),
   .I2(level2_in[140]),
   .I3(level2_in[141]),
   .I4(level2_in[142]),
   .I5(level2_in[143])
);

LUT6 #(
   .INIT(64'hf8fff495f8fff495)  
) LUT6_inst9312 (
   .O(to_level1[24]),
   .I0(level2_in[144]),
   .I1(level2_in[145]),
   .I2(level2_in[146]),
   .I3(level2_in[147]),
   .I4(level2_in[148]),
   .I5(level2_in[149])
);

LUT6 #(
   .INIT(64'ha6e684d5a6e684d5)  
) LUT6_inst9313 (
   .O(to_level1[25]),
   .I0(level2_in[150]),
   .I1(level2_in[151]),
   .I2(level2_in[152]),
   .I3(level2_in[153]),
   .I4(level2_in[154]),
   .I5(level2_in[155])
);

LUT6 #(
   .INIT(64'hb462adfeb462adfe)  
) LUT6_inst9314 (
   .O(to_level1[26]),
   .I0(level2_in[156]),
   .I1(level2_in[157]),
   .I2(level2_in[158]),
   .I3(level2_in[159]),
   .I4(level2_in[160]),
   .I5(level2_in[161])
);

LUT6 #(
   .INIT(64'h1eeaf7331eeaf733)  
) LUT6_inst9315 (
   .O(to_level1[27]),
   .I0(level2_in[162]),
   .I1(level2_in[163]),
   .I2(level2_in[164]),
   .I3(level2_in[165]),
   .I4(level2_in[166]),
   .I5(level2_in[167])
);

LUT6 #(
   .INIT(64'hbff585eabff585ea)  
) LUT6_inst9316 (
   .O(to_level1[28]),
   .I0(level2_in[168]),
   .I1(level2_in[169]),
   .I2(level2_in[170]),
   .I3(level2_in[171]),
   .I4(level2_in[172]),
   .I5(level2_in[173])
);

LUT6 #(
   .INIT(64'hdf4d6b59df4d6b59)  
) LUT6_inst9317 (
   .O(to_level1[29]),
   .I0(level2_in[174]),
   .I1(level2_in[175]),
   .I2(level2_in[176]),
   .I3(level2_in[177]),
   .I4(level2_in[178]),
   .I5(level2_in[179])
);

LUT6 #(
   .INIT(64'hdf7066f7df7066f7)  
) LUT6_inst9318 (
   .O(to_level1[30]),
   .I0(level2_in[180]),
   .I1(level2_in[181]),
   .I2(level2_in[182]),
   .I3(level2_in[183]),
   .I4(level2_in[184]),
   .I5(level2_in[185])
);

LUT6 #(
   .INIT(64'h5fcf397b5fcf397b)  
) LUT6_inst9319 (
   .O(to_level1[31]),
   .I0(level2_in[186]),
   .I1(level2_in[187]),
   .I2(level2_in[188]),
   .I3(level2_in[189]),
   .I4(level2_in[190]),
   .I5(level2_in[191])
);

LUT6 #(
   .INIT(64'hcf44ca21cf44ca21)  
) LUT6_inst9320 (
   .O(to_level1[32]),
   .I0(level2_in[192]),
   .I1(level2_in[193]),
   .I2(level2_in[194]),
   .I3(level2_in[195]),
   .I4(level2_in[196]),
   .I5(level2_in[197])
);

LUT6 #(
   .INIT(64'hf7001e8ef7001e8e)  
) LUT6_inst9321 (
   .O(to_level1[33]),
   .I0(level2_in[198]),
   .I1(level2_in[199]),
   .I2(level2_in[200]),
   .I3(level2_in[201]),
   .I4(level2_in[202]),
   .I5(level2_in[203])
);

LUT6 #(
   .INIT(64'h1e390ce71e390ce7)  
) LUT6_inst9322 (
   .O(to_level1[34]),
   .I0(level2_in[204]),
   .I1(level2_in[205]),
   .I2(level2_in[206]),
   .I3(level2_in[207]),
   .I4(level2_in[208]),
   .I5(level2_in[209])
);

LUT6 #(
   .INIT(64'h23cbcedf23cbcedf)  
) LUT6_inst9323 (
   .O(to_level1[35]),
   .I0(level2_in[210]),
   .I1(level2_in[211]),
   .I2(level2_in[212]),
   .I3(level2_in[213]),
   .I4(level2_in[214]),
   .I5(level2_in[215])
);
////////////// level 1 starts below:/n
LUT6 #(
   .INIT(64'h78ba1a6a78ba1a6a)  
) LUT6_inst9324 (
   .O(to_level0[0]),
   .I0(level1_in[0]),
   .I1(level1_in[1]),
   .I2(level1_in[2]),
   .I3(level1_in[3]),
   .I4(level1_in[4]),
   .I5(level1_in[5])
);

LUT6 #(
   .INIT(64'h6503c3c16503c3c1)  
) LUT6_inst9325 (
   .O(to_level0[1]),
   .I0(level1_in[6]),
   .I1(level1_in[7]),
   .I2(level1_in[8]),
   .I3(level1_in[9]),
   .I4(level1_in[10]),
   .I5(level1_in[11])
);

LUT6 #(
   .INIT(64'hd01a25a1d01a25a1)  
) LUT6_inst9326 (
   .O(to_level0[2]),
   .I0(level1_in[12]),
   .I1(level1_in[13]),
   .I2(level1_in[14]),
   .I3(level1_in[15]),
   .I4(level1_in[16]),
   .I5(level1_in[17])
);

LUT6 #(
   .INIT(64'h751ac337751ac337)  
) LUT6_inst9327 (
   .O(to_level0[3]),
   .I0(level1_in[18]),
   .I1(level1_in[19]),
   .I2(level1_in[20]),
   .I3(level1_in[21]),
   .I4(level1_in[22]),
   .I5(level1_in[23])
);

LUT6 #(
   .INIT(64'h67735aa867735aa8)  
) LUT6_inst9328 (
   .O(to_level0[4]),
   .I0(level1_in[24]),
   .I1(level1_in[25]),
   .I2(level1_in[26]),
   .I3(level1_in[27]),
   .I4(level1_in[28]),
   .I5(level1_in[29])
);

LUT6 #(
   .INIT(64'h88b98d7888b98d78)  
) LUT6_inst9329 (
   .O(to_level0[5]),
   .I0(level1_in[30]),
   .I1(level1_in[31]),
   .I2(level1_in[32]),
   .I3(level1_in[33]),
   .I4(level1_in[34]),
   .I5(level1_in[35])
);
////////////// level 0 starts below:/n
LUT6 #(
   .INIT(64'hcb0e1a4acb0e1a4a)  
) LUT6_inst9330 (
   .O(data_out_temp),
   .I0(level0_in[0]),
   .I1(level0_in[1]),
   .I2(level0_in[2]),
   .I3(level0_in[3]),
   .I4(level0_in[4]),
   .I5(level0_in[5])
);

endmodule