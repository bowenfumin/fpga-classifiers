module lut_5level_tree4(
                       input       rx_fifo_clock ,
                       input       rx_fifo_resetn,
                       input       [576:0] data_in,
                       input       data_valid,
                       output      data_out     
                       );
wire    [576:0] InputBits;
wire    gates_1, gates_2, gates_3, gates_4, gates_5, gates_6, gates_7, gates_8, gates_9, gates_10, gates_11, gates_12, gates_13, gates_14, gates_15, gates_16, gates_17, gates_18, gates_19, gates_20, gates_21, gates_22, gates_23, gates_24, gates_25, gates_26, gates_27, gates_28, gates_29, gates_30, gates_31, gates_32, gates_33, gates_34, gates_35, gates_36, gates_37, gates_38, gates_39, gates_40, gates_41, gates_42, gates_43, gates_44, gates_45, gates_46, gates_47, gates_48, gates_49, gates_50, gates_51, gates_52, gates_53, gates_54, gates_55, gates_56, gates_57, gates_58, gates_59, gates_60, gates_61, gates_62, gates_63, gates_64, gates_65, gates_66, gates_67, gates_68, gates_69, gates_70, gates_71, gates_72, gates_73, gates_74, gates_75, gates_76, gates_77, gates_78, gates_79, gates_80, gates_81, gates_82, gates_83, gates_84, gates_85, gates_86, gates_87, gates_88, gates_89, gates_90, gates_91, gates_92, gates_93, gates_94, gates_95, gates_96, gates_97, gates_98, gates_99, gates_100, gates_101, gates_102, gates_103, gates_104, gates_105, gates_106, gates_107, gates_108, gates_109, gates_110, gates_111, gates_112, gates_113, gates_114, gates_115, gates_116, gates_117, gates_118, gates_119, gates_120, gates_121, gates_122, gates_123, gates_124, gates_125, gates_126, gates_127, gates_128, gates_129, gates_130, gates_131, gates_132, gates_133, gates_134, gates_135, gates_136, gates_137, gates_138, gates_139, gates_140, gates_141, gates_142, gates_143, gates_144, gates_145, gates_146, gates_147, gates_148, gates_149, gates_150, gates_151, gates_152, gates_153, gates_154, gates_155, gates_156, gates_157, gates_158, gates_159, gates_160, gates_161, gates_162, gates_163, gates_164, gates_165, gates_166, gates_167, gates_168, gates_169, gates_170, gates_171, gates_172, gates_173, gates_174, gates_175, gates_176, gates_177, gates_178, gates_179, gates_180, gates_181, gates_182, gates_183, gates_184, gates_185, gates_186, gates_187, gates_188, gates_189, gates_190, gates_191, gates_192, gates_193, gates_194, gates_195, gates_196, gates_197, gates_198, gates_199, gates_200, gates_201, gates_202, gates_203, gates_204, gates_205, gates_206, gates_207, gates_208, gates_209, gates_210, gates_211, gates_212, gates_213, gates_214, gates_215, gates_216, gates_217, gates_218, gates_219, gates_220, gates_221, gates_222, gates_223, gates_224, gates_225, gates_226, gates_227, gates_228, gates_229, gates_230, gates_231, gates_232, gates_233, gates_234, gates_235, gates_236, gates_237, gates_238, gates_239, gates_240, gates_241, gates_242, gates_243, gates_244, gates_245, gates_246, gates_247, gates_248, gates_249, gates_250, gates_251, gates_252, gates_253, gates_254, gates_255, gates_256, gates_257, gates_258, gates_259, gates_260, gates_261, gates_262, gates_263, gates_264, gates_265, gates_266, gates_267, gates_268, gates_269, gates_270, gates_271, gates_272, gates_273, gates_274, gates_275, gates_276, gates_277, gates_278, gates_279, gates_280, gates_281, gates_282, gates_283, gates_284, gates_285, gates_286, gates_287, gates_288, gates_289, gates_290, gates_291, gates_292, gates_293, gates_294, gates_295, gates_296, gates_297, gates_298, gates_299, gates_300, gates_301, gates_302, gates_303, gates_304, gates_305, gates_306, gates_307, gates_308, gates_309, gates_310, gates_311, gates_312, gates_313, gates_314, gates_315, gates_316, gates_317, gates_318, gates_319, gates_320, gates_321, gates_322, gates_323, gates_324, gates_325, gates_326, gates_327, gates_328, gates_329, gates_330, gates_331, gates_332, gates_333, gates_334, gates_335, gates_336, gates_337, gates_338, gates_339, gates_340, gates_341, gates_342, gates_343, gates_344, gates_345, gates_346, gates_347, gates_348, gates_349, gates_350, gates_351, gates_352, gates_353, gates_354, gates_355, gates_356, gates_357, gates_358, gates_359, gates_360, gates_361, gates_362, gates_363, gates_364, gates_365, gates_366, gates_367, gates_368, gates_369, gates_370, gates_371, gates_372, gates_373, gates_374, gates_375, gates_376, gates_377, gates_378, gates_379, gates_380, gates_381, gates_382, gates_383, gates_384, gates_385, gates_386, gates_387, gates_388, gates_389, gates_390, gates_391, gates_392, gates_393, gates_394, gates_395, gates_396, gates_397, gates_398, gates_399, gates_400, gates_401, gates_402, gates_403, gates_404, gates_405, gates_406, gates_407, gates_408, gates_409, gates_410, gates_411, gates_412, gates_413, gates_414, gates_415, gates_416, gates_417, gates_418, gates_419, gates_420, gates_421, gates_422, gates_423, gates_424, gates_425, gates_426, gates_427, gates_428, gates_429, gates_430, gates_431, gates_432, gates_433, gates_434, gates_435, gates_436, gates_437, gates_438, gates_439, gates_440, gates_441, gates_442, gates_443, gates_444, gates_445, gates_446, gates_447, gates_448, gates_449, gates_450, gates_451, gates_452, gates_453, gates_454, gates_455, gates_456, gates_457, gates_458, gates_459, gates_460, gates_461, gates_462, gates_463, gates_464, gates_465, gates_466, gates_467, gates_468, gates_469, gates_470, gates_471, gates_472, gates_473, gates_474, gates_475, gates_476, gates_477, gates_478, gates_479, gates_480, gates_481, gates_482, gates_483, gates_484, gates_485, gates_486, gates_487, gates_488, gates_489, gates_490, gates_491, gates_492, gates_493, gates_494, gates_495, gates_496, gates_497, gates_498, gates_499, gates_500, gates_501, gates_502, gates_503, gates_504, gates_505, gates_506, gates_507, gates_508, gates_509, gates_510, gates_511, gates_512, gates_513, gates_514, gates_515, gates_516, gates_517, gates_518, gates_519, gates_520, gates_521, gates_522, gates_523, gates_524, gates_525, gates_526, gates_527, gates_528, gates_529, gates_530, gates_531, gates_532, gates_533, gates_534, gates_535, gates_536, gates_537, gates_538, gates_539, gates_540, gates_541, gates_542, gates_543, gates_544, gates_545, gates_546, gates_547, gates_548, gates_549, gates_550, gates_551, gates_552, gates_553, gates_554, gates_555, gates_556, gates_557, gates_558, gates_559, gates_560, gates_561, gates_562, gates_563, gates_564, gates_565, gates_566, gates_567, gates_568, gates_569, gates_570, gates_571, gates_572, gates_573, gates_574, gates_575, gates_576, gates_577, gates_578, gates_579, gates_580, gates_581, gates_582, gates_583, gates_584, gates_585, gates_586, gates_587, gates_588, gates_589, gates_590, gates_591, gates_592, gates_593, gates_594, gates_595, gates_596, gates_597, gates_598, gates_599, gates_600, gates_601, gates_602, gates_603, gates_604, gates_605, gates_606, gates_607, gates_608, gates_609, gates_610, gates_611, gates_612, gates_613, gates_614, gates_615, gates_616, gates_617, gates_618, gates_619, gates_620, gates_621, gates_622, gates_623, gates_624, gates_625, gates_626, gates_627, gates_628, gates_629, gates_630, gates_631, gates_632, gates_633, gates_634, gates_635, gates_636, gates_637, gates_638, gates_639, gates_640, gates_641, gates_642, gates_643, gates_644, gates_645, gates_646, gates_647, gates_648, gates_649, gates_650, gates_651, gates_652, gates_653, gates_654, gates_655, gates_656, gates_657, gates_658, gates_659, gates_660, gates_661, gates_662, gates_663, gates_664, gates_665, gates_666, gates_667, gates_668, gates_669, gates_670, gates_671, gates_672, gates_673, gates_674, gates_675, gates_676, gates_677, gates_678, gates_679, gates_680, gates_681, gates_682, gates_683, gates_684, gates_685, gates_686, gates_687, gates_688, gates_689, gates_690, gates_691, gates_692, gates_693, gates_694, gates_695, gates_696, gates_697, gates_698, gates_699, gates_700, gates_701, gates_702, gates_703, gates_704, gates_705, gates_706, gates_707, gates_708, gates_709, gates_710, gates_711, gates_712, gates_713, gates_714, gates_715, gates_716, gates_717, gates_718, gates_719, gates_720, gates_721, gates_722, gates_723, gates_724, gates_725, gates_726, gates_727, gates_728, gates_729, gates_730, gates_731, gates_732, gates_733, gates_734, gates_735, gates_736, gates_737, gates_738, gates_739, gates_740, gates_741, gates_742, gates_743, gates_744, gates_745, gates_746, gates_747, gates_748, gates_749, gates_750, gates_751, gates_752, gates_753, gates_754, gates_755, gates_756, gates_757, gates_758, gates_759, gates_760, gates_761, gates_762, gates_763, gates_764, gates_765, gates_766, gates_767, gates_768, gates_769, gates_770, gates_771, gates_772, gates_773, gates_774, gates_775, gates_776, gates_777, gates_778, gates_779, gates_780, gates_781, gates_782, gates_783, gates_784, gates_785, gates_786, gates_787, gates_788, gates_789, gates_790, gates_791, gates_792, gates_793, gates_794, gates_795, gates_796, gates_797, gates_798, gates_799, gates_800, gates_801, gates_802, gates_803, gates_804, gates_805, gates_806, gates_807, gates_808, gates_809, gates_810, gates_811, gates_812, gates_813, gates_814, gates_815, gates_816, gates_817, gates_818, gates_819, gates_820, gates_821, gates_822, gates_823, gates_824, gates_825, gates_826, gates_827, gates_828, gates_829, gates_830, gates_831, gates_832, gates_833, gates_834, gates_835, gates_836, gates_837, gates_838, gates_839, gates_840, gates_841, gates_842, gates_843, gates_844, gates_845, gates_846, gates_847, gates_848, gates_849, gates_850, gates_851, gates_852, gates_853, gates_854, gates_855, gates_856, gates_857, gates_858, gates_859, gates_860, gates_861, gates_862, gates_863, gates_864, gates_865, gates_866, gates_867, gates_868, gates_869, gates_870, gates_871, gates_872, gates_873, gates_874, gates_875, gates_876, gates_877, gates_878, gates_879, gates_880, gates_881, gates_882, gates_883, gates_884, gates_885, gates_886, gates_887, gates_888, gates_889, gates_890, gates_891, gates_892, gates_893, gates_894, gates_895, gates_896, gates_897, gates_898, gates_899, gates_900, gates_901, gates_902, gates_903, gates_904, gates_905, gates_906, gates_907, gates_908, gates_909, gates_910, gates_911, gates_912, gates_913, gates_914, gates_915, gates_916, gates_917, gates_918, gates_919, gates_920, gates_921, gates_922, gates_923, gates_924, gates_925, gates_926, gates_927, gates_928, gates_929, gates_930, gates_931, gates_932, gates_933, gates_934, gates_935, gates_936, gates_937, gates_938, gates_939, gates_940, gates_941, gates_942, gates_943, gates_944, gates_945, gates_946, gates_947, gates_948, gates_949, gates_950, gates_951, gates_952, gates_953, gates_954, gates_955, gates_956, gates_957, gates_958, gates_959, gates_960, gates_961, gates_962, gates_963, gates_964, gates_965, gates_966, gates_967, gates_968, gates_969, gates_970, gates_971, gates_972, gates_973, gates_974, gates_975, gates_976, gates_977, gates_978, gates_979, gates_980, gates_981, gates_982, gates_983, gates_984, gates_985, gates_986, gates_987, gates_988, gates_989, gates_990, gates_991, gates_992, gates_993, gates_994, gates_995, gates_996, gates_997, gates_998, gates_999, gates_1000, gates_1001, gates_1002, gates_1003, gates_1004, gates_1005, gates_1006, gates_1007, gates_1008, gates_1009, gates_1010, gates_1011, gates_1012, gates_1013, gates_1014, gates_1015, gates_1016, gates_1017, gates_1018, gates_1019, gates_1020, gates_1021, gates_1022, gates_1023, gates_1024, gates_1025, gates_1026, gates_1027, gates_1028, gates_1029, gates_1030, gates_1031, gates_1032, gates_1033, gates_1034, gates_1035, gates_1036, gates_1037, gates_1038, gates_1039, gates_1040, gates_1041, gates_1042, gates_1043, gates_1044, gates_1045, gates_1046, gates_1047, gates_1048, gates_1049, gates_1050, gates_1051, gates_1052, gates_1053, gates_1054, gates_1055, gates_1056, gates_1057, gates_1058, gates_1059, gates_1060, gates_1061, gates_1062, gates_1063, gates_1064, gates_1065, gates_1066, gates_1067, gates_1068, gates_1069, gates_1070, gates_1071, gates_1072, gates_1073, gates_1074, gates_1075, gates_1076, gates_1077, gates_1078, gates_1079, gates_1080, gates_1081, gates_1082, gates_1083, gates_1084, gates_1085, gates_1086, gates_1087, gates_1088, gates_1089, gates_1090, gates_1091, gates_1092, gates_1093, gates_1094, gates_1095, gates_1096, gates_1097, gates_1098, gates_1099, gates_1100, gates_1101, gates_1102, gates_1103, gates_1104, gates_1105, gates_1106, gates_1107, gates_1108, gates_1109, gates_1110, gates_1111, gates_1112, gates_1113, gates_1114, gates_1115, gates_1116, gates_1117, gates_1118, gates_1119, gates_1120, gates_1121, gates_1122, gates_1123, gates_1124, gates_1125, gates_1126, gates_1127, gates_1128, gates_1129, gates_1130, gates_1131, gates_1132, gates_1133, gates_1134, gates_1135, gates_1136, gates_1137, gates_1138, gates_1139, gates_1140, gates_1141, gates_1142, gates_1143, gates_1144, gates_1145, gates_1146, gates_1147, gates_1148, gates_1149, gates_1150, gates_1151, gates_1152, gates_1153, gates_1154, gates_1155, gates_1156, gates_1157, gates_1158, gates_1159, gates_1160, gates_1161, gates_1162, gates_1163, gates_1164, gates_1165, gates_1166, gates_1167, gates_1168, gates_1169, gates_1170, gates_1171, gates_1172, gates_1173, gates_1174, gates_1175, gates_1176, gates_1177, gates_1178, gates_1179, gates_1180, gates_1181, gates_1182, gates_1183, gates_1184, gates_1185, gates_1186, gates_1187, gates_1188, gates_1189, gates_1190, gates_1191, gates_1192, gates_1193, gates_1194, gates_1195, gates_1196, gates_1197, gates_1198, gates_1199, gates_1200, gates_1201, gates_1202, gates_1203, gates_1204, gates_1205, gates_1206, gates_1207, gates_1208, gates_1209, gates_1210, gates_1211, gates_1212, gates_1213, gates_1214, gates_1215, gates_1216, gates_1217, gates_1218, gates_1219, gates_1220, gates_1221, gates_1222, gates_1223, gates_1224, gates_1225, gates_1226, gates_1227, gates_1228, gates_1229, gates_1230, gates_1231, gates_1232, gates_1233, gates_1234, gates_1235, gates_1236, gates_1237, gates_1238, gates_1239, gates_1240, gates_1241, gates_1242, gates_1243, gates_1244, gates_1245, gates_1246, gates_1247, gates_1248, gates_1249, gates_1250, gates_1251, gates_1252, gates_1253, gates_1254, gates_1255, gates_1256, gates_1257, gates_1258, gates_1259, gates_1260, gates_1261, gates_1262, gates_1263, gates_1264, gates_1265, gates_1266, gates_1267, gates_1268, gates_1269, gates_1270, gates_1271, gates_1272, gates_1273, gates_1274, gates_1275, gates_1276, gates_1277, gates_1278, gates_1279, gates_1280, gates_1281, gates_1282, gates_1283, gates_1284, gates_1285, gates_1286, gates_1287, gates_1288, gates_1289, gates_1290, gates_1291, gates_1292, gates_1293, gates_1294, gates_1295, gates_1296, gates_1297, gates_1298, gates_1299, gates_1300, gates_1301, gates_1302, gates_1303, gates_1304, gates_1305, gates_1306, gates_1307, gates_1308, gates_1309, gates_1310, gates_1311, gates_1312, gates_1313, gates_1314, gates_1315, gates_1316, gates_1317, gates_1318, gates_1319, gates_1320, gates_1321, gates_1322, gates_1323, gates_1324, gates_1325, gates_1326, gates_1327, gates_1328, gates_1329, gates_1330, gates_1331, gates_1332, gates_1333, gates_1334, gates_1335, gates_1336, gates_1337, gates_1338, gates_1339, gates_1340, gates_1341, gates_1342, gates_1343, gates_1344, gates_1345, gates_1346, gates_1347, gates_1348, gates_1349, gates_1350, gates_1351, gates_1352, gates_1353, gates_1354, gates_1355, gates_1356, gates_1357, gates_1358, gates_1359, gates_1360, gates_1361, gates_1362, gates_1363, gates_1364, gates_1365, gates_1366, gates_1367, gates_1368, gates_1369, gates_1370, gates_1371, gates_1372, gates_1373, gates_1374, gates_1375, gates_1376, gates_1377, gates_1378, gates_1379, gates_1380, gates_1381, gates_1382, gates_1383, gates_1384, gates_1385, gates_1386, gates_1387, gates_1388, gates_1389, gates_1390, gates_1391, gates_1392, gates_1393, gates_1394, gates_1395, gates_1396, gates_1397, gates_1398, gates_1399, gates_1400, gates_1401, gates_1402, gates_1403, gates_1404, gates_1405, gates_1406, gates_1407, gates_1408, gates_1409, gates_1410, gates_1411, gates_1412, gates_1413, gates_1414, gates_1415, gates_1416, gates_1417, gates_1418, gates_1419, gates_1420, gates_1421, gates_1422, gates_1423, gates_1424, gates_1425, gates_1426, gates_1427, gates_1428, gates_1429, gates_1430, gates_1431, gates_1432, gates_1433, gates_1434, gates_1435, gates_1436, gates_1437, gates_1438, gates_1439, gates_1440, gates_1441, gates_1442, gates_1443, gates_1444, gates_1445, gates_1446, gates_1447, gates_1448, gates_1449, gates_1450, gates_1451, gates_1452, gates_1453, gates_1454, gates_1455, gates_1456, gates_1457, gates_1458, gates_1459, gates_1460, gates_1461, gates_1462, gates_1463, gates_1464, gates_1465, gates_1466, gates_1467, gates_1468, gates_1469, gates_1470, gates_1471, gates_1472, gates_1473, gates_1474, gates_1475, gates_1476, gates_1477, gates_1478, gates_1479, gates_1480, gates_1481, gates_1482, gates_1483, gates_1484, gates_1485, gates_1486, gates_1487, gates_1488, gates_1489, gates_1490, gates_1491, gates_1492, gates_1493, gates_1494, gates_1495, gates_1496, gates_1497, gates_1498, gates_1499, gates_1500, gates_1501, gates_1502, gates_1503, gates_1504, gates_1505, gates_1506, gates_1507, gates_1508, gates_1509, gates_1510, gates_1511, gates_1512, gates_1513, gates_1514, gates_1515, gates_1516, gates_1517, gates_1518, gates_1519, gates_1520, gates_1521, gates_1522, gates_1523, gates_1524, gates_1525, gates_1526, gates_1527, gates_1528, gates_1529, gates_1530, gates_1531, gates_1532, gates_1533, gates_1534, gates_1535, gates_1536, gates_1537, gates_1538, gates_1539, gates_1540, gates_1541, gates_1542, gates_1543, gates_1544, gates_1545, gates_1546, gates_1547, gates_1548, gates_1549, gates_1550, gates_1551, gates_1552, gates_1553, gates_1554, gates_1555;

assign  InputBits = data_in;
//assign  data_out = data_valid & gates[807];
assign  data_out = data_valid & gates_1422;

LUT6 #(
   .INIT(64'b0111000100000010101111010110010111111000101011000001010111110100)  
) LUT6_1 (
   .O(gates_29),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1110100100011111010101010110101110111001011100011011111000110110)  
) LUT6_2 (
   .O(gates_124),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0101011010001111011001011101010111001001010101110101111000100010)  
) LUT6_3 (
   .O(gates_1412),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0001100000101111100101101101101101110000101100110101101000110011)  
) LUT6_4 (
   .O(gates_780),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0000100110100111000111001010011011101101010110111110000010010100)  
) LUT6_5 (
   .O(gates_1003),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1010000010110100111110011000100110110010010111110000001111100110)  
) LUT6_6 (
   .O(gates_709),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0100010100001001001111100001101100110011011000100101000100010010)  
) LUT6_7 (
   .O(gates_1173),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000110100001111110001110001100111111000110000000110101000111101)  
) LUT6_8 (
   .O(gates_1250),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0011101000011110000011111110101100110100000001011011101100101110)  
) LUT6_9 (
   .O(gates_1415),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0000110001010001110000100111000100101110001000011011100111100011)  
) LUT6_10 (
   .O(gates_86),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0011100100111000010010110100100000101001001010001100100001001111)  
) LUT6_11 (
   .O(gates_76),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b1010101001110000111100110100001111000000101010001110101110000110)  
) LUT6_12 (
   .O(gates_1266),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1111111100010010100110010000111010011001110000100011010101011000)  
) LUT6_13 (
   .O(gates_1051),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0100011100101100001110111011001001101110001001100100101111100001)  
) LUT6_14 (
   .O(gates_1451),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0000010101010100101110000010111011001100110000111010100111111100)  
) LUT6_15 (
   .O(gates_309),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0011100010101100110011010011010001011100000100111100110110000101)  
) LUT6_16 (
   .O(gates_155),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0111100100101110101011001110000010010101010001100100010010001000)  
) LUT6_17 (
   .O(gates_588),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1001010110100011010110110101110001010000011000010100110000010101)  
) LUT6_18 (
   .O(gates_1352),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001000011001010001000001001100110011101101001101111011011110011)  
) LUT6_19 (
   .O(gates_148),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0001011001001011111101110001110000100011101010111000000011111101)  
) LUT6_20 (
   .O(gates_1210),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0110111011101011111110100110000010000110100010100110000101001110)  
) LUT6_21 (
   .O(gates_1153),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1100010000000110111011001001101101101100011001101101111111100111)  
) LUT6_22 (
   .O(gates_205),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1101101100100100101110000011100101000110000011000111111000001110)  
) LUT6_23 (
   .O(gates_527),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100101101101110111101111110101010100110100011110100011001010111)  
) LUT6_24 (
   .O(gates_20),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1110101101011001001011100000011110101010111100010100110100110101)  
) LUT6_25 (
   .O(gates_1334),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1111010001110010100111011101010110100101000101110110011010001101)  
) LUT6_26 (
   .O(gates_160),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1110110101101101100000010010100001011111111101110011000010010111)  
) LUT6_27 (
   .O(gates_606),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1001001111100100100000101100100110100010010100001011101110000010)  
) LUT6_28 (
   .O(gates_1354),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0010111000010111000100110000011111000110111010111100010110011011)  
) LUT6_29 (
   .O(gates_1066),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0011110101000000110110011100101101110110010010100110100011101010)  
) LUT6_30 (
   .O(gates_187),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1111001100110000110101110100110010111001000000011001101100110010)  
) LUT6_31 (
   .O(gates_1127),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1111010101001010110010111001101000010011011011101100010000011000)  
) LUT6_32 (
   .O(gates_80),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1101000000010101111010110001000100100010011100110010110111110001)  
) LUT6_33 (
   .O(gates_854),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010111000111000000110111111111000000100110000001010010011000110)  
) LUT6_34 (
   .O(gates_656),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0011100000001110011101011101101001110111100101000001000001111111)  
) LUT6_35 (
   .O(gates_1247),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1001111110010011111101010110111110001100010010110100010010101110)  
) LUT6_36 (
   .O(gates_1447),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0110011000011100101100110100110000001001111111111000011110101001)  
) LUT6_37 (
   .O(gates_1207),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1111110001001011000010111110011011001000100101110000111001100100)  
) LUT6_38 (
   .O(gates_298),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0101100011110010010001010110101101110101111000111101101000001011)  
) LUT6_39 (
   .O(gates_785),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1110010110000100111100110100111111001010101100010001000110000100)  
) LUT6_40 (
   .O(gates_226),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1101011100010000011001011011111100110011100001101000100011000000)  
) LUT6_41 (
   .O(gates_315),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1011010010100111101110100110111111100001101001101110101001111000)  
) LUT6_42 (
   .O(gates_671),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1010100101000001110111100101001111011110011111101111111111111001)  
) LUT6_43 (
   .O(gates_69),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1001111111001001010001001011001000011100110110000111100100100011)  
) LUT6_44 (
   .O(gates_478),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1011010110011111010011110011100011011101001010001011011010011010)  
) LUT6_45 (
   .O(gates_1100),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1000001110011011011001010100010010010011010111011100111011000111)  
) LUT6_46 (
   .O(gates_1479),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1001011101010001011111001010001001000011100010010011100100100111)  
) LUT6_47 (
   .O(gates_547),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0000011100000010011000110100101101101110110110011010101101001100)  
) LUT6_48 (
   .O(gates_1359),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0011011000011110101100100110010001101110000000101000110110010010)  
) LUT6_49 (
   .O(gates_435),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1110110011011000011110111100001100001100001101010101000110110010)  
) LUT6_50 (
   .O(gates_330),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1001110000000001110110001101010111100111001111110000111110111010)  
) LUT6_51 (
   .O(gates_409),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0110000101111100110111000101011101000101101000000000000100001111)  
) LUT6_52 (
   .O(gates_270),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0100111111010110001101111001110000100111100001011011101010000011)  
) LUT6_53 (
   .O(gates_1436),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1001101101011000010101110000010101100011111000011100100101010111)  
) LUT6_54 (
   .O(gates_1133),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0111010010011101011101011101110011000100011001110100101101110110)  
) LUT6_55 (
   .O(gates_240),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0001111111100101001000110110011010100100010111010111101100111110)  
) LUT6_56 (
   .O(gates_1289),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0100100011110101000110111101110011111100010100101111010011000001)  
) LUT6_57 (
   .O(gates_27),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0110001010000100000011111001000000101110100011011111100001000010)  
) LUT6_58 (
   .O(gates_183),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1100001010000101011011001111011011011001000111101001100000100110)  
) LUT6_59 (
   .O(gates_636),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1000010010110110001101010111100001100001111111011011100101100101)  
) LUT6_60 (
   .O(gates_745),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b1000001111010011001000001100110011010001110111000100001101110001)  
) LUT6_61 (
   .O(gates_1208),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1001000010110100001111101111011111101110000010101111001111110000)  
) LUT6_62 (
   .O(gates_1312),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1101101100010111011010011111011101100000111101000001100001110101)  
) LUT6_63 (
   .O(gates_1272),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0110100011100000010010111001000001101000011111001011101101101011)  
) LUT6_64 (
   .O(gates_1098),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0011011001100111111110110100110000011111001000100101000111100101)  
) LUT6_65 (
   .O(gates_149),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0110111001000111110100101011000010001011101010101011010110111100)  
) LUT6_66 (
   .O(gates_1249),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1111111110111010111101000101101010010011010001001100101000111101)  
) LUT6_67 (
   .O(gates_687),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0111101111000011001001011010000001110001101010011010001101111001)  
) LUT6_68 (
   .O(gates_888),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b1110010110111011011111100111000111010101110010011100001011101000)  
) LUT6_69 (
   .O(gates_874),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0000100100111001110110101101001101110000001111101000010101101010)  
) LUT6_70 (
   .O(gates_649),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0001010000101011011000001100000011000000001101011010000111101110)  
) LUT6_71 (
   .O(gates_1503),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1101100010000011101000100100000110011011000100101111110101111111)  
) LUT6_72 (
   .O(gates_1043),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b1001001111111100001100010010101110100001000111101110010010001001)  
) LUT6_73 (
   .O(gates_1425),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0010111000010001110000010110110011001011011001110100010100100100)  
) LUT6_74 (
   .O(gates_586),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1011011111100110001110000010111101110111000001101010101101010100)  
) LUT6_75 (
   .O(gates_136),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0010001110011101110111101100001010000110111010001111010111000000)  
) LUT6_76 (
   .O(gates_180),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1100100100001110110001000011100011010010101011111000111000010101)  
) LUT6_77 (
   .O(gates_1146),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0101000011001011111011000011111010011001111100101111100001010010)  
) LUT6_78 (
   .O(gates_1472),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0111011000110110111111001001101001101011001010001110100000101101)  
) LUT6_79 (
   .O(gates_530),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0110001100000100100010101011111110000100011011000111111011000111)  
) LUT6_80 (
   .O(gates_998),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0110111001101110111100111001011000010010011011101100111110100010)  
) LUT6_81 (
   .O(gates_456),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0101010000101101010110010110000010110100110110101110011111011010)  
) LUT6_82 (
   .O(gates_246),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1110010100010100001110010010110110010010000110110100101011010101)  
) LUT6_83 (
   .O(gates_233),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b0101011000101100011000100000000010001101011111000111000101000111)  
) LUT6_84 (
   .O(gates_1199),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1001011000110001010010111100100011000000010011101111011110001001)  
) LUT6_85 (
   .O(gates_863),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0001100001101111000110101111010011110010110101010111101000010100)  
) LUT6_86 (
   .O(gates_711),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b1001011010000110110110100111111101100110000110001001000011100101)  
) LUT6_87 (
   .O(gates_1406),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0110001011001000100100001011101000111010110000100011001010111000)  
) LUT6_88 (
   .O(gates_1327),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1101010001111011001100010011100001111000101001001110101110101011)  
) LUT6_89 (
   .O(gates_581),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0101011001010110111101110001100000001100111100101100000101110110)  
) LUT6_90 (
   .O(gates_765),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0011010011110100011000110111100101101011101101111000101011110001)  
) LUT6_91 (
   .O(gates_403),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0111100100000011010111110110010100011011111100000000010000001001)  
) LUT6_92 (
   .O(gates_960),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0101001111001011110100111100111001111011011000001010110111100100)  
) LUT6_93 (
   .O(gates_1530),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0100110111000101101011110011011111110101000101000101000000100101)  
) LUT6_94 (
   .O(gates_554),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1001110010110010000100000101001100000010011011111010010101011010)  
) LUT6_95 (
   .O(gates_1304),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0100001101101111011100110001110010010111110011110010101010111001)  
) LUT6_96 (
   .O(gates_1476),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000010011010001000101000111110001101110100011010000110101100110)  
) LUT6_97 (
   .O(gates_806),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0011010001010100100110011110101110011100011010001001001000011000)  
) LUT6_98 (
   .O(gates_1362),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b1011001001110111100111011001000111000100111010010001110101110110)  
) LUT6_99 (
   .O(gates_1259),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1100010000111010100110110100101000100000010111001010010010100011)  
) LUT6_100 (
   .O(gates_1388),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1001001001000110011000111111011011100001110100000001110101010000)  
) LUT6_101 (
   .O(gates_1209),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1001111001001110011101001011101101011100100111101010010100101110)  
) LUT6_102 (
   .O(gates_1337),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1111110100010101111010101000010101001111011101111111110001011001)  
) LUT6_103 (
   .O(gates_775),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0110100101111110011001111100000100110000001101011110111000111001)  
) LUT6_104 (
   .O(gates_207),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1000110111100000111100110111110100111110111100000110111101100011)  
) LUT6_105 (
   .O(gates_702),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0010000000100011010110010001110110101110100011001010101110110110)  
) LUT6_106 (
   .O(gates_1096),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1000010110011110000101011111001100110100100111000010111001110100)  
) LUT6_107 (
   .O(gates_294),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b1110111001100001010010000111010011100101111100001001011100100011)  
) LUT6_108 (
   .O(gates_1387),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1011101010010111011111101011010101101111011000101000010110000000)  
) LUT6_109 (
   .O(gates_243),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0010100101111001000001001101111011101111100000011001110000010011)  
) LUT6_110 (
   .O(gates_371),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1001111000110000100110110000001100011000001011100100100100111011)  
) LUT6_111 (
   .O(gates_1375),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1110100010101000100111110000111001101100111000111011000011001001)  
) LUT6_112 (
   .O(gates_164),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1101011010111000010100100110111100010100010011000111110010111111)  
) LUT6_113 (
   .O(gates_432),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1000000000011100110000000100101101110010100000111100111001010000)  
) LUT6_114 (
   .O(gates_381),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0111101010011000011010110011101100010000001010001000101101101110)  
) LUT6_115 (
   .O(gates_408),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0110101110000111111110011101110111011011101101011101000010011101)  
) LUT6_116 (
   .O(gates_1302),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0110000011011111001101101011011110000001010100101011110010000101)  
) LUT6_117 (
   .O(gates_912),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1011001111011100001100000000001000001000100001001101111111110100)  
) LUT6_118 (
   .O(gates_555),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1001111011011110111110110011000010011000011011110101010101011101)  
) LUT6_119 (
   .O(gates_261),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0001111111011001000111101111000011000000010110101111011000000110)  
) LUT6_120 (
   .O(gates_523),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0000110000010010001101110010011100010011011000111111001100001101)  
) LUT6_121 (
   .O(gates_971),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1100000000100100010101111111101100101000010001000000101111100101)  
) LUT6_122 (
   .O(gates_147),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0001001011000111000001101010101101111000001111001110100011110111)  
) LUT6_123 (
   .O(gates_55),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0100011010011101101100001000101000101100011100011111000111101010)  
) LUT6_124 (
   .O(gates_917),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0111101000001010000000010110100111110111101110011011111111000010)  
) LUT6_125 (
   .O(gates_12),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0000101011110101111001110001110111010100111000100001001001000001)  
) LUT6_126 (
   .O(gates_582),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0010110011110010000100101000110011100001100101010001100111011010)  
) LUT6_127 (
   .O(gates_499),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1111000010000001010011110100100001011001010011010110100001011110)  
) LUT6_128 (
   .O(gates_166),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1100010010000110101111010101100000000001000111101010101100111101)  
) LUT6_129 (
   .O(gates_119),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1110101101100101111000001100011100001100010111000101101100001011)  
) LUT6_130 (
   .O(gates_116),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1000100101100001101010010111010101011111111101010110111011111001)  
) LUT6_131 (
   .O(gates_313),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1001011111101011111011000110000101001011010100101011110011010000)  
) LUT6_132 (
   .O(gates_672),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b1011101000100001100011000110011110001100111101110010110101111011)  
) LUT6_133 (
   .O(gates_747),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0101101010111011001001001110111011001111110010100011001111100110)  
) LUT6_134 (
   .O(gates_1397),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0100010100001110010111110100010010000010011110011011010111110001)  
) LUT6_135 (
   .O(gates_157),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0110111000110001110001111110110001010011110111110010111111000010)  
) LUT6_136 (
   .O(gates_282),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0100010011101011110001010110101100010100001110001111100111011110)  
) LUT6_137 (
   .O(gates_297),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0100001001000000111100011101000000011110000110101011110000011101)  
) LUT6_138 (
   .O(gates_1507),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1000001100111001000011101101110100001100110011111000011110111000)  
) LUT6_139 (
   .O(gates_61),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0100111101000011110010100100110111111100100011100001010000010000)  
) LUT6_140 (
   .O(gates_993),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0010111100110111010111001111001111011110100000001110010110111000)  
) LUT6_141 (
   .O(gates_1309),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010001111001001001111011110101001011111011011011000101000001111)  
) LUT6_142 (
   .O(gates_673),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1000011100010000001000010111110010111000100110111110000100101111)  
) LUT6_143 (
   .O(gates_1462),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0011010110100111011001101001100110110011100010000011010000000111)  
) LUT6_144 (
   .O(gates_682),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0011011110001101000011100001110111100011101001011110110101000011)  
) LUT6_145 (
   .O(gates_1251),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1011001100110100010100011010110000000011011100100001000011111110)  
) LUT6_146 (
   .O(gates_897),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1111100011011111111000110000110010111101010000110001010001011110)  
) LUT6_147 (
   .O(gates_571),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1011000011110010101101101110110110100001010001110001101111010001)  
) LUT6_148 (
   .O(gates_1411),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b1100101000101010101110011110000010011101110111000000111111010011)  
) LUT6_149 (
   .O(gates_1058),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1100000000100011001000010111101001100011110101111101010110111000)  
) LUT6_150 (
   .O(gates_455),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0000110011110101001001100001001011100101100101000000011110101011)  
) LUT6_151 (
   .O(gates_1267),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1101001110110111000101100101011000111100110111011100110101101000)  
) LUT6_152 (
   .O(gates_319),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0110011100011000011010001100010011101010110100101111010000000000)  
) LUT6_153 (
   .O(gates_884),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0000100110010111000101111101010110111111001111111000001101011110)  
) LUT6_154 (
   .O(gates_263),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1001110100001011111111011000001000010001110100000100001000110111)  
) LUT6_155 (
   .O(gates_1416),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1110000111101111011011110001001111100110111100011111000110101011)  
) LUT6_156 (
   .O(gates_1092),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0100010101010101110001000111110000100001010111110110101000010110)  
) LUT6_157 (
   .O(gates_1294),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0110101011100111101001101101111000110101111010010001100000000000)  
) LUT6_158 (
   .O(gates_1215),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1111101001011011110000000001000100110100000111011000011110100110)  
) LUT6_159 (
   .O(gates_678),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0000001101001000110111011011001100010111111110000101100001001101)  
) LUT6_160 (
   .O(gates_1271),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0000111111110000101011010110111111111001110000100011100111111001)  
) LUT6_161 (
   .O(gates_327),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0101011110011011000110011011100111101000000111100100001011011011)  
) LUT6_162 (
   .O(gates_904),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1111001101101010010110101001100111111111111100110110111111100101)  
) LUT6_163 (
   .O(gates_1290),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b1001001101011100111010001001101010111111011000111110101101001110)  
) LUT6_164 (
   .O(gates_735),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0111101011100001001000000010101010101110110001010100000100010101)  
) LUT6_165 (
   .O(gates_722),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0101110100100010001101111100000001010010011001101011010111111111)  
) LUT6_166 (
   .O(gates_1522),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0011010100000110101010001100011110101010001110011101100000100010)  
) LUT6_167 (
   .O(gates_1118),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0100010100011001100001100011100110101000100011000000000011100000)  
) LUT6_168 (
   .O(gates_1385),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b1110010010000111100110110011001001011100011011001100000111100001)  
) LUT6_169 (
   .O(gates_1493),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1011100100110110100010001010010111001011110111101010010001110011)  
) LUT6_170 (
   .O(gates_326),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b0110100000101111100110100011011100010000000111110110101111001110)  
) LUT6_171 (
   .O(gates_1489),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0011010111010101010101010011111101101011001100011100011101111101)  
) LUT6_172 (
   .O(gates_359),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1111111001101010010101010000111001011001100000110000101111001001)  
) LUT6_173 (
   .O(gates_230),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1111110100111101111111000100011111000001111011100001111001101011)  
) LUT6_174 (
   .O(gates_13),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1000111101110101100100100011001101110001010111100111101001011111)  
) LUT6_175 (
   .O(gates_16),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1110110101111101100111010010110011010000100000011010001100000010)  
) LUT6_176 (
   .O(gates_428),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0001011000110010110101101101010101100111100011100000010100011101)  
) LUT6_177 (
   .O(gates_669),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1011101000000001100100100011010111110101001111101001011000101000)  
) LUT6_178 (
   .O(gates_595),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0010010101000111000001000000111011001111100101000000001111000000)  
) LUT6_179 (
   .O(gates_501),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1101110000100111010110101100011000001100110010110101100001101011)  
) LUT6_180 (
   .O(gates_1030),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1110111011101000101100011101111101110101100011001011010111011001)  
) LUT6_181 (
   .O(gates_474),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0000000011010110111100101111100111100111111001101000110110000001)  
) LUT6_182 (
   .O(gates_1303),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0010100000101011111000111111111011101000011101111111000100001010)  
) LUT6_183 (
   .O(gates_1028),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000000001111100001001000011110100111110000001101110100111011100)  
) LUT6_184 (
   .O(gates_1161),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0110011100010011011101100101010110111011101001001101110010111000)  
) LUT6_185 (
   .O(gates_1514),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0001010011100001010011110011110100111110110010000100100010010111)  
) LUT6_186 (
   .O(gates_195),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1010101001111101010100010111111010101110001100101011010000010100)  
) LUT6_187 (
   .O(gates_387),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0111010101111111010100101111101011111101010100100011110000001100)  
) LUT6_188 (
   .O(gates_632),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0011000000001011111011110100111000110110010100101101011100110010)  
) LUT6_189 (
   .O(gates_105),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1001100001010011011001101010000010101101011100111101101000000001)  
) LUT6_190 (
   .O(gates_50),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0011000101001111101011111100110011110110101000010000001101100011)  
) LUT6_191 (
   .O(gates_1147),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1000000111110010000101001101100101100011111011001110100001110100)  
) LUT6_192 (
   .O(gates_1527),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b1110110001100101001001101011100100101111010100000110011110110110)  
) LUT6_193 (
   .O(gates_289),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1000001011101101100100101000100000000110011011110010011101001101)  
) LUT6_194 (
   .O(gates_725),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0011101100100010011100010111001010011000100010001100111000101100)  
) LUT6_195 (
   .O(gates_1046),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0011110011111101011100000101100001000011110000100010111101101110)  
) LUT6_196 (
   .O(gates_1163),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1011001111010000010010101111111000111110111011011100111000011010)  
) LUT6_197 (
   .O(gates_1305),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b0110001111010111010011111011100111101111110011100100111111010000)  
) LUT6_198 (
   .O(gates_1433),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0011001010110100000101000010011101011100011100101010000010001110)  
) LUT6_199 (
   .O(gates_287),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0001101101010111011101011101110010111110011000000001010101001100)  
) LUT6_200 (
   .O(gates_962),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0111111000000100000001010100010101011110100000100011111000110101)  
) LUT6_201 (
   .O(gates_1370),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0011000001110001000110100010111100100011110100000100100010011100)  
) LUT6_202 (
   .O(gates_56),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1101010100011011101111100101100010011010000001000011110001000100)  
) LUT6_203 (
   .O(gates_522),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0001110100101011011100000001000010100010001010111001011010001110)  
) LUT6_204 (
   .O(gates_391),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1001000000110100000110001010100001001001001001111011000001110101)  
) LUT6_205 (
   .O(gates_668),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0110110111001011010011001101111001001000000011001110000001011110)  
) LUT6_206 (
   .O(gates_949),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1000110000111001101100110000000011100001101111011000001000111100)  
) LUT6_207 (
   .O(gates_700),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1010001100010000101111100011011111110100101000100000111000001111)  
) LUT6_208 (
   .O(gates_1072),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0100110100110000000001110110010111111000001110010110100010110111)  
) LUT6_209 (
   .O(gates_740),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0010001111000111100110100001010010101010110010110111011111010001)  
) LUT6_210 (
   .O(gates_1206),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0101010001101001000101100101111011101000011100110110010001111100)  
) LUT6_211 (
   .O(gates_1383),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0110110100011001101001010110100111100111010101011000011101011111)  
) LUT6_212 (
   .O(gates_93),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1001100100001101100111100100000011011101000010001010010111111100)  
) LUT6_213 (
   .O(gates_503),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0100001010100001001101100101000111011000001010000111010110000010)  
) LUT6_214 (
   .O(gates_1320),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1000011111011011110101001101101011001001110001010111100010101000)  
) LUT6_215 (
   .O(gates_1306),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0011010001111000100101010100100100101101010001110111101111001001)  
) LUT6_216 (
   .O(gates_177),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0001000111100110000110001011001001110110111111110100111110110000)  
) LUT6_217 (
   .O(gates_314),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0011011111011110101101010101111101010101011100111111001101101100)  
) LUT6_218 (
   .O(gates_879),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0011110101001011000100000101011000010000110110011110010001001011)  
) LUT6_219 (
   .O(gates_926),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1101100100010000001101110110111111000100110101101101101001011001)  
) LUT6_220 (
   .O(gates_19),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b1110110000000001101100111001101100111000001000000011011010101100)  
) LUT6_221 (
   .O(gates_1341),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0100001010101010110111001011011111110001001011101010111000001110)  
) LUT6_222 (
   .O(gates_997),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0111110110100000111011101100011100001001111101011101011000011010)  
) LUT6_223 (
   .O(gates_1018),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0110101110111111011111111110001100010110000111101111001111101001)  
) LUT6_224 (
   .O(gates_938),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b0001011110001010100101100110001000010101110100000001000100111100)  
) LUT6_225 (
   .O(gates_422),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1011000000010011111000101101000011011001011011111001110011100001)  
) LUT6_226 (
   .O(gates_652),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1111100100111111001101101100010011001000010111001111111100111000)  
) LUT6_227 (
   .O(gates_1116),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0000000011100001111001110110010110001101001010000100010100111111)  
) LUT6_228 (
   .O(gates_1548),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0101001001110110000111010010000011010111110101100101101010100011)  
) LUT6_229 (
   .O(gates_457),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1101010011101111011000010101001010100110001011010011000111111001)  
) LUT6_230 (
   .O(gates_987),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0001101010101110010010011111110001011000011111111011110000011000)  
) LUT6_231 (
   .O(gates_14),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1000010101001101110101101000001110010110100111000000010000001101)  
) LUT6_232 (
   .O(gates_249),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0100001010101111100010010111100010011011110010111011101000101100)  
) LUT6_233 (
   .O(gates_1549),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1110000010001100110000101101101101001100010010100010100101110100)  
) LUT6_234 (
   .O(gates_1245),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1111000000101001110111101101101000111111010100010111010101001111)  
) LUT6_235 (
   .O(gates_639),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0101100110111010101101010010111000000110110100001111001110000011)  
) LUT6_236 (
   .O(gates_186),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1111100100111100001010010001011001011111011010010000011111111010)  
) LUT6_237 (
   .O(gates_57),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1101111100110110010111100001001001010011111110001000101001111001)  
) LUT6_238 (
   .O(gates_881),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0001101011000100101100011100100111011000111001000000001001010001)  
) LUT6_239 (
   .O(gates_188),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0101001111010111101001011100010110101101111011100001100011001111)  
) LUT6_240 (
   .O(gates_1317),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0111011010001001101011010111011111010100101111001101101100110101)  
) LUT6_241 (
   .O(gates_316),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1011110001111101111100011101000100101110100001110000101100101001)  
) LUT6_242 (
   .O(gates_1380),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0101100011100100000010001001101010100001110100111010101100100100)  
) LUT6_243 (
   .O(gates_730),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0101101010111000111110001011010111111111000001100100110000100111)  
) LUT6_244 (
   .O(gates_984),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0100001010111000001001100110100000001110100100100000011111011010)  
) LUT6_245 (
   .O(gates_750),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1001011111011011111111010101010000000100011111110110001110000100)  
) LUT6_246 (
   .O(gates_349),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b1101000111001000011000011001111000111100011100010010101000001001)  
) LUT6_247 (
   .O(gates_1089),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0001110010000101000101100101011011110101100100001111110010111000)  
) LUT6_248 (
   .O(gates_1461),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1011011011100101110101000010000011001110110010011001110011101100)  
) LUT6_249 (
   .O(gates_625),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1011001011101101000111100010101101110110110001101010100011101100)  
) LUT6_250 (
   .O(gates_1135),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0111010010100000111111000010111100010101101110000000100011001001)  
) LUT6_251 (
   .O(gates_442),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1011111111100011100100101101011001110111010100101110110001100110)  
) LUT6_252 (
   .O(gates_1457),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0100011000011011001010001100110100011110101110111000011001101111)  
) LUT6_253 (
   .O(gates_792),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1000110100011101100000111000011010011011101100111011011000111101)  
) LUT6_254 (
   .O(gates_411),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0010011101100110100000110010101100111111010110010100011001010000)  
) LUT6_255 (
   .O(gates_1402),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b1001000100110010100011010100110111011010111001011111011110001101)  
) LUT6_256 (
   .O(gates_1277),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b1001100001010001111101000010011001010001011000000011110110100011)  
) LUT6_257 (
   .O(gates_693),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1100011101100001010010011100011111000010100110001110101100010001)  
) LUT6_258 (
   .O(gates_450),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0011100011110011111101000110000101010001110100011110010011110101)  
) LUT6_259 (
   .O(gates_793),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0001111100010011010100010000010111001100110101111011100000001111)  
) LUT6_260 (
   .O(gates_531),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0010000100010011111001010011011000110011011110000110110111111011)  
) LUT6_261 (
   .O(gates_1237),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0100000001011110011000100101110011111110001101011110010111011010)  
) LUT6_262 (
   .O(gates_1177),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1010010110011111101011100101110010111101101100100011001001110001)  
) LUT6_263 (
   .O(gates_470),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0100000011101001101001010000000100000011011101111001000000101100)  
) LUT6_264 (
   .O(gates_1367),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0110000011111010001011010100000101101110000011001110111101110100)  
) LUT6_265 (
   .O(gates_1270),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1101101111110100110000001001110100100110000000000110010100011100)  
) LUT6_266 (
   .O(gates_798),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1101110000001000000110100011010001000100001010000000101101001001)  
) LUT6_267 (
   .O(gates_659),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1001101100011000010110010100011001011100101110010011001011011000)  
) LUT6_268 (
   .O(gates_942),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0011000011101100110111001001101110110101010011011100100100111001)  
) LUT6_269 (
   .O(gates_118),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1101111011001111000000011100010100101000010110101101010000101011)  
) LUT6_270 (
   .O(gates_1346),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0010011010000110000110011111010011111101111000010100010111110010)  
) LUT6_271 (
   .O(gates_406),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0100011101001011000111101100100101111111011010100010100111010011)  
) LUT6_272 (
   .O(gates_1498),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1101100000010111011101100000101011110111000101111010001110011010)  
) LUT6_273 (
   .O(gates_208),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0110100001000110000001100101111001110000011011111101101110000101)  
) LUT6_274 (
   .O(gates_386),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1101100110100000100010101111001000101011010010111010011111010111)  
) LUT6_275 (
   .O(gates_665),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1001001001101100101001101100110111011110000101100010100101000101)  
) LUT6_276 (
   .O(gates_824),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1100100110010100101000001011010100111100010000111010111100101010)  
) LUT6_277 (
   .O(gates_404),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b1110111010100011001111101000100111000011110001110110000110001110)  
) LUT6_278 (
   .O(gates_200),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b1100010110000100111001110011111110000110000000110010011101010001)  
) LUT6_279 (
   .O(gates_536),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0101100100001011010101110000001100111110100100011100110011010011)  
) LUT6_280 (
   .O(gates_1145),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1111101001001110000110011000101000111010111001010101001101101000)  
) LUT6_281 (
   .O(gates_647),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0010000000010101010111010101111001111010011101001110000100011001)  
) LUT6_282 (
   .O(gates_587),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0111101000010000010001100000000110110011010010101111100011001011)  
) LUT6_283 (
   .O(gates_460),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1110010011101111100001110000010001111110111110101010001100100111)  
) LUT6_284 (
   .O(gates_357),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0110001000001011101111011001000010100001100011110101100001111101)  
) LUT6_285 (
   .O(gates_902),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1110111100100000001000001001011011101101100011010010110001100111)  
) LUT6_286 (
   .O(gates_1418),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0000011110011110101110110100010010000000011010100011101011100111)  
) LUT6_287 (
   .O(gates_1170),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1110110000000000010101010011000100010010011101001101110111011101)  
) LUT6_288 (
   .O(gates_1403),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b1101100001101100010001111001101000001110001111111011011100101110)  
) LUT6_289 (
   .O(gates_444),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1010100110011011111011110001111101100101110001011111110010111000)  
) LUT6_290 (
   .O(gates_648),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0011001110110110010010000011000111111001001011100110010101110100)  
) LUT6_291 (
   .O(gates_440),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1101100101111111000111000110111111111011111111010010101001011100)  
) LUT6_292 (
   .O(gates_710),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0001001000110111110001101111100001010011010101110000011000001110)  
) LUT6_293 (
   .O(gates_212),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1001000100100110001110001001110111101000010100001011101100100010)  
) LUT6_294 (
   .O(gates_1299),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0000111111011001110100001010011011100000111110010101010010111101)  
) LUT6_295 (
   .O(gates_719),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1111010010100010100111100001101010011011110011110111111100001110)  
) LUT6_296 (
   .O(gates_414),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0000010110011000000110010110110110110101010011111001100001001011)  
) LUT6_297 (
   .O(gates_1296),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b1010101101001001101101110011100100100101110011111010101110110011)  
) LUT6_298 (
   .O(gates_940),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1101000001110000001010001111100101001011001000100011101001110100)  
) LUT6_299 (
   .O(gates_269),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0010101000100101000001101111111101000001011001010010011110010001)  
) LUT6_300 (
   .O(gates_1474),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b0011000000110011100110100100000101110010000001010000000000111111)  
) LUT6_301 (
   .O(gates_189),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0100011110010000110010110100111000101000111111111000001101101011)  
) LUT6_302 (
   .O(gates_1495),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1011100101101101110100010011100101111001000111110001111111010001)  
) LUT6_303 (
   .O(gates_680),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1010101001101010101011000011101110101101010000000100010111011100)  
) LUT6_304 (
   .O(gates_2),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0111011011111000111001010110000000110001101011011011110000001110)  
) LUT6_305 (
   .O(gates_895),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0101111010110100010011000100110111000100101110111011001000011101)  
) LUT6_306 (
   .O(gates_1232),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0000011011101011111011100111101110011001001011111011001101010011)  
) LUT6_307 (
   .O(gates_941),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0111010111000110100000110011101010111001010100010000101000100101)  
) LUT6_308 (
   .O(gates_677),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0111011001110110110010011100000100111110110000001001001101001010)  
) LUT6_309 (
   .O(gates_1038),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0010110110101001000011001100001011110000100011010011101101100101)  
) LUT6_310 (
   .O(gates_48),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1110001011110001111000110100100111001000101101011000111010010001)  
) LUT6_311 (
   .O(gates_217),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100100010011011100001010101000010010110010000010011111010100010)  
) LUT6_312 (
   .O(gates_924),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0011010110011111111011001110111000100011010111010011111010010011)  
) LUT6_313 (
   .O(gates_512),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1111000010111010110110100110110101101000000001101110101100011110)  
) LUT6_314 (
   .O(gates_1450),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1000001000100101010100000001111001001010000010001111110010101010)  
) LUT6_315 (
   .O(gates_1534),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1011001001011000101110000111101010100110111010110110010100101000)  
) LUT6_316 (
   .O(gates_1355),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0000100101010110100101110010011101110011110100001010100011011011)  
) LUT6_317 (
   .O(gates_1045),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b1001111001001001100010110111011100111110110101001100000000010101)  
) LUT6_318 (
   .O(gates_951),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1110010101110101000000110110011110000000101011011111010111000110)  
) LUT6_319 (
   .O(gates_223),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1010101111000001000111111010101010101001100010011000011010111011)  
) LUT6_320 (
   .O(gates_137),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1110000010100010101101010011001111011011111111110010101111101010)  
) LUT6_321 (
   .O(gates_1228),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010001100110100111111100011111100000001001000111001011110111100)  
) LUT6_322 (
   .O(gates_1478),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0100110001111110001101101100011100011100001111010000011110111111)  
) LUT6_323 (
   .O(gates_1537),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0110110010101001000111111110001010001010001100111100000001110110)  
) LUT6_324 (
   .O(gates_1252),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b1101010000011100100000111010111110001111011010110000000001011010)  
) LUT6_325 (
   .O(gates_265),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1011011010011011000011110100010100001010101000111100011001000001)  
) LUT6_326 (
   .O(gates_510),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b1100101000101000101011010100001111111101111101000111011011010010)  
) LUT6_327 (
   .O(gates_58),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1110000111110000000111101011100010011110101000000111001101101100)  
) LUT6_328 (
   .O(gates_63),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1011010011011101000001001100001011101101101011100100010001110100)  
) LUT6_329 (
   .O(gates_161),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1110110100111001001111101111101011010110000000000101110100010011)  
) LUT6_330 (
   .O(gates_1231),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0101011000000111010000100000010001001111011110111111000000100101)  
) LUT6_331 (
   .O(gates_485),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0100100100101001111110111100001111000010100100000111011011101010)  
) LUT6_332 (
   .O(gates_1326),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0100000111100111010000001100110000111100111001100011010011001000)  
) LUT6_333 (
   .O(gates_1081),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1001101000101101100010100001010110111010111100110011001010111000)  
) LUT6_334 (
   .O(gates_4),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1000000100110110000010111000010100101101110001110100111101010101)  
) LUT6_335 (
   .O(gates_1547),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b1100011101110000111011000000000111010010100000000100100000110110)  
) LUT6_336 (
   .O(gates_836),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1110001001100010010110000000100110110001010001011001101011101010)  
) LUT6_337 (
   .O(gates_84),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0111101000000011000011111010011001010001010110001000101000101111)  
) LUT6_338 (
   .O(gates_462),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1111010110101010111100100101100101010011101001110100111011011000)  
) LUT6_339 (
   .O(gates_850),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1110011000111010010011011001011101110101000000101101011101000111)  
) LUT6_340 (
   .O(gates_752),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0000011001011101111010000101111111110101110111110101000110111100)  
) LUT6_341 (
   .O(gates_275),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1110010001010101110010011011100101000100000100010100100101101100)  
) LUT6_342 (
   .O(gates_622),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0100110001100010110101000110011011110011101100001001110011011001)  
) LUT6_343 (
   .O(gates_1369),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0011010101111000010111000001100111000100000011111111111110100000)  
) LUT6_344 (
   .O(gates_489),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0001010101110001010010110100000000111010110000110110010110000101)  
) LUT6_345 (
   .O(gates_548),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1101100110000100011010110100100011110110111101100001111111101011)  
) LUT6_346 (
   .O(gates_544),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1101011110011000010100110101110101111100111011011111001111111010)  
) LUT6_347 (
   .O(gates_1042),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0011000010100100000111111010111000010001010000110100010101101010)  
) LUT6_348 (
   .O(gates_906),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0100110010000001000010000011000101110101101001101000101111010101)  
) LUT6_349 (
   .O(gates_1330),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1000111001110100100011100001111110110001110001101011011110010101)  
) LUT6_350 (
   .O(gates_401),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0110001000111000111010100100111010101001010000000001011100110101)  
) LUT6_351 (
   .O(gates_1053),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0011110010011001001111101111101011001001011100011101001000111101)  
) LUT6_352 (
   .O(gates_256),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0101100101011010111101011000111100010110101000000001100000000111)  
) LUT6_353 (
   .O(gates_128),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0101001011001011000110011101111010011111001110001111101000010110)  
) LUT6_354 (
   .O(gates_1318),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1100010100111101001100111011001001101100001001100111010100101000)  
) LUT6_355 (
   .O(gates_823),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0111111010000111011110111001000101000111000110110111011100000100)  
) LUT6_356 (
   .O(gates_708),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0011101001111100000110111011111111000110010000111100010110101101)  
) LUT6_357 (
   .O(gates_866),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1110110000100101110011101111000110101001000001100111000101011001)  
) LUT6_358 (
   .O(gates_1134),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1111110011101001110011110100011111010001001101001010001000101010)  
) LUT6_359 (
   .O(gates_1444),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0011110001010001001101110010000011010101000101111010110001100011)  
) LUT6_360 (
   .O(gates_362),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0110111000101001111011101000110001111101001011010010101001001110)  
) LUT6_361 (
   .O(gates_1499),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0010110010001011011101011100011000011011110010110111111001111000)  
) LUT6_362 (
   .O(gates_449),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1110101010111110011000001001110011100000001001011101110001111001)  
) LUT6_363 (
   .O(gates_341),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0100000000011010000110000111100001111011010100101111010111111101)  
) LUT6_364 (
   .O(gates_1496),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1110101011111000101011110111100011111010011110100100000111000000)  
) LUT6_365 (
   .O(gates_103),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1011010001000010111101001011100000110000010101001111000011000000)  
) LUT6_366 (
   .O(gates_799),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0011011001010001011001110000111101011111011011010011101010010100)  
) LUT6_367 (
   .O(gates_1463),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1001100100110000011011010011101110010111100001110000001100011001)  
) LUT6_368 (
   .O(gates_616),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1000100000011000011100100101101001101110100100111110001000111110)  
) LUT6_369 (
   .O(gates_412),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1111011110101000101010111111000110001010100100001110000111011000)  
) LUT6_370 (
   .O(gates_504),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1101110010100011001110111101101100110001110001111000001011011001)  
) LUT6_371 (
   .O(gates_848),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1111101101110001110110110001011110111111001100101110000001100001)  
) LUT6_372 (
   .O(gates_9),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0000011010111110100110011011101111001101100010101010100100011011)  
) LUT6_373 (
   .O(gates_1242),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0001011001101100011010011011011100111110000111010101111010000000)  
) LUT6_374 (
   .O(gates_1176),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b1101110000001011010101001011010101100101010010101001110111010111)  
) LUT6_375 (
   .O(gates_1233),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b1001010010101101001011010001011111100110001111111111111100110111)  
) LUT6_376 (
   .O(gates_1090),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1010010010100101100000110101100100011001011110001011010110111011)  
) LUT6_377 (
   .O(gates_279),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1110111101111010001001000011011110100100100110001000010011111100)  
) LUT6_378 (
   .O(gates_1344),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0001010100100011111110000000011110111111100111101011001100010000)  
) LUT6_379 (
   .O(gates_1192),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0000010100101001101110001001110011111000010101100111100011010101)  
) LUT6_380 (
   .O(gates_959),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1101010110010000100111100010011000000111101001110001000100011001)  
) LUT6_381 (
   .O(gates_870),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0000001001001101000111001111110001010000110111000000010011100001)  
) LUT6_382 (
   .O(gates_953),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0111111101101101011000010110001101001001101101110010100100110000)  
) LUT6_383 (
   .O(gates_840),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1100010110011101110111110111010010001101111011101001010000111110)  
) LUT6_384 (
   .O(gates_736),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b1001010111010010101100000110000000110000100000111011000011100011)  
) LUT6_385 (
   .O(gates_1288),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1111011001010010101010010110011011011111100001001110110001011100)  
) LUT6_386 (
   .O(gates_1099),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0010101111111001011110011101111001101101010101011010110100101000)  
) LUT6_387 (
   .O(gates_1102),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1100001100111110100011000111001100001101001101100100010100101011)  
) LUT6_388 (
   .O(gates_1545),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1101111011010011101000100110001011101111111001000011110000110110)  
) LUT6_389 (
   .O(gates_1469),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1001000011001001111010100000110101110010100100001111100110011001)  
) LUT6_390 (
   .O(gates_376),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1000000101011011110100111010001010110000100110011001100000011000)  
) LUT6_391 (
   .O(gates_607),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0011011010000110000010111100010110101011101110000111001111000100)  
) LUT6_392 (
   .O(gates_1185),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0010011001101111010000100001001100011001111010010100010011000101)  
) LUT6_393 (
   .O(gates_333),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b1110100100100101000000010001011101010101100110001111000110001110)  
) LUT6_394 (
   .O(gates_108),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1101001111000010001001110010001001010001101000110100110100101100)  
) LUT6_395 (
   .O(gates_1504),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b1001000001111110010111100001100011000010101000101101111001100100)  
) LUT6_396 (
   .O(gates_248),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1010101111101011000100010010011001010101010101010100110010011001)  
) LUT6_397 (
   .O(gates_1165),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b1111001001111000001000001100010000011110011111011101111101110101)  
) LUT6_398 (
   .O(gates_1160),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1110010000001000000101011101011000110011011101111011011010000110)  
) LUT6_399 (
   .O(gates_96),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1100111010000110001100010111100011010000011000010101000000101110)  
) LUT6_400 (
   .O(gates_885),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0110111111010010110100100110001000001100101101111100110110011100)  
) LUT6_401 (
   .O(gates_363),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0110100001010111010110111000110011000111101101011110101011110010)  
) LUT6_402 (
   .O(gates_90),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001010000100100111011110001100111001000001010101100001101100111)  
) LUT6_403 (
   .O(gates_968),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b1011110101001011010110001011011100100110001010011110010110000101)  
) LUT6_404 (
   .O(gates_1284),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1100111011010011010001000110110110100111100100000100011100100001)  
) LUT6_405 (
   .O(gates_322),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0010010011010010010011011000010010110000011000100101011110000001)  
) LUT6_406 (
   .O(gates_1222),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b0001001011111110001000011011111100110000111101010110011001001101)  
) LUT6_407 (
   .O(gates_575),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1001000001101000110000011011100100000111011100110001111100100111)  
) LUT6_408 (
   .O(gates_1060),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0101011001000001000011000111001110111100110100011000010011110011)  
) LUT6_409 (
   .O(gates_1526),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0111001000101000110011010000110110010011001011001000000000001100)  
) LUT6_410 (
   .O(gates_934),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0100010010011010100010110101101110010010111101110010011100101000)  
) LUT6_411 (
   .O(gates_25),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1101010111000111011100111000110100111110110111111110110011001011)  
) LUT6_412 (
   .O(gates_1512),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0110001001000011111010101110011001111010110101011001100001001000)  
) LUT6_413 (
   .O(gates_835),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0111001010101111111110001010001101101110101010101011001001110100)  
) LUT6_414 (
   .O(gates_209),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0101011101000101000111100101101101100000011110101111001010000100)  
) LUT6_415 (
   .O(gates_1332),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0011001111101011110000111001000001001101100001100111110100100110)  
) LUT6_416 (
   .O(gates_766),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1101001011101100000100001001111001000100100111110111001001001100)  
) LUT6_417 (
   .O(gates_1009),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1001010011110111110111010011100110111011000111101111000000010100)  
) LUT6_418 (
   .O(gates_609),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1101100111111110110011010100011101000101000000010111001111100010)  
) LUT6_419 (
   .O(gates_291),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0111101100110100010010010101001111111001010100100101010111111011)  
) LUT6_420 (
   .O(gates_585),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b1011010000111110100100010011011101111100010010101100100000001100)  
) LUT6_421 (
   .O(gates_117),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0111001000111000100110101111010100100111111110101110011000001101)  
) LUT6_422 (
   .O(gates_1427),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0110000110010110111111101110000001100101000111011111010100000110)  
) LUT6_423 (
   .O(gates_1347),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1100100010010111101010101101010000011101111010110001011111011000)  
) LUT6_424 (
   .O(gates_334),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0101000010010111101011011101001011001000011011011111001110010001)  
) LUT6_425 (
   .O(gates_340),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1100001011011111101011001010111000001111100100000110001011111000)  
) LUT6_426 (
   .O(gates_1027),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1101011001111101011101000110110100011011111111101100110010010110)  
) LUT6_427 (
   .O(gates_173),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1110101001000011010010101111011010010100010001001101100100100110)  
) LUT6_428 (
   .O(gates_982),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1110111111111100110101001001000100011011010110101110100111000100)  
) LUT6_429 (
   .O(gates_467),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0000001001000011101000000111010101110001011101010110011101010110)  
) LUT6_430 (
   .O(gates_880),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0110010100100100010110110101000100100110011010101110010000110100)  
) LUT6_431 (
   .O(gates_1382),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0100100010001000011010000000110100011101001111000000010110000010)  
) LUT6_432 (
   .O(gates_681),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001000011110100000011100111101101001010010001111000100111000011)  
) LUT6_433 (
   .O(gates_620),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1011000110101010010011101111110110101101001111101100000001101000)  
) LUT6_434 (
   .O(gates_153),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1010111001100000000100001101001110010101001001110001110010100110)  
) LUT6_435 (
   .O(gates_570),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1111000101100000111001101110000000000110111110010110101110100011)  
) LUT6_436 (
   .O(gates_549),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0111111100111000100011101100100000010001110100011001010110010111)  
) LUT6_437 (
   .O(gates_425),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0100110010110111111100001000110111001000001000110101111001101111)  
) LUT6_438 (
   .O(gates_1482),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0011001101110000010100000011101001100111000001100101000101000111)  
) LUT6_439 (
   .O(gates_1298),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1000111001111110000010101100001100001000001111111010100010011111)  
) LUT6_440 (
   .O(gates_1084),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1001101010011001101101011011111001001000011000001110011100001011)  
) LUT6_441 (
   .O(gates_804),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0110011011000011011010101111010010011010010101011000001100000011)  
) LUT6_442 (
   .O(gates_5),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0111111101100000101100111100001000100000100000101101100011010110)  
) LUT6_443 (
   .O(gates_1532),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1100111100111111000011010011100101101101111001000100110100010110)  
) LUT6_444 (
   .O(gates_1389),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b1011101000010010010001011001101010110011010000001011100101110010)  
) LUT6_445 (
   .O(gates_916),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1100001011010101110111110000010100111000101110011011110110001010)  
) LUT6_446 (
   .O(gates_1248),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1111011101010100001011010010001100110010100110000111001001011101)  
) LUT6_447 (
   .O(gates_862),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0111011111110100111000000001011010100101111100100001100111011011)  
) LUT6_448 (
   .O(gates_936),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0010000011101000011011011111010001001110110100000011010101001101)  
) LUT6_449 (
   .O(gates_583),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0000101100001010100010001000011111010100101001001101110011011111)  
) LUT6_450 (
   .O(gates_1115),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1000011111111100011110100001100110101011101100010001101110101110)  
) LUT6_451 (
   .O(gates_1539),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0011110101010011000010110011110011010010001111110110011111011000)  
) LUT6_452 (
   .O(gates_1438),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b1010001111010110000110111010111000001001001011110000100111011011)  
) LUT6_453 (
   .O(gates_631),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1011110001010101001011100000011010001011010011101100000011111111)  
) LUT6_454 (
   .O(gates_1508),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1010000011100000111111111000101001111101010011010101000001110110)  
) LUT6_455 (
   .O(gates_1175),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1111111000110011011110010010010011010011110110010101100100100111)  
) LUT6_456 (
   .O(gates_892),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0010111001001110111101010110100010111110011000110100001011001000)  
) LUT6_457 (
   .O(gates_762),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1101111101111001011101101010110100011101010101110101111010001001)  
) LUT6_458 (
   .O(gates_805),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1001001011000101010010011101111000110000001111000101010110101101)  
) LUT6_459 (
   .O(gates_1443),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1000011010001101110100000011100110100000110100100010001110001011)  
) LUT6_460 (
   .O(gates_382),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0011010010101100110100011011111110000111001000100000011011111000)  
) LUT6_461 (
   .O(gates_1432),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1111011010100011111001100010100111110100010010001101111110110110)  
) LUT6_462 (
   .O(gates_1393),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0110111101110001000110101110110100111011010001010111000111101001)  
) LUT6_463 (
   .O(gates_78),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1010111001011001000001110100100111110101011111111010010011110011)  
) LUT6_464 (
   .O(gates_1157),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1100011000101010001100111100001110010001010101100110110101000001)  
) LUT6_465 (
   .O(gates_1188),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1010010111001000110010011101100010101011010010111111101000101000)  
) LUT6_466 (
   .O(gates_262),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0110001111000011010011100011111001011100000001001110011011011010)  
) LUT6_467 (
   .O(gates_537),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b0100011110101111101111100000010000010001111000011000110101001111)  
) LUT6_468 (
   .O(gates_507),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1100110011010100001011000001101111100000100010010100100101100001)  
) LUT6_469 (
   .O(gates_808),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0001001000001100010010000011100101111111001010101110101111011111)  
) LUT6_470 (
   .O(gates_42),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0101010011010101001011001111101010101001011111010010101100010010)  
) LUT6_471 (
   .O(gates_380),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0010001011001111000101100111111100010001101100101110100011111011)  
) LUT6_472 (
   .O(gates_491),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1011000111111000100010111111010001110100010111011110001101010110)  
) LUT6_473 (
   .O(gates_563),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0100100110110101010101101101101010111110101111101001111001110110)  
) LUT6_474 (
   .O(gates_1446),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1011010100011110010010111100001100000100111011101101011110001101)  
) LUT6_475 (
   .O(gates_239),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0000010110011001011111010010000110001010011001100000000001011111)  
) LUT6_476 (
   .O(gates_592),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1110100011000111101000000110011001111110111001100000001100000110)  
) LUT6_477 (
   .O(gates_1225),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1010101100100001100111111000010011111100001010111000000100001101)  
) LUT6_478 (
   .O(gates_224),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1010011101101100110000000011111110000010001111101101000011000111)  
) LUT6_479 (
   .O(gates_600),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1010100001110100011001000101010100011100101011001100011000000010)  
) LUT6_480 (
   .O(gates_141),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b1100111111011111011101000100001011001010111111100100111101001001)  
) LUT6_481 (
   .O(gates_308),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1011011100111110011010100100000100000001001100100111111011111011)  
) LUT6_482 (
   .O(gates_274),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b1100110000111101100111000000010100100111111001010110011101010010)  
) LUT6_483 (
   .O(gates_1465),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0010010010101100001001101100110100011000000111101000010100101111)  
) LUT6_484 (
   .O(gates_374),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0100110011011101110100001011110100101111010011101111000110110111)  
) LUT6_485 (
   .O(gates_299),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1010001100100010110110101011010011101010101101000110001010001100)  
) LUT6_486 (
   .O(gates_1541),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0111100101101111011011000000110001110000100010001000111000100101)  
) LUT6_487 (
   .O(gates_945),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1011100111101001000001110011001011011011011011111100100011111100)  
) LUT6_488 (
   .O(gates_1401),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1010101110101100100101111110010101000111100010010101111000010001)  
) LUT6_489 (
   .O(gates_847),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0100110111000110111000100100101011111110011000010111011110101101)  
) LUT6_490 (
   .O(gates_1070),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0101010100111011110000001001000001100001001000110000011000001010)  
) LUT6_491 (
   .O(gates_914),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0100011011100001110111011010000100000010111101111000111101001111)  
) LUT6_492 (
   .O(gates_1137),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1101000101111001111011011000000011011101111000010011100111110011)  
) LUT6_493 (
   .O(gates_1052),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0001110100010110010100100010111110000100011001001110010001010001)  
) LUT6_494 (
   .O(gates_858),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0101001101000001001111011111001011001010110101001100111101101011)  
) LUT6_495 (
   .O(gates_1529),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0011001110001111110001010001110111001101000101111100111000111111)  
) LUT6_496 (
   .O(gates_40),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1000011001101011110000001001110000000001111100100000100000011111)  
) LUT6_497 (
   .O(gates_293),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1101010010111111010011001100110100101001110011010101100000110100)  
) LUT6_498 (
   .O(gates_172),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0110011010001001000011001001011000000001000010011010000101010111)  
) LUT6_499 (
   .O(gates_1417),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b1110110000011100001110110111010110010001101111011001101010101101)  
) LUT6_500 (
   .O(gates_72),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1100011100010001111100111111111010111111010101111100011000000101)  
) LUT6_501 (
   .O(gates_332),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1110011100101011010011100111110011111110111111010111001000101100)  
) LUT6_502 (
   .O(gates_1220),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1110111101001111010011110011101111000111001101010110001111010111)  
) LUT6_503 (
   .O(gates_869),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100110111000011001011001100101011011101101010111111001100000111)  
) LUT6_504 (
   .O(gates_728),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1001110000000101000000101011111000101000011010001111000010100110)  
) LUT6_505 (
   .O(gates_1293),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1101100101011010001010000010111000001010000001110010001001101111)  
) LUT6_506 (
   .O(gates_932),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1011111110010110100000110100000110001100000101001111001000100111)  
) LUT6_507 (
   .O(gates_1279),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0111000010010111101100010101001110111001110111011001101010101001)  
) LUT6_508 (
   .O(gates_1219),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0110101011010101111101011101111001010111001110011100000110111000)  
) LUT6_509 (
   .O(gates_46),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0000100101000111010010000110010001011111010100000000010111110110)  
) LUT6_510 (
   .O(gates_828),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1011000110101000110001101111000101110110011000100111010011001001)  
) LUT6_511 (
   .O(gates_1536),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1101101010101001001011101101000001001001100010010110101101111011)  
) LUT6_512 (
   .O(gates_244),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1000000111011101110110100001111001101111101001001010010110001110)  
) LUT6_513 (
   .O(gates_520),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0101100010111000100111010100010010000100100010011110100011110111)  
) LUT6_514 (
   .O(gates_1077),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1100000110111111001111111110011001110000010110010111010101100001)  
) LUT6_515 (
   .O(gates_1104),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0110101001001010110111111101100110011001011111110010010110011010)  
) LUT6_516 (
   .O(gates_115),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0110101001111111111000101011001111000001010011110111011101100010)  
) LUT6_517 (
   .O(gates_1286),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1101010001000100000111011001000011111110010100000110111101100011)  
) LUT6_518 (
   .O(gates_324),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0100100100000111010010110010001000101001100010001101011101010100)  
) LUT6_519 (
   .O(gates_1343),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1100010110111100101000010001110001101000000110011011110010010001)  
) LUT6_520 (
   .O(gates_1459),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1110010001110001001110100011101111101011100011101100110010011111)  
) LUT6_521 (
   .O(gates_106),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1011101100100001101011000000100101011001111000011111111010110000)  
) LUT6_522 (
   .O(gates_703),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1101111101110001110010111010010110111110011001011011110011100011)  
) LUT6_523 (
   .O(gates_1156),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0101101111000110111111010010100010110000001001101100101101011100)  
) LUT6_524 (
   .O(gates_516),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1101101101110001110110000101101000111100100111010110000111001101)  
) LUT6_525 (
   .O(gates_102),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010000000111110110011010110010010100001011010101010111010110111)  
) LUT6_526 (
   .O(gates_323),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0101011011000101000100000000111001110101010001010100000001110000)  
) LUT6_527 (
   .O(gates_1128),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0011100000100100101100100001101011001101010000101101011110101110)  
) LUT6_528 (
   .O(gates_1458),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0110001011001000000001110111010111101000100001110110011001111001)  
) LUT6_529 (
   .O(gates_167),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1101000111011101010110111000111000110111111000100001000000001101)  
) LUT6_530 (
   .O(gates_667),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0110100101001101001000110011111001010011011000000010100000100000)  
) LUT6_531 (
   .O(gates_713),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1010110111110010111100111101001001001101111001110111010011011001)  
) LUT6_532 (
   .O(gates_1148),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b1100000110101011111010011010101100010110000011101000001011010000)  
) LUT6_533 (
   .O(gates_214),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1001101001011011001010010100111001010001111110001111010111111100)  
) LUT6_534 (
   .O(gates_1390),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0100001111100100000101101101111000111001110000000001110110000111)  
) LUT6_535 (
   .O(gates_966),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0110101000011001100000110010111001111111000000100000111010110110)  
) LUT6_536 (
   .O(gates_580),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1011110101011010111000000001100101011010011110001110011100101100)  
) LUT6_537 (
   .O(gates_871),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1010011100001011111011111100010100101110101010101111000101010110)  
) LUT6_538 (
   .O(gates_825),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1110111111100000110110111100101101010010011011101000101111110010)  
) LUT6_539 (
   .O(gates_815),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0010011100110110011110011011110101000111110100110100100000100100)  
) LUT6_540 (
   .O(gates_1353),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0101001111011001110011100101010100110111101110001001010111100010)  
) LUT6_541 (
   .O(gates_135),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1000011110111010101101111001010110100111100001110100100001110001)  
) LUT6_542 (
   .O(gates_461),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0001100010011000101001111110001000000101110011001110111001100010)  
) LUT6_543 (
   .O(gates_961),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0011101101011110001110110011100101001001101100111100010111111000)  
) LUT6_544 (
   .O(gates_886),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0001110101111000011111011100011011010000011001101110110011111110)  
) LUT6_545 (
   .O(gates_1358),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0011011111001110110010101000010001101100010111100011110010000011)  
) LUT6_546 (
   .O(gates_769),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0011111001100000111010001011101001110111010010101000100001010011)  
) LUT6_547 (
   .O(gates_1056),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b1101100111000001110111110000101000100010110110100111110001000001)  
) LUT6_548 (
   .O(gates_1183),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0101001110010001000011000101110100111100101011111111010010011111)  
) LUT6_549 (
   .O(gates_1204),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0011110110110101000010100111101100110001011011000011110100110100)  
) LUT6_550 (
   .O(gates_1502),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1000110011111000011100110100011010011100111110110111000111000111)  
) LUT6_551 (
   .O(gates_487),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1110001010100010010100100101111011011111001011111000011100000110)  
) LUT6_552 (
   .O(gates_1360),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0100110110001010011110101011011110011000000100000110101000000100)  
) LUT6_553 (
   .O(gates_1048),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0100110100010010001100100110101000000010101100101000010011110110)  
) LUT6_554 (
   .O(gates_1105),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b0010011101000001010100100010000101010101001000101111001000000000)  
) LUT6_555 (
   .O(gates_225),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1011001011110100010101011001110000111001000011100100101111000001)  
) LUT6_556 (
   .O(gates_1139),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1000111010000011000010010010011001001101101110011100111000111010)  
) LUT6_557 (
   .O(gates_185),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0111010101001001100100110100011000001001010010000001010000010110)  
) LUT6_558 (
   .O(gates_1239),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1001101110010100000010010100100100110011110110101100110110011110)  
) LUT6_559 (
   .O(gates_1282),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0011011111111011000010011011000010101000110011000100011000101001)  
) LUT6_560 (
   .O(gates_889),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1111011000011011110110000110111110101001110110111010100000100101)  
) LUT6_561 (
   .O(gates_715),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0110101110101001001011001100000110000100100010100011010011111111)  
) LUT6_562 (
   .O(gates_1230),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0010100011000010000111101010001000100111001001101001001001100000)  
) LUT6_563 (
   .O(gates_1340),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1010011010010000100010001100110001110101011011011001000101101111)  
) LUT6_564 (
   .O(gates_1240),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1011011110001111011110000001001111011000011100100010001001000110)  
) LUT6_565 (
   .O(gates_561),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0011001011111000111011111000101101101110011111101001010001011011)  
) LUT6_566 (
   .O(gates_851),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0100000101101110000010100110000001101001101011100010010010010010)  
) LUT6_567 (
   .O(gates_238),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0110111100001001001011101001101000101011000011111010010000001001)  
) LUT6_568 (
   .O(gates_1445),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0010111010100001111011000001010110011001010110011010011110001000)  
) LUT6_569 (
   .O(gates_87),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0100001001101010100010010110100000100000001101010101110000001000)  
) LUT6_570 (
   .O(gates_152),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0001011101011100001101000010100011101111110001000101011110010111)  
) LUT6_571 (
   .O(gates_1313),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1100000000000100101010111000101001011101111000010001011010111110)  
) LUT6_572 (
   .O(gates_416),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0010000011001001001010101100101100001111100001011010011111111011)  
) LUT6_573 (
   .O(gates_443),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0110001001010001010100010111100010011001010000100111010010000100)  
) LUT6_574 (
   .O(gates_159),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0011011110001111110110100100100000001000111001100100011010100010)  
) LUT6_575 (
   .O(gates_618),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0111000100000000011011010010111011101011001001001110101001110111)  
) LUT6_576 (
   .O(gates_62),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000111001111011010010101100101010010000010010001010100010000111)  
) LUT6_577 (
   .O(gates_782),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0010011111101110010111000011000101010000000010011100010000011001)  
) LUT6_578 (
   .O(gates_329),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0110100100101100001111001101010111000010101101000010111101000111)  
) LUT6_579 (
   .O(gates_1292),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0101000110100111110101001101100010001010111111001000101011100101)  
) LUT6_580 (
   .O(gates_70),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0100001100100111110101010011011111100110110010001110111010101011)  
) LUT6_581 (
   .O(gates_643),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1111110111010101001011000111111000011100011100111000000110001101)  
) LUT6_582 (
   .O(gates_1325),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1011010001110000101010111010010011001101101100001011101110110010)  
) LUT6_583 (
   .O(gates_1180),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000001011101101010011000011101011011001101101010010101010001100)  
) LUT6_584 (
   .O(gates_498),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0110010101110111011010110000110100001000010111010111001010001010)  
) LUT6_585 (
   .O(gates_145),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0110101010110011000001000111011001011101011101101111111111101010)  
) LUT6_586 (
   .O(gates_60),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0010111010110011111010010001000100101001001111001010100101011001)  
) LUT6_587 (
   .O(gates_1324),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b1101110010110011100011101110110001101110000000101011011101101111)  
) LUT6_588 (
   .O(gates_613),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1111011110011011101001110011001110010010111010111011011100000011)  
) LUT6_589 (
   .O(gates_85),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0110000101100101100111110010100100010111111101000110110101111011)  
) LUT6_590 (
   .O(gates_1399),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0001011000100100100101000000100001101101011011110001101111000110)  
) LUT6_591 (
   .O(gates_488),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1001011001100001100111011111111100001001110000000111011010010110)  
) LUT6_592 (
   .O(gates_420),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1110101111111110001011111100101011111001111010101101011111011100)  
) LUT6_593 (
   .O(gates_203),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1101011001001100100110010010011111100011100110001100011010010011)  
) LUT6_594 (
   .O(gates_1364),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0001011001010000111010101100110000001110010100100010001101110001)  
) LUT6_595 (
   .O(gates_281),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b1100000110110111010010011110010010101000111101101101000011011101)  
) LUT6_596 (
   .O(gates_1119),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0001101100100110011101110010000011001011111101010011111101010010)  
) LUT6_597 (
   .O(gates_666),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0110011001011010101010010010110100010010001111001111101001100111)  
) LUT6_598 (
   .O(gates_1186),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1111100101000010011110011100001100111000000100100111100000000101)  
) LUT6_599 (
   .O(gates_181),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0101110000110111100101000001100010111100100010010010000110110110)  
) LUT6_600 (
   .O(gates_952),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1100111001101000101101110000110001001010111010011000000001100100)  
) LUT6_601 (
   .O(gates_112),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1000011000001010111111101000011001010101100111011011001001110010)  
) LUT6_602 (
   .O(gates_655),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1011010001101101100111111000001011111000111110001001100100010111)  
) LUT6_603 (
   .O(gates_1255),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1110110100100011100101111000100001111111111100110111111000110001)  
) LUT6_604 (
   .O(gates_121),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b1011000110010110001011000100110110010110010011000100001100110101)  
) LUT6_605 (
   .O(gates_1328),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0110011010110111010111111010111011010110101111111001001100010101)  
) LUT6_606 (
   .O(gates_896),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1010110001010101100001001001110101011011100011110000100011101101)  
) LUT6_607 (
   .O(gates_441),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1010100001011011000000001100000001001011110001110111010111111100)  
) LUT6_608 (
   .O(gates_1002),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b0111100111111001110110001000011010010001110011110001100011110010)  
) LUT6_609 (
   .O(gates_471),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0011110011001001010100110111010111001110101111100010101101100010)  
) LUT6_610 (
   .O(gates_670),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1010110110001111110011000101100111001100111111011000100100001111)  
) LUT6_611 (
   .O(gates_690),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0001101001000101011110100001001010001010000010000110000100111000)  
) LUT6_612 (
   .O(gates_519),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0110001001000110100001001100101110100111011000100110010000000000)  
) LUT6_613 (
   .O(gates_957),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0000000110100111001000010010101000101101100001101110100000110101)  
) LUT6_614 (
   .O(gates_1342),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0000101110011001111000001110011111101111001001111001010000010100)  
) LUT6_615 (
   .O(gates_572),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0000111101010101001110010111110110000110010001100001000000011111)  
) LUT6_616 (
   .O(gates_1087),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1010011000110011111100000100011101001011110101101010100001010101)  
) LUT6_617 (
   .O(gates_905),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0011010111001001111100010000001000110101001011110101010001001001)  
) LUT6_618 (
   .O(gates_675),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1100100100011110001011100001010000111011011110111111000101011110)  
) LUT6_619 (
   .O(gates_304),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1011111100010100000110000001011101000110011101011000000111100110)  
) LUT6_620 (
   .O(gates_640),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0001000000000100110001001000101100101010100010111001001110000011)  
) LUT6_621 (
   .O(gates_415),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1100000111100111001010000100000110000010111101100001100110001110)  
) LUT6_622 (
   .O(gates_514),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0111011100110111101000111000001010001010001100011110111000101111)  
) LUT6_623 (
   .O(gates_254),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0100000011111010000110000110000011100100001110000101011100001001)  
) LUT6_624 (
   .O(gates_973),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0110010001110100100101100100010010110010101101101111000101100110)  
) LUT6_625 (
   .O(gates_723),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1100011100101100110101100100001001111100101100111011101011100011)  
) LUT6_626 (
   .O(gates_901),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1111111010011111110000110011111111110011110110001001001100111111)  
) LUT6_627 (
   .O(gates_1026),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0111101111110001100101111111110100011001111010111000110010111110)  
) LUT6_628 (
   .O(gates_1063),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0001000101010110010011111000011010011010011011001000100111001000)  
) LUT6_629 (
   .O(gates_1083),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1111101010001100110111011010100110111100111110000000011011001111)  
) LUT6_630 (
   .O(gates_421),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0010100111110011011110110111100111000001000100011111001000001010)  
) LUT6_631 (
   .O(gates_231),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1110000001101110110010011000001000110010100000000101000001001111)  
) LUT6_632 (
   .O(gates_1201),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1010000010011101111111101101000101111100010111110111110010101111)  
) LUT6_633 (
   .O(gates_1315),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0101010100110111010010110101000000101000001111111110011110000000)  
) LUT6_634 (
   .O(gates_228),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1111101110001010110110010110010111001011000001111111100000110110)  
) LUT6_635 (
   .O(gates_1551),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0001011101000110100111010010100001010110010000000010111010000110)  
) LUT6_636 (
   .O(gates_893),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b1111110101011010011101111001111100101110000000010100000100010101)  
) LUT6_637 (
   .O(gates_343),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0010111001000011010000110000011100100010111101011100000001100000)  
) LUT6_638 (
   .O(gates_464),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1111110011100000100000010101110111100111100000001000101000101001)  
) LUT6_639 (
   .O(gates_610),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0000000000000001010001011110010111100001001000100100100111000110)  
) LUT6_640 (
   .O(gates_477),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0110111011001110001101011110110001001001101011011110100011111110)  
) LUT6_641 (
   .O(gates_41),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1101010100111101001111110100011111001010111011110111001011001000)  
) LUT6_642 (
   .O(gates_1297),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1111101110010111100010000101000111010110100001100101011001000101)  
) LUT6_643 (
   .O(gates_1550),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0101101001100101010010101001110101011110011000001110111010001111)  
) LUT6_644 (
   .O(gates_345),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0000011000100110111010011001111000010110100001101101010101011010)  
) LUT6_645 (
   .O(gates_624),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1000010111000001001001010010100011110000001110111010001000001000)  
) LUT6_646 (
   .O(gates_1490),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0011001111111110100000001001011011010110110010011110010001101011)  
) LUT6_647 (
   .O(gates_1466),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0100100101001110100011000101110000111110101110100101001101110001)  
) LUT6_648 (
   .O(gates_578),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b1110001111001000011110001101000010110011010001010110001110010010)  
) LUT6_649 (
   .O(gates_683),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0000001011101110011011010101101111000011011101000101111100110011)  
) LUT6_650 (
   .O(gates_738),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1011101010101011011011011100101001100110001110011000110011000110)  
) LUT6_651 (
   .O(gates_1381),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0100000101110011011100100000101110100011111111001101011110000100)  
) LUT6_652 (
   .O(gates_8),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1110100001001011101100101001100011010110101110100110001011110110)  
) LUT6_653 (
   .O(gates_686),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0111101100010000011101001000000111101111010001111101000110111111)  
) LUT6_654 (
   .O(gates_852),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0000111111101010111001101010000111111011001000111111101100011111)  
) LUT6_655 (
   .O(gates_944),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1100100010100000001001001110100110111110001000000100010011010001)  
) LUT6_656 (
   .O(gates_676),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0101011100110101010111011110110100010111100011100110001001001110)  
) LUT6_657 (
   .O(gates_1125),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1001010010011001100000101110000010001000100101011110000100011001)  
) LUT6_658 (
   .O(gates_95),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0110101000010000100011110100010110001010101110100001000101001010)  
) LUT6_659 (
   .O(gates_990),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1111010110010110110011011001101000111100111111000101010101001010)  
) LUT6_660 (
   .O(gates_542),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1001111010110111010110001100010011111000101110110110001111011110)  
) LUT6_661 (
   .O(gates_729),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0101011010100001001101010101011011111001110110101110000100011111)  
) LUT6_662 (
   .O(gates_176),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0010001011111010011100110001100011101100111001011101011111010101)  
) LUT6_663 (
   .O(gates_890),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0010111000111011110101010100000100011010011000000111110011110101)  
) LUT6_664 (
   .O(gates_1485),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1100111011100101001111001010111000000101111101101010000001110111)  
) LUT6_665 (
   .O(gates_935),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0110010111010011100111111001011011001011010010110011110110111010)  
) LUT6_666 (
   .O(gates_277),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1100001001111001010100101101010001101011001101110001111010111100)  
) LUT6_667 (
   .O(gates_7),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0010001101100100010111100110100111111101010001011011010001100010)  
) LUT6_668 (
   .O(gates_1517),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1100011100100001110010110001001100010101111110110000010110110111)  
) LUT6_669 (
   .O(gates_844),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0011101010100110001100110011110111010000100010111101111011101100)  
) LUT6_670 (
   .O(gates_1376),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1101111101110111110111101000110100110111001011011101100000001001)  
) LUT6_671 (
   .O(gates_1391),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0010001010011010000100011000011110110110100110100010111000011010)  
) LUT6_672 (
   .O(gates_196),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0010000111000110000111001100011010011100001011001110111010000101)  
) LUT6_673 (
   .O(gates_426),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0011101110010010011101111000100001111011101111010000010010110000)  
) LUT6_674 (
   .O(gates_1223),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0100011101011011011010101001111000000100010111101100101000100000)  
) LUT6_675 (
   .O(gates_1500),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0011100001000011000100110011001011101010000001100010111101011010)  
) LUT6_676 (
   .O(gates_1138),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1011000110010011010100000000011001101000011010001100110111111101)  
) LUT6_677 (
   .O(gates_335),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1100101110101001101010010011110101110001110000110001101111010010)  
) LUT6_678 (
   .O(gates_1464),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1001010011110111111000010001110011101110110100000100110010111100)  
) LUT6_679 (
   .O(gates_1349),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0111110010010001110000001101111101010010111001010111010010100001)  
) LUT6_680 (
   .O(gates_726),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1001000110111010010110101101110100001010100011011001100101001010)  
) LUT6_681 (
   .O(gates_479),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b1011110011000110001011010101111101010110001001010001010110011010)  
) LUT6_682 (
   .O(gates_350),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0010101111011000111010101000100110100101101101010000010100001000)  
) LUT6_683 (
   .O(gates_493),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0100011010010011101110011101110011101001010111000100100001000001)  
) LUT6_684 (
   .O(gates_831),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b0111100000010011011010101011011110111010111011010010111101110110)  
) LUT6_685 (
   .O(gates_37),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0110000010111001101010001111100011000100010000100011000101001111)  
) LUT6_686 (
   .O(gates_405),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0101011101001111010100011010101111111000011100110011010100110110)  
) LUT6_687 (
   .O(gates_1420),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1000011001111110100110000000110011100111111001010001000010011001)  
) LUT6_688 (
   .O(gates_306),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1110100001011101010100010011000011110111101100101111111101001100)  
) LUT6_689 (
   .O(gates_99),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1011010011110010011011100100110100101110110111100000011000001010)  
) LUT6_690 (
   .O(gates_567),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0110100011001001001111110111000111001011011001101111100010001001)  
) LUT6_691 (
   .O(gates_518),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b1110110100111110111111111000101010000000111100010101001110000011)  
) LUT6_692 (
   .O(gates_1338),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1010100111010010001010011010011100110111101000001110110010101011)  
) LUT6_693 (
   .O(gates_651),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1101011000000101011100011000011010000100100100111010110101011001)  
) LUT6_694 (
   .O(gates_744),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1011101101011011111100101111010110100110110000001111100100000011)  
) LUT6_695 (
   .O(gates_490),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1010100101100000101100100001101100001001101100100000100111000000)  
) LUT6_696 (
   .O(gates_143),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1000001110110111100110110110001101101001010000000110110110001011)  
) LUT6_697 (
   .O(gates_437),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0010111011111011101100100000101000000010111001110001000100101010)  
) LUT6_698 (
   .O(gates_975),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1010010001011110110001110110010010000101000001101000010100011011)  
) LUT6_699 (
   .O(gates_1421),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0010100000100101001111111111010000111000101100110110111000001011)  
) LUT6_700 (
   .O(gates_1308),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0111101110111110011100000100111011010001101110011011101100001011)  
) LUT6_701 (
   .O(gates_1316),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b1100100101001111001001101100000000010100010000110011100010011010)  
) LUT6_702 (
   .O(gates_579),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0010101000111010111100000110100011110101110110001000000000101110)  
) LUT6_703 (
   .O(gates_727),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1110011101101100110011011001000010011111111110110010011110000011)  
) LUT6_704 (
   .O(gates_1405),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1100100111001110111000001110000011110110011011110100110000001011)  
) LUT6_705 (
   .O(gates_290),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010000010110001111100101111111000001100100110100101011100110011)  
) LUT6_706 (
   .O(gates_977),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1001011011000100110101100111011000110110101100011011010000011100)  
) LUT6_707 (
   .O(gates_303),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1110101101101000000010011100101000000111011111101011101101101011)  
) LUT6_708 (
   .O(gates_867),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0110101000110110010101101000010111000000101100011001100111100000)  
) LUT6_709 (
   .O(gates_1172),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0110100011000100110000000001101010011001101101001110000010100010)  
) LUT6_710 (
   .O(gates_356),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0100011100010010101110000010111111100101010110000110010001001101)  
) LUT6_711 (
   .O(gates_553),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0101000010000100110011111101101001010011000111000011010101000001)  
) LUT6_712 (
   .O(gates_480),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0110110001100100100000001011011001011001000110100101001111011011)  
) LUT6_713 (
   .O(gates_192),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0001110100000100001000001000000111001010010011100110110110001011)  
) LUT6_714 (
   .O(gates_1033),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0011001100110001100101101111011101011010111110111100100110011111)  
) LUT6_715 (
   .O(gates_861),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1010101010110010111011111100010010100100000101100010111100100100)  
) LUT6_716 (
   .O(gates_1032),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000000000011000000001010111110011111110000100010000010111010101)  
) LUT6_717 (
   .O(gates_59),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0010101110011011110010010000101001010101111100010000010000101001)  
) LUT6_718 (
   .O(gates_1295),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1011000111010100101000101110110100111011001011001100110000100000)  
) LUT6_719 (
   .O(gates_247),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b1011100100000010110001111010000010000110101110010100100101110101)  
) LUT6_720 (
   .O(gates_569),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0111011001011111111011010101111011101010011010001100111100000110)  
) LUT6_721 (
   .O(gates_385),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0001111101111001011001111110001010000010001100011011100111001011)  
) LUT6_722 (
   .O(gates_1213),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0101000110101000011011000101000110001011010001011100001010111110)  
) LUT6_723 (
   .O(gates_1136),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1100000000011101111110111111000010110100000000010111100111010011)  
) LUT6_724 (
   .O(gates_761),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0100111111001111010001111111011111101000001100001011101010011000)  
) LUT6_725 (
   .O(gates_1285),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0100010101111110011001000111011100100101100111110000000000000110)  
) LUT6_726 (
   .O(gates_826),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0000000101111101100001101001110001110000000001110111111011111110)  
) LUT6_727 (
   .O(gates_922),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1110010101111011110010111101001001001101111101100001111100111101)  
) LUT6_728 (
   .O(gates_505),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0111010001000011011010011110110110111100111010111000101010011011)  
) LUT6_729 (
   .O(gates_842),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0000000001010011000000110011111000110000100000010111011010000011)  
) LUT6_730 (
   .O(gates_781),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1100011000001001110100000011001100101001011010001010100001011000)  
) LUT6_731 (
   .O(gates_251),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1011111101001111000010010111011100000101110000001100101110101111)  
) LUT6_732 (
   .O(gates_320),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b1111000110110011001100011101011001000100011101011100101110100000)  
) LUT6_733 (
   .O(gates_283),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0000010000100111000010111001111100011101011110111101000110000001)  
) LUT6_734 (
   .O(gates_1178),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0011011010000000011100011111011011101100011100101010011001001000)  
) LUT6_735 (
   .O(gates_978),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0111000111110111111110111111011110111100110000010110001111001011)  
) LUT6_736 (
   .O(gates_34),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b1011010101101000001111010100110010110101000010011011101101010100)  
) LUT6_737 (
   .O(gates_1212),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0100010011011000110001111111000110110000010001101101111111001010)  
) LUT6_738 (
   .O(gates_1091),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0000101100000001101001001011000110000011000011111011000110101100)  
) LUT6_739 (
   .O(gates_699),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0010011011101101011011010110001011111110100101010011001110111011)  
) LUT6_740 (
   .O(gates_229),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0010010011100011000100000111101011101110000111110101100010000100)  
) LUT6_741 (
   .O(gates_384),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1001111110110011100101010010100010100001000001101100101010110101)  
) LUT6_742 (
   .O(gates_541),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0101001101110101111010001011010000000100001000100010010110001010)  
) LUT6_743 (
   .O(gates_378),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1001110110011111011000000101010011010110011001000111011101010101)  
) LUT6_744 (
   .O(gates_377),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0010010100010110001110000011100111011101000111101001001011001101)  
) LUT6_745 (
   .O(gates_252),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0000011010111101111110001110101111100101010100000110110100001110)  
) LUT6_746 (
   .O(gates_1468),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b0110100110100011100001100110001010000011001100010100010011011001)  
) LUT6_747 (
   .O(gates_1034),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1011010101011000011111101011101001011110000110100001101110011000)  
) LUT6_748 (
   .O(gates_833),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0010100101101010011001000001011100100101101000111001111000011010)  
) LUT6_749 (
   .O(gates_1074),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0000110011110001101011111011010101011011111101001111101101111111)  
) LUT6_750 (
   .O(gates_1361),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0001000000011100010101110011110000110111001010101111101000001110)  
) LUT6_751 (
   .O(gates_64),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1000110011010100110000100000010100100010101010000100101101110001)  
) LUT6_752 (
   .O(gates_1203),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0110001010010011110100101001001110001010000100001110101011000111)  
) LUT6_753 (
   .O(gates_768),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1011010001011010001010010000001011011111010001101010011001001110)  
) LUT6_754 (
   .O(gates_28),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1110001000110110011101100100000110111010010101000001100000001011)  
) LUT6_755 (
   .O(gates_560),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1011010111110000001100110110100101110010000001111100101001010011)  
) LUT6_756 (
   .O(gates_1182),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1110110011111110001000001110011011110011010100111100110011101001)  
) LUT6_757 (
   .O(gates_342),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0000010111010001010001001110011000001000100111001101010101101001)  
) LUT6_758 (
   .O(gates_1211),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0001010001111010100011001111100110011010111101000110101101001111)  
) LUT6_759 (
   .O(gates_937),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b1100101011101110100011001110111111001001110100010110000100001100)  
) LUT6_760 (
   .O(gates_1054),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1000100100110100111010010110101101001000110001100110111100110011)  
) LUT6_761 (
   .O(gates_35),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1111000100100001101101011000011101001100110000100110000101000010)  
) LUT6_762 (
   .O(gates_838),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1000000000100001101010011111111111101110010111011010001010111100)  
) LUT6_763 (
   .O(gates_1435),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1000011011101001100000001000100010110011110110100100000010010101)  
) LUT6_764 (
   .O(gates_608),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0110011000110000101101011110100010011000110101011100011101010011)  
) LUT6_765 (
   .O(gates_468),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0001000111101101111110011101011101000011111101111101101111110111)  
) LUT6_766 (
   .O(gates_1477),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1011100110001011111011100111010110010110110100111100011101110111)  
) LUT6_767 (
   .O(gates_111),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0001111001100011001111011010011100010101110011011011010001111111)  
) LUT6_768 (
   .O(gates_1473),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0100000111100011010000110010010010001110100011001000100110011101)  
) LUT6_769 (
   .O(gates_1120),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0100011111110110001011011100100001111111110100000001111111001111)  
) LUT6_770 (
   .O(gates_1130),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0000111011011011100011100101111110000100010011111110010110110110)  
) LUT6_771 (
   .O(gates_1394),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0110100101000110000111000000011110010010001010101000011110000011)  
) LUT6_772 (
   .O(gates_1200),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0100001011001011001001110011100001111111101101000010101010101101)  
) LUT6_773 (
   .O(gates_1029),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b0101010001111000000101100100000101011100101101100000001111000101)  
) LUT6_774 (
   .O(gates_1467),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1111100111110001110011110100001100110111111111101001010000111100)  
) LUT6_775 (
   .O(gates_127),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1000100011011011000001011010011100110101001111110001011101010011)  
) LUT6_776 (
   .O(gates_144),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0011101001100111010011100100010110101010110011100010101011001000)  
) LUT6_777 (
   .O(gates_494),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0101111010010001100011100111000111011001010011010111000011001111)  
) LUT6_778 (
   .O(gates_767),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0011111001001101110000100101000111000001001110010100111111001001)  
) LUT6_779 (
   .O(gates_1065),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0110001010110110100101111010111101110101001111011001000010110011)  
) LUT6_780 (
   .O(gates_171),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1001001011100111110111111100111100010100001010000000110011100100)  
) LUT6_781 (
   .O(gates_565),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b1011100111011111100101100111001101110111110010100111000001111011)  
) LUT6_782 (
   .O(gates_17),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0111010100100111001100110100110110011101110101110010000001011001)  
) LUT6_783 (
   .O(gates_392),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0100001110000011001000011010001011101111101010001010010111100010)  
) LUT6_784 (
   .O(gates_165),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1100100101111010110111001001110101101111100000111000000101101000)  
) LUT6_785 (
   .O(gates_1181),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1011111000110110101000001111110100000100110011010111101110001001)  
) LUT6_786 (
   .O(gates_701),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001100000100110100100010000010001100001000110011101101101110000)  
) LUT6_787 (
   .O(gates_198),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0010100011010101000000110100001111111101110101101101110101100000)  
) LUT6_788 (
   .O(gates_550),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0011001011010100110110100111101010010011010010110010010011111100)  
) LUT6_789 (
   .O(gates_156),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1010111001111100011110110101010010011000010100011100101101010010)  
) LUT6_790 (
   .O(gates_841),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b0101110001011100010011111101101011110001110101110000010111110010)  
) LUT6_791 (
   .O(gates_1440),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0101100011111010011010111101001101100101100110101000011010110011)  
) LUT6_792 (
   .O(gates_748),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1010110011000110110110011101011100101011011110110101100001100100)  
) LUT6_793 (
   .O(gates_1226),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0011001110001100100011001111001011101101111010010111101010000110)  
) LUT6_794 (
   .O(gates_126),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0101101010010110000001101010110001111100110010010010001110111111)  
) LUT6_795 (
   .O(gates_1005),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1111100110010101010010000001001100001011101010010101101110000001)  
) LUT6_796 (
   .O(gates_1449),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0000110101101100010001001000011101101000000111111110101010010000)  
) LUT6_797 (
   .O(gates_864),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0000010110010011010001101000100011111011100001000110111011110101)  
) LUT6_798 (
   .O(gates_1101),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1001110011010111010000110010101000110101101101010101101000000101)  
) LUT6_799 (
   .O(gates_1535),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0011011000110100101000110000000000110011101010110101110001110001)  
) LUT6_800 (
   .O(gates_1314),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1101010111101111011010111100110011101100001000100101110010100101)  
) LUT6_801 (
   .O(gates_43),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1001101101011001111111101101010100001101110110110000110000110100)  
) LUT6_802 (
   .O(gates_1198),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0010101001111001000001011101101100111010111101110011011100010000)  
) LUT6_803 (
   .O(gates_1414),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0001111000101111010001001010010001010101011000011001001010110001)  
) LUT6_804 (
   .O(gates_369),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0011011000111010011011011110101111001111100011010111110100001101)  
) LUT6_805 (
   .O(gates_1121),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1001000000010111010110011011110100010011010000101010100011110010)  
) LUT6_806 (
   .O(gates_433),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0101000110010011011001001010101011011111111011011110111110111101)  
) LUT6_807 (
   .O(gates_109),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0111001110001100000101010111101010011110010110111111010111001001)  
) LUT6_808 (
   .O(gates_336),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1000111000110011100001100101101000011101110111010101001000011011)  
) LUT6_809 (
   .O(gates_1523),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0111001111111110101111000100110001001110110110110110000000100101)  
) LUT6_810 (
   .O(gates_446),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1000100001101100111101101101000110000001111101100111100100001101)  
) LUT6_811 (
   .O(gates_796),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0000010000001101100101111111011110110111111101110001110010100101)  
) LUT6_812 (
   .O(gates_697),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0000100111110101100011100111111001101101100100000011111000111111)  
) LUT6_813 (
   .O(gates_795),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0010110111100001011000011100010110010010110011010101011001110000)  
) LUT6_814 (
   .O(gates_691),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0111110000111001001000001101101001001001000011001010111100101111)  
) LUT6_815 (
   .O(gates_178),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0111110100000010110001101100000011100000110110111001100010110000)  
) LUT6_816 (
   .O(gates_994),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1010111111111011101101010000110000010111111111000011000100000001)  
) LUT6_817 (
   .O(gates_1039),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1100100100010000000011110110101110100001111110001111111001000101)  
) LUT6_818 (
   .O(gates_801),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1010100111101000011110000100101000001001001001101011111111100011)  
) LUT6_819 (
   .O(gates_355),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1111101000111110111110111000101111001001000101111110110000000010)  
) LUT6_820 (
   .O(gates_626),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0000110011100111100001000100110011100011000010110110000010001011)  
) LUT6_821 (
   .O(gates_513),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0100010010010001011000010100101000000101100111100110011001111111)  
) LUT6_822 (
   .O(gates_163),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b1100011101101100100010011011110111100000110111011011100101000101)  
) LUT6_823 (
   .O(gates_930),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1001010100101000110001001110010001011101010010100011000111011101)  
) LUT6_824 (
   .O(gates_331),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0010011010010011011001000011111101010010110101110110010000001011)  
) LUT6_825 (
   .O(gates_1448),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b0111001010001011000010111010010100110011100011101100111101011100)  
) LUT6_826 (
   .O(gates_6),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0111011111111100110100111100001101011001001000000011101110001111)  
) LUT6_827 (
   .O(gates_142),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0110000101111001001001001000100000011111111101111100100001011111)  
) LUT6_828 (
   .O(gates_94),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b1010001001001100011111111110000010111111100111001101110001000111)  
) LUT6_829 (
   .O(gates_430),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0010110101111000101111001011110001111000000010011101110110010001)  
) LUT6_830 (
   .O(gates_1010),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0011101111101001101100101001111111111101001000111010110110011011)  
) LUT6_831 (
   .O(gates_1335),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b1001000110100101000010010001011010100001110000001001011000100011)  
) LUT6_832 (
   .O(gates_1424),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b1010101001111110101001001011010001101000111000101101101000100000)  
) LUT6_833 (
   .O(gates_394),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0110011000000101011110000010100011111110101000010011011000111111)  
) LUT6_834 (
   .O(gates_206),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0011011011101001001111001111101001101011111101111000001011100011)  
) LUT6_835 (
   .O(gates_497),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0100010010000010111100001001111011110001110111001010010011001111)  
) LUT6_836 (
   .O(gates_985),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b1011010011000100011000000010011110001100011001101010111000010011)  
) LUT6_837 (
   .O(gates_1122),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1100001011110110011010111101000110110110011100001001010010000110)  
) LUT6_838 (
   .O(gates_1516),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0100100101110001011100100001001010011011000000011110110111001000)  
) LUT6_839 (
   .O(gates_694),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0101010101011010110100110100010111010100101001111010010010111110)  
) LUT6_840 (
   .O(gates_746),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0110101001011110010110101100011000000101010110011111001101100101)  
) LUT6_841 (
   .O(gates_1017),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1010100011010011011100111111110011000010101000011110011010111000)  
) LUT6_842 (
   .O(gates_1193),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b0000111101010011000100000011011001111001011110111011011000011001)  
) LUT6_843 (
   .O(gates_257),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0010011110000001100010011110010000100100111101100111100001001111)  
) LUT6_844 (
   .O(gates_972),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0000111000110001101111111110011111111111001011111001111101000111)  
) LUT6_845 (
   .O(gates_469),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b0010010100000111111100110000001000000000111100010111100100110100)  
) LUT6_846 (
   .O(gates_1241),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0110000100100101010001111101011110001011100000010010111000110110)  
) LUT6_847 (
   .O(gates_1506),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1000101011010101100011100000001000011111010011100100100110010011)  
) LUT6_848 (
   .O(gates_822),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0111001010110010101000000010011101000010111010011110011010111000)  
) LUT6_849 (
   .O(gates_948),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1111111000101000000011110111010100000010100110101110001111010010)  
) LUT6_850 (
   .O(gates_182),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0010101101011010011000101000101011101110111001110000011100111100)  
) LUT6_851 (
   .O(gates_908),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b0000001011010011110101100110001101110000100010111100110100110001)  
) LUT6_852 (
   .O(gates_15),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0010110111001001111000010000000000111111010111000010000000100001)  
) LUT6_853 (
   .O(gates_114),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b1001110000011001011010110111000110100100000110001100010100101111)  
) LUT6_854 (
   .O(gates_1106),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0011011110001010110100111011001010111011101110000110110100111001)  
) LUT6_855 (
   .O(gates_448),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0001101110101110011011001010100001010010011000011111110011100110)  
) LUT6_856 (
   .O(gates_857),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1010101001110010110011011100011000011010111111100010111001001000)  
) LUT6_857 (
   .O(gates_1430),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0001100111100000111010100101011011001110111000110110010110110111)  
) LUT6_858 (
   .O(gates_465),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0001101000010101000011001111011010111011100100000010000110011100)  
) LUT6_859 (
   .O(gates_1481),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1100010001010000110101110100001011110110110010010000111101010000)  
) LUT6_860 (
   .O(gates_264),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1010101001001110001101111000001011110100100111110010101001000111)  
) LUT6_861 (
   .O(gates_241),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1010110110010110111101101000011110011010001011001111010110010101)  
) LUT6_862 (
   .O(gates_344),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b0101110110111010001011111000010001101111000000110011110011011010)  
) LUT6_863 (
   .O(gates_98),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0101010110110000001011011011001000011000011000001001000101100000)  
) LUT6_864 (
   .O(gates_1455),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000000101010011001101000110101001101110110111101010111010011000)  
) LUT6_865 (
   .O(gates_1528),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b0000100000110111010100100110101010011100111011101100010011000000)  
) LUT6_866 (
   .O(gates_24),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b1100101011111011010001000011101001100101000000101100000001000001)  
) LUT6_867 (
   .O(gates_552),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1100101001111100100100111001010100101011111110011101101010001100)  
) LUT6_868 (
   .O(gates_872),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0111101101001000011011110001001000000000001100001110100001111101)  
) LUT6_869 (
   .O(gates_1409),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b0111110010011100101010010100000011001001000101111110010110001010)  
) LUT6_870 (
   .O(gates_635),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0000101001011111111000011100111100011001000100001010011000100111)  
) LUT6_871 (
   .O(gates_1379),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1101111110001110010010111100110011000110011101011010101011100001)  
) LUT6_872 (
   .O(gates_366),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b0100111010101111101010111101011011001010010011000110110100010010)  
) LUT6_873 (
   .O(gates_1143),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0100110101110000111000000100010110001110001100101100101111100011)  
) LUT6_874 (
   .O(gates_533),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1010011010011001100001101101001110101001110111101000001101000010)  
) LUT6_875 (
   .O(gates_979),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0001110010101110000100011000101011011110100101011100001100011101)  
) LUT6_876 (
   .O(gates_310),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1110010001011101000111000000010100111111000101110111011111011011)  
) LUT6_877 (
   .O(gates_939),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0101100100001100111110101011001001000101011011111110010101101101)  
) LUT6_878 (
   .O(gates_150),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1100111111110110011011110100010001101000010110001011110110011010)  
) LUT6_879 (
   .O(gates_1123),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0011110011000000111100100000110111111100000110101100110011011100)  
) LUT6_880 (
   .O(gates_1404),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0110011011111111011100100111011111001000110010100010110101100110)  
) LUT6_881 (
   .O(gates_919),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0001100110010000000111001111110111010100101010001000011000001000)  
) LUT6_882 (
   .O(gates_445),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0001101010001000101010101001010000111101001111111101001010101111)  
) LUT6_883 (
   .O(gates_300),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0010111001101111101101010010011111110110010010111011110000100110)  
) LUT6_884 (
   .O(gates_1190),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0010111000010111011000001100111011110111011101001001101001010111)  
) LUT6_885 (
   .O(gates_1126),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0101101010111000100001101010101010001010010000011000001101110010)  
) LUT6_886 (
   .O(gates_1229),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1111111001000111001111001111110100011000000101000011010111100110)  
) LUT6_887 (
   .O(gates_1235),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0111111100111000001010111110101100010001101011010101111110001110)  
) LUT6_888 (
   .O(gates_1013),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0000100100001111110100000010011011011010110010001011001100101001)  
) LUT6_889 (
   .O(gates_741),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0011011101001001001100000110010010001000111000001111110100101101)  
) LUT6_890 (
   .O(gates_873),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1000111001001111011100111101100100110101111011001100000110100001)  
) LUT6_891 (
   .O(gates_318),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1101101111111100000000011111111111010011101000110110000001011000)  
) LUT6_892 (
   .O(gates_786),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0010001000011110111101001001011011110111011111101010011111011110)  
) LUT6_893 (
   .O(gates_696),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0010010001100001100111111111100011100110111010111011011011011000)  
) LUT6_894 (
   .O(gates_969),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0101111111100110111101000110110001000110111000000011001111000010)  
) LUT6_895 (
   .O(gates_1168),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1010001001110011110001111100111100111011100010111010100100010100)  
) LUT6_896 (
   .O(gates_1275),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1111111110010110001010101111011001111000000100001111000101000010)  
) LUT6_897 (
   .O(gates_1470),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0100000100011110101100100001011000011101011100111100010101001110)  
) LUT6_898 (
   .O(gates_168),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0111000000111111111111011000111100100000101001011100011010010101)  
) LUT6_899 (
   .O(gates_521),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0100100000010100001011111000111010110100000001011100110111111100)  
) LUT6_900 (
   .O(gates_1080),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0000011011110100000011110000101111111101100101011100010110011111)  
) LUT6_901 (
   .O(gates_417),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0011101101110110001001001100010001001011011000000110110011110010)  
) LUT6_902 (
   .O(gates_1413),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b1000101100001010010011110111000010100100000001111011100101000000)  
) LUT6_903 (
   .O(gates_245),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0100000101001011000001001101010001010110000101000101100010000101)  
) LUT6_904 (
   .O(gates_612),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0001001001010101000111001110110101111010100101010100010100101010)  
) LUT6_905 (
   .O(gates_1480),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1010100000111111110100011001010011011101101011001101000101110011)  
) LUT6_906 (
   .O(gates_688),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1001000001110101000010000011000000100010010101011110010101111010)  
) LUT6_907 (
   .O(gates_679),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1001011010000100101011110001111010110100110100100001000111110001)  
) LUT6_908 (
   .O(gates_473),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b0111000010010101101011111001100101001101001010110100111111110011)  
) LUT6_909 (
   .O(gates_603),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0110101010111011010010010111111100101100010101101010001110010110)  
) LUT6_910 (
   .O(gates_1088),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0110100100001110110100111010101101010001100010000000110010010110)  
) LUT6_911 (
   .O(gates_692),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0011000111010001010100011000100011111110110010000010001111111100)  
) LUT6_912 (
   .O(gates_819),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1001110111101010101000110000011011101001100110011000011011110011)  
) LUT6_913 (
   .O(gates_928),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1100001111010110100101011110000110011100100000000010100101011101)  
) LUT6_914 (
   .O(gates_1484),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1000101001001101000101110001000001111001100010111100001000010110)  
) LUT6_915 (
   .O(gates_1274),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1011100010001001001000111000001010111101100001101110110101011111)  
) LUT6_916 (
   .O(gates_1187),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b1011111100101110011011010000011011011000011010111111011010010000)  
) LUT6_917 (
   .O(gates_809),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0011111101010010101111111100011010010011010000111000111010100101)  
) LUT6_918 (
   .O(gates_1202),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b1011110111100011101000001011010010111000010111001001101110000011)  
) LUT6_919 (
   .O(gates_763),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0111100011101000010000101110011010100101110110001010101010101000)  
) LUT6_920 (
   .O(gates_358),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b1011111111110010001101100101000101110010111000000101101100110101)  
) LUT6_921 (
   .O(gates_1059),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1100101010101101101000000101001111000011000010101010100001101100)  
) LUT6_922 (
   .O(gates_1423),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0001101100100010001101001000010101100011100110010010001111100011)  
) LUT6_923 (
   .O(gates_1169),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1101011111001011010010111100011110110000011110111110000110010000)  
) LUT6_924 (
   .O(gates_627),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0011000011011010110010011000000100001100011100010110011111011000)  
) LUT6_925 (
   .O(gates_75),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1010010010101010011001010010011010011000010110100010010000011010)  
) LUT6_926 (
   .O(gates_123),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0111000110100001000101010110100001101011010110100110110000001001)  
) LUT6_927 (
   .O(gates_734),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b1001000000100010110010110010010010111100001001000100001100110101)  
) LUT6_928 (
   .O(gates_829),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b1010000111011000101010110111011001010001011111010110010011111110)  
) LUT6_929 (
   .O(gates_773),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0101001111111010111100111000000001100100001100101011110100111111)  
) LUT6_930 (
   .O(gates_365),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0000010101001110101101011100001010111110001001110001011000111011)  
) LUT6_931 (
   .O(gates_1372),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b1111001100111000101011101100001110101001001101111001001111001001)  
) LUT6_932 (
   .O(gates_1356),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0111100101001111011110011101101110000001111001110100011000111100)  
) LUT6_933 (
   .O(gates_1205),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0110110000110000010001000101101110000011010111100001101001110000)  
) LUT6_934 (
   .O(gates_131),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b0100000000100111101001110011001100100110111100101100000110000100)  
) LUT6_935 (
   .O(gates_253),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1110100001011011111001100001001111110111010001100110001100000110)  
) LUT6_936 (
   .O(gates_995),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0010110110000110110101110011110010001010010001001110001100011010)  
) LUT6_937 (
   .O(gates_907),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1100010000011111010010010111000010110001011110110011010010000001)  
) LUT6_938 (
   .O(gates_184),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1111001011011010010000111011001100100101010100011010100000010100)  
) LUT6_939 (
   .O(gates_1144),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0011000110111011001001000010011110011010100011110111011111100000)  
) LUT6_940 (
   .O(gates_818),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0010101110000011111111110011001111111000001101000000101000111011)  
) LUT6_941 (
   .O(gates_1439),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1011001111010110110111010100100101010000110010101100110111101010)  
) LUT6_942 (
   .O(gates_1497),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1010111011001011110110010101110111101111000001101010010101110111)  
) LUT6_943 (
   .O(gates_1112),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1010001010011011001011111000010000111111110100000011011111110001)  
) LUT6_944 (
   .O(gates_23),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0010001110001011011011000101011001010011011011010110011000111001)  
) LUT6_945 (
   .O(gates_771),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b1011111100111111111011000010100001110010100101100111011011111010)  
) LUT6_946 (
   .O(gates_788),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1100011111011000001111010001111110111010110001011110111110101111)  
) LUT6_947 (
   .O(gates_1336),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1110110101100101110111000000110010001011001110111001100001111110)  
) LUT6_948 (
   .O(gates_1486),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0111101011010110010110000011100010000001101000001111110010100011)  
) LUT6_949 (
   .O(gates_784),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b1000101001110100111111111111101010001110010010010111110110101000)  
) LUT6_950 (
   .O(gates_817),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b1110001110011100110100010011110100001010101101010101110111101100)  
) LUT6_951 (
   .O(gates_757),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0010111101000111111110001000000001110101110110100001010100100101)  
) LUT6_952 (
   .O(gates_875),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b0011110000100000100111011111110011100000000001000111011000011100)  
) LUT6_953 (
   .O(gates_1000),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0011110001011000000000001101011011001011011000101001101011111111)  
) LUT6_954 (
   .O(gates_1124),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1111010101001110011111111110111101101101111000010010100110011000)  
) LUT6_955 (
   .O(gates_760),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1011010011100101001011000011010010101100000000110001110010010101)  
) LUT6_956 (
   .O(gates_89),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1111001011111101101100101001101011011000111100110000000110000001)  
) LUT6_957 (
   .O(gates_986),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1000100101001101100110010111100111110001110110000101111000110001)  
) LUT6_958 (
   .O(gates_1386),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1100001101110101011000100110111011100001111111011111001110011101)  
) LUT6_959 (
   .O(gates_1460),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1000100101111010101110011110111001011001100001101101001010011100)  
) LUT6_960 (
   .O(gates_1023),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b1000010101001011100010111000110000011110110001101010101011010010)  
) LUT6_961 (
   .O(gates_360),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1010100101010101111010100011110010010110011010000000100010010001)  
) LUT6_962 (
   .O(gates_1377),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0110001010011101110011011110000100001001110111010010010010101001)  
) LUT6_963 (
   .O(gates_630),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1100100111001100001010011001111010010110100001111111011111111001)  
) LUT6_964 (
   .O(gates_878),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1011100110111011001001011001010011000100111001111100101001101000)  
) LUT6_965 (
   .O(gates_589),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1011001101000110111001011000010111011001111101100011111100001110)  
) LUT6_966 (
   .O(gates_1429),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1111111000001111101000101000110000000000001001101001100010110101)  
) LUT6_967 (
   .O(gates_1246),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1000011100100110010011101010001001101110001000010111110100100001)  
) LUT6_968 (
   .O(gates_1396),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1000111010101010010100000101110010001001100111010010101110100110)  
) LUT6_969 (
   .O(gates_967),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0110110100101101110000000100001111110000110010000100101111011001)  
) LUT6_970 (
   .O(gates_534),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0011110010101111010101100001000101010001110000001110000001111110)  
) LUT6_971 (
   .O(gates_1164),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0001000100011001011010011111100111101111111011011011110011000001)  
) LUT6_972 (
   .O(gates_1392),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1110010110000000010010010110100100100000000101001101000001010100)  
) LUT6_973 (
   .O(gates_1524),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0011101001110011101001001010000110000000101100010110000101000001)  
) LUT6_974 (
   .O(gates_674),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1011000010011100111010111011000001100000010101000110111011110101)  
) LUT6_975 (
   .O(gates_1086),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0001010100001010001101101001010000010011010001011010000101011001)  
) LUT6_976 (
   .O(gates_1494),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1110110100001001010011010100000100010001101010111010111000101100)  
) LUT6_977 (
   .O(gates_1552),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1101110101011110011101000111001100001011111100110000010010001010)  
) LUT6_978 (
   .O(gates_154),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1110011001100000001001001001001000010110000110110101000000010110)  
) LUT6_979 (
   .O(gates_1348),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0010011011010011100011000001011101100000001101100111001101011110)  
) LUT6_980 (
   .O(gates_1140),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0001011010000001011111111000110110010101100010011101111000000011)  
) LUT6_981 (
   .O(gates_1129),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b1101000111000110000011101101101101100011101111001001010001100011)  
) LUT6_982 (
   .O(gates_234),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b0101001011110001011101000010000000101010101110110100011101001101)  
) LUT6_983 (
   .O(gates_1149),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1111001011110100010110010010000101011011101000101001110000110111)  
) LUT6_984 (
   .O(gates_615),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0101011101001100111100101001111010111111011001110010111101110100)  
) LUT6_985 (
   .O(gates_1453),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1111111100011100111010011011111100001001111011000101001010011110)  
) LUT6_986 (
   .O(gates_1456),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1001101001001100011000111001011100101101001010101001111010010100)  
) LUT6_987 (
   .O(gates_325),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0110111101000110101010100011100110101000101101100111001110001000)  
) LUT6_988 (
   .O(gates_402),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b0101101100110100001100100100101000000100101111100101110011100010)  
) LUT6_989 (
   .O(gates_1378),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0010101110101100100111101010000100101010001101100001110110100110)  
) LUT6_990 (
   .O(gates_44),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0111110000000000101010010110110000111100000000100000011101011111)  
) LUT6_991 (
   .O(gates_911),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1101101000111100110000000100011000110111011000110000101010111100)  
) LUT6_992 (
   .O(gates_26),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b0110110100001001110100110100110010001111000001011000010100101001)  
) LUT6_993 (
   .O(gates_1107),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010101101010100010110111010101101111000000010010111100111110101)  
) LUT6_994 (
   .O(gates_1218),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0010110000000000001100101110111000100100001111100010100011010100)  
) LUT6_995 (
   .O(gates_965),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1100111110101100000101111100101000010011010001011000011001110001)  
) LUT6_996 (
   .O(gates_1049),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b1111101001100000110010111111011000010110110101111101011111011000)  
) LUT6_997 (
   .O(gates_1322),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1100010000100000010111000101101100101100110011111100110110001000)  
) LUT6_998 (
   .O(gates_321),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b1111001000110101010111111100101000111101100101010001010110010100)  
) LUT6_999 (
   .O(gates_227),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1000010000001001001000111010100100110111111100001001100000100100)  
) LUT6_1000 (
   .O(gates_543),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b0100110010010000011011111101110011010101010000010111010110111100)  
) LUT6_1001 (
   .O(gates_1),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b0010011111001000110010011110010101010110010110110001011110101111)  
) LUT6_1002 (
   .O(gates_749),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1110001000100110101010000010110011110101000001101000011011011110)  
) LUT6_1003 (
   .O(gates_438),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1010001100101010000101110011110001111000101011010110011001010100)  
) LUT6_1004 (
   .O(gates_1384),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1001010010101011101010011100000100111110111010111011100000000010)  
) LUT6_1005 (
   .O(gates_413),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010110001110010100010111001011000001110011001000001010101010011)  
) LUT6_1006 (
   .O(gates_492),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1001010111001001010110100000110011100110100100100111010101010010)  
) LUT6_1007 (
   .O(gates_770),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0110010000000110101001011101111101101010000110011111110001100000)  
) LUT6_1008 (
   .O(gates_482),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1010000000011001001111110101110001011001011101110011001010101011)  
) LUT6_1009 (
   .O(gates_1410),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1111110010111101101011000001101000011010000010111100101011111001)  
) LUT6_1010 (
   .O(gates_891),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0001101001110100100111110100010100010111101010110100111001001001)  
) LUT6_1011 (
   .O(gates_1321),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b0000001110110000100010101000111010100100101111010001100011011100)  
) LUT6_1012 (
   .O(gates_146),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0111001010111100011101000011010001011110010101101000110010110110)  
) LUT6_1013 (
   .O(gates_1329),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0001100110000001011111101101111111010111011111100101100000101111)  
) LUT6_1014 (
   .O(gates_898),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0011101011011000111100001000110101100101100111000001110000010001)  
) LUT6_1015 (
   .O(gates_950),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0101100110111011000001100100000101110001111011101110111010110010)  
) LUT6_1016 (
   .O(gates_947),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0001110101110100101011001011011100100110110001111000010111010011)  
) LUT6_1017 (
   .O(gates_1323),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1001001111111110101010111111001011111000100000101001000011100001)  
) LUT6_1018 (
   .O(gates_954),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b1100000000100101000101110111010111010100110100010111111000101111)  
) LUT6_1019 (
   .O(gates_1269),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1100100011111101100100110011011100011110000101110111111001011001)  
) LUT6_1020 (
   .O(gates_388),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0000101000110111000111100100110101010000001100001000110000010000)  
) LUT6_1021 (
   .O(gates_370),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b0011000011001110011101101011110010011001001100001111110000001000)  
) LUT6_1022 (
   .O(gates_814),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1011111111000100001010001000001111011111101110000000001111001100)  
) LUT6_1023 (
   .O(gates_846),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0001000001100000100110101101010100000011100011110010001110000111)  
) LUT6_1024 (
   .O(gates_1431),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b1101100101111111111011110001110010011000111110000001101110110001)  
) LUT6_1025 (
   .O(gates_204),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1001110000110111111010110001101110111000100001110011010111111111)  
) LUT6_1026 (
   .O(gates_900),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b1110100111110101111010001101101000110010111100111110000000000010)  
) LUT6_1027 (
   .O(gates_213),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0101100010010001100000101111110111011011101100110000101000000010)  
) LUT6_1028 (
   .O(gates_237),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0000000110010011101000001011010110000101101000000101000000101001)  
) LUT6_1029 (
   .O(gates_577),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1100101001000011010001001110011101101110011000111100100101110010)  
) LUT6_1030 (
   .O(gates_1224),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1101110000011000000010001110101100000011110000010011100110110101)  
) LUT6_1031 (
   .O(gates_272),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1001001010011110000100010101000000011000000101110001100111001111)  
) LUT6_1032 (
   .O(gates_574),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b1101111111111100110100000011100110001011100111000100000011001101)  
) LUT6_1033 (
   .O(gates_1044),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0111011001001001101110110110100001100111100100101100001101110011)  
) LUT6_1034 (
   .O(gates_250),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b0001011110000011000100011101010000110111011001101111101111100011)  
) LUT6_1035 (
   .O(gates_120),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b0010001000000000011110101110000110011001001100110111011100110011)  
) LUT6_1036 (
   .O(gates_1441),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0110001111101010111010011101000101011111010110001000111101101000)  
) LUT6_1037 (
   .O(gates_1167),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1001000100010010010000110101000011010100111110010010101011111110)  
) LUT6_1038 (
   .O(gates_732),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0011000010001000001100011010000000010001000101100000010110011000)  
) LUT6_1039 (
   .O(gates_807),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b0111101111011111100011011000000101110111000001001101101010001011)  
) LUT6_1040 (
   .O(gates_1509),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1101011010011101101011110110111011110010000101110011001110001011)  
) LUT6_1041 (
   .O(gates_395),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0010110101111100011001100010110110000011011100000011001000000101)  
) LUT6_1042 (
   .O(gates_190),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0010101010101011100100001101000000001011011100100111000110001111)  
) LUT6_1043 (
   .O(gates_255),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b0001001101001101011001110111000001101111101101011100011100100100)  
) LUT6_1044 (
   .O(gates_1426),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0011101010001011011110111111000010111110000111001001110101110100)  
) LUT6_1045 (
   .O(gates_712),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b0111101100100110000001001011000101000001001011110010001010100000)  
) LUT6_1046 (
   .O(gates_882),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0011001100100110111011110010111011001111110101011011101100110100)  
) LUT6_1047 (
   .O(gates_1491),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0011010100100000101111001100011000100010000100100100000011010100)  
) LUT6_1048 (
   .O(gates_1142),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1101001101011110010000011100010101001011001001101111011011000110)  
) LUT6_1049 (
   .O(gates_235),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0001000010011000001110100010110010001101011100001000001001001001)  
) LUT6_1050 (
   .O(gates_1064),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0000011100000100100111110110111001010101011011100001011000100110)  
) LUT6_1051 (
   .O(gates_280),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b0110011000001101101101100011110000100010100010001011010001001110)  
) LUT6_1052 (
   .O(gates_179),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1011111010011010001101101110110101111101101100001000110010101101)  
) LUT6_1053 (
   .O(gates_140),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0010101000001100110101010011100110010101100111000001000111100001)  
) LUT6_1054 (
   .O(gates_170),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1000001110010111010110001100110110110011000100111100011000000000)  
) LUT6_1055 (
   .O(gates_367),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1110001100101010010110000110100001001101101011000001010001010111)  
) LUT6_1056 (
   .O(gates_532),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0000010011111001000111001101110010111110011111110100010110000101)  
) LUT6_1057 (
   .O(gates_855),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1110011100000100111100001100101010000100000000111001111100010111)  
) LUT6_1058 (
   .O(gates_375),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0101111100101111101001101101010101100001100110111101101001000100)  
) LUT6_1059 (
   .O(gates_638),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1110111011110001110001110101000111011001010000100110101110101000)  
) LUT6_1060 (
   .O(gates_1001),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0111000110101101100011111000100001101110111101001010011110010100)  
) LUT6_1061 (
   .O(gates_481),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b0001110010000100101010110011101111100000011111101010111010110110)  
) LUT6_1062 (
   .O(gates_65),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1110110010000111010011110100100010101111011010110000101011110100)  
) LUT6_1063 (
   .O(gates_495),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0001110001010101110010100111001001111000110110110100010100101011)  
) LUT6_1064 (
   .O(gates_1007),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1000001101001010010101011010011000110100010000101010110101101110)  
) LUT6_1065 (
   .O(gates_79),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b1001011101101111000010000110111100000001101001100000111101100101)  
) LUT6_1066 (
   .O(gates_859),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b0101111001001011110101111000100010001011011101010110000101111111)  
) LUT6_1067 (
   .O(gates_1518),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0010111001110110000011100100010011000101100111010010111011101001)  
) LUT6_1068 (
   .O(gates_260),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1111101101100101101111011110100001111011101010010101001101101001)  
) LUT6_1069 (
   .O(gates_129),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0001111100100000001100000010010111110111000010001110000000011001)  
) LUT6_1070 (
   .O(gates_361),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1010110010010010001000010001110000010001110000010111010100100000)  
) LUT6_1071 (
   .O(gates_1278),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0011001111010111110001011101111011110100010111111001111111011101)  
) LUT6_1072 (
   .O(gates_923),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1011011110001011000011011011011110000111100011001011100100101010)  
) LUT6_1073 (
   .O(gates_1022),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b1011001010000111011001010000111110110111110010010111110000100111)  
) LUT6_1074 (
   .O(gates_718),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1010011011010001100111100000001010011110001000011001110011010000)  
) LUT6_1075 (
   .O(gates_1008),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0000110101101011010110110011110100000010001110010111010101111110)  
) LUT6_1076 (
   .O(gates_653),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1100111110011010000000011010111100000100101110011001010011001100)  
) LUT6_1077 (
   .O(gates_32),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0000111110000101100000110010101101011111011011110010101001110000)  
) LUT6_1078 (
   .O(gates_1184),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1000101111100011110000001100000101011011111101101001001101001111)  
) LUT6_1079 (
   .O(gates_657),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b0011010100101011010011110010101111100001100001111000001000110110)  
) LUT6_1080 (
   .O(gates_66),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0010010110101110011011001011010010111001110000111000100100100110)  
) LUT6_1081 (
   .O(gates_790),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b0101010101001011100100011010011111010010111110110111101001111010)  
) LUT6_1082 (
   .O(gates_614),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1100111010000000000101111100100000101101110010001001001110110110)  
) LUT6_1083 (
   .O(gates_980),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0010100001101001000100100111000001100101111011111000111011001001)  
) LUT6_1084 (
   .O(gates_36),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b1001011111010111100000110000110110101111010010011011000010010111)  
) LUT6_1085 (
   .O(gates_100),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b1100110101111011111001101011001111010111111101000010100000000011)  
) LUT6_1086 (
   .O(gates_453),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b0111010001010001011000101111000011100011011010010011111010010111)  
) LUT6_1087 (
   .O(gates_38),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1011100101100001111000111101101011001011010000110101111010001110)  
) LUT6_1088 (
   .O(gates_1214),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1000001000100110010100110110100010110010110010010011110011010100)  
) LUT6_1089 (
   .O(gates_45),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0011000010001001110110110011101011100101000100110110100100011000)  
) LUT6_1090 (
   .O(gates_1345),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b0011001110110110001001101010100010010111011100011010101010011010)  
) LUT6_1091 (
   .O(gates_278),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b0100000010000100110110110110101111110001101111010110110000011111)  
) LUT6_1092 (
   .O(gates_800),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0011001001111100000101110001011101100000110111111011110000011111)  
) LUT6_1093 (
   .O(gates_1546),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1000000010110001000010000011101000110101000100101101001001000010)  
) LUT6_1094 (
   .O(gates_759),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b0011001111100101010010000111111100101011011101011000010010011010)  
) LUT6_1095 (
   .O(gates_820),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0011001011001111110100010101011110001100101000101101000101010110)  
) LUT6_1096 (
   .O(gates_1071),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1010101011100000001100000100010011110010010110101010000110011111)  
) LUT6_1097 (
   .O(gates_943),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1110010000011011010010100011011101101100001110100011000101101010)  
) LUT6_1098 (
   .O(gates_399),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b0001011101101111100101110100000110111111101111010011001110110111)  
) LUT6_1099 (
   .O(gates_743),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1101010001110010111010101101101110011111010000011000011000011010)  
) LUT6_1100 (
   .O(gates_568),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1011100101001001010000110011100011001011010010111101100001000101)  
) LUT6_1101 (
   .O(gates_1374),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b0101101000101110011000100010011011111100110111000010011011110001)  
) LUT6_1102 (
   .O(gates_509),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1010110000110110110110000011111001011000110000010101101110110101)  
) LUT6_1103 (
   .O(gates_1109),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b1101011111001111010101110100010100110100000001001000010000110110)  
) LUT6_1104 (
   .O(gates_1166),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0001101100000010001011100110010110001110010000000000010101011110)  
) LUT6_1105 (
   .O(gates_451),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b0001011101100011100111110011111010011010111101111111010000111101)  
) LUT6_1106 (
   .O(gates_539),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b1101010000001010010111101001110101110011001101101111101011100110)  
) LUT6_1107 (
   .O(gates_1019),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1010110100010111000001001000100100111110010111111101000010101011)  
) LUT6_1108 (
   .O(gates_393),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0011001010101010111101010110000001010101101101110101110001001010)  
) LUT6_1109 (
   .O(gates_222),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b0001111001011010000000010010000111110000001100110111000110101100)  
) LUT6_1110 (
   .O(gates_753),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b1000000001011001011101100001011011011000001111111101101010100100)  
) LUT6_1111 (
   .O(gates_1057),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b1111001111110001000001010011110101000010001001111100000010000101)  
) LUT6_1112 (
   .O(gates_396),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0001000110000011001010001000010111100111010001100001101110011001)  
) LUT6_1113 (
   .O(gates_133),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1100111110101101111011111001110111001111000110001100010001010101)  
) LUT6_1114 (
   .O(gates_351),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0100000011100000100000011000100000011011100100010010011101111001)  
) LUT6_1115 (
   .O(gates_689),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b0111101010010011001110000011111001000000100111011011000000111100)  
) LUT6_1116 (
   .O(gates_1159),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0011001111111001000100011011101100010111110011011111001010101111)  
) LUT6_1117 (
   .O(gates_933),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1001011111010100001011000111110001001001011101011101110111010000)  
) LUT6_1118 (
   .O(gates_1037),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b0001100001001111011000100110011110111001110101010000001101000111)  
) LUT6_1119 (
   .O(gates_1236),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b1010010010111001000110111010101100111010111000110001010000000001)  
) LUT6_1120 (
   .O(gates_1350),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0011101111100100100010000110011110101001011010000001000000100101)  
) LUT6_1121 (
   .O(gates_996),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b0110001011101111000011011010000001000000010100000101011101110110)  
) LUT6_1122 (
   .O(gates_1171),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0110001000001100101100011110010001110100000110010101100010100000)  
) LUT6_1123 (
   .O(gates_317),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0000101000101110101111001011000011100110011010101111110001011000)  
) LUT6_1124 (
   .O(gates_220),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0010101110001000111101000110111001110001000001001100101101010100)  
) LUT6_1125 (
   .O(gates_797),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b1010000100011100110010101111111100000011001000101100111010000010)  
) LUT6_1126 (
   .O(gates_598),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1011010000011101000111110110001001111100100001001001001010111001)  
) LUT6_1127 (
   .O(gates_1111),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b1110110001001100101100010001001011011101101011000001010110000101)  
) LUT6_1128 (
   .O(gates_122),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0111011000010101101111011001111111100101110011111111010110000100)  
) LUT6_1129 (
   .O(gates_390),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b1011110000010110001001001100001001110000010110101111010111010000)  
) LUT6_1130 (
   .O(gates_970),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1000111101001111101011000101001111010010101010001000111011110110)  
) LUT6_1131 (
   .O(gates_810),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1000010100001010101111010111110111001111110010000001011000100100)  
) LUT6_1132 (
   .O(gates_307),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b0000101110000101011100110111011100110011111111001111110110011100)  
) LUT6_1133 (
   .O(gates_739),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1110111111001100101001100000101101110101011011010001011101100010)  
) LUT6_1134 (
   .O(gates_1300),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b1000101001111000001000001110010111010001110000000010101101001001)  
) LUT6_1135 (
   .O(gates_778),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1111001010000010100001010100000110011100100000011100101010100110)  
) LUT6_1136 (
   .O(gates_383),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b1000010111110001100111000011000000000110111111110111011100101000)  
) LUT6_1137 (
   .O(gates_1492),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0001000110111011100000010101000000110010110010000101111011111011)  
) LUT6_1138 (
   .O(gates_1194),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b1010110110110110000000101011001111110111100001011010011111011111)  
) LUT6_1139 (
   .O(gates_591),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b0101101001100110100000011000100001100001010100111101000100110001)  
) LUT6_1140 (
   .O(gates_22),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b1001010110011100101101000101111111011100111100110010100100110100)  
) LUT6_1141 (
   .O(gates_1263),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b1101010011111011011100111111010010001011101001100110101100111001)  
) LUT6_1142 (
   .O(gates_955),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0000001110101011000010011001011111011110110010010110101010110011)  
) LUT6_1143 (
   .O(gates_11),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b1100101110111111110010011111011001100001001101100011000001000001)  
) LUT6_1144 (
   .O(gates_566),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1101111000110111101110011010001010101101101011100111101010100101)  
) LUT6_1145 (
   .O(gates_1197),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b1110110101000100001111110001001100100101110001111000110011010011)  
) LUT6_1146 (
   .O(gates_496),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b0111001101000100111100110110101001001111001100011001111100001001)  
) LUT6_1147 (
   .O(gates_169),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1101010110110010011001000001011001011001001110100011111010010010)  
) LUT6_1148 (
   .O(gates_459),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b0010001011110010010101010000111111101110110101101111001011111011)  
) LUT6_1149 (
   .O(gates_664),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b1010110001000110100100101010001000011011000000100101011001110101)  
) LUT6_1150 (
   .O(gates_1268),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1101100101001011111111000101011101011001111101111110010001010011)  
) LUT6_1151 (
   .O(gates_1400),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b0010110011111110000010010011110101100101010100111110001010001001)  
) LUT6_1152 (
   .O(gates_107),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0100001111111001011010000011000100100010001110101010100101111011)  
) LUT6_1153 (
   .O(gates_756),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1000011011010101000001000000011100001001000110101111110111110110)  
) LUT6_1154 (
   .O(gates_305),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b0011001100010010100001001001100010101000111100101001111010111001)  
) LUT6_1155 (
   .O(gates_617),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b1101001101011111111110000110100001001101000100010110101111001101)  
) LUT6_1156 (
   .O(gates_1195),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b1001111000010101110110001111110100100101001100010010010111011111)  
) LUT6_1157 (
   .O(gates_839),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1010010001001101000111111100100010001001110011111101101100110000)  
) LUT6_1158 (
   .O(gates_424),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b1011000010111111001011000001000001010001010111101110010101011010)  
) LUT6_1159 (
   .O(gates_463),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b1111101100000010000001010000011100010001100011000111101100110100)  
) LUT6_1160 (
   .O(gates_276),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1010011110011100011011100111111010011011001100010000001100111100)  
) LUT6_1161 (
   .O(gates_597),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0111001010100101110111111111110011000011110000000111111110000111)  
) LUT6_1162 (
   .O(gates_1082),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1011110110010111110110100110100001010010100000110010010000010001)  
) LUT6_1163 (
   .O(gates_1113),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b1100011101111010000000111011011101110101000100010000011010001101)  
) LUT6_1164 (
   .O(gates_1555),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b1011001111101110000111010011011000101000100100100101000110010100)  
) LUT6_1165 (
   .O(gates_1331),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b1101000011110111001011010000110011000111101111011010100110010110)  
) LUT6_1166 (
   .O(gates_1310),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b1010001011101110000110101110011001100101010010101010100101001000)  
) LUT6_1167 (
   .O(gates_1021),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b0111011110001111111001001011111011010010000111111111101000001011)  
) LUT6_1168 (
   .O(gates_1365),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b1011100000101010000010001000010110110110011100000111101001010110)  
) LUT6_1169 (
   .O(gates_484),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0010111101011000111010001000110110110011100010000110111010101110)  
) LUT6_1170 (
   .O(gates_913),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b0001111001101001011001110101110000111011000111111111101011110010)  
) LUT6_1171 (
   .O(gates_389),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b1110000011000101111000111000001111100101000100110101110110010000)  
) LUT6_1172 (
   .O(gates_1373),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b1001110101001001010101001111010010100111010100100101001110111101)  
) LUT6_1173 (
   .O(gates_1258),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0110010101000001111001110100010010011110111010110110000001111111)  
) LUT6_1174 (
   .O(gates_1154),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b1110011110000111011100100000011001100100010011100000101010010001)  
) LUT6_1175 (
   .O(gates_705),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100010001111011010110001111101010101011100000111100000010111000)  
) LUT6_1176 (
   .O(gates_1543),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b0111011111110110101001101000110110011011010111110101010100110111)  
) LUT6_1177 (
   .O(gates_328),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1110110111011101101000001110000010010001011001000011010110011010)  
) LUT6_1178 (
   .O(gates_1036),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b0011110101000000111000011000111011011011010000010011100111000010)  
) LUT6_1179 (
   .O(gates_1158),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b0011110001000000111100101110011011011011111000000011101000111011)  
) LUT6_1180 (
   .O(gates_68),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b1100111010111000011110111111011010010000000111011100101001100001)  
) LUT6_1181 (
   .O(gates_584),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0100111110101101101000100010110001111100111011110110000110001111)  
) LUT6_1182 (
   .O(gates_268),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1011101110000001010111001101110101110000000010010110111010010100)  
) LUT6_1183 (
   .O(gates_1069),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b0001000100110011000010000100101101111101001110101001000000010000)  
) LUT6_1184 (
   .O(gates_1538),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b1101001100110010110000110110111000000001110011111101000000010101)  
) LUT6_1185 (
   .O(gates_1062),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b1111110011011111010101110001110101001100110111010111100110011011)  
) LUT6_1186 (
   .O(gates_30),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1101101010101111100110010000101111111011001110101111010111001001)  
) LUT6_1187 (
   .O(gates_3),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1110000010000111101101100011000110101010111011001110100001001000)  
) LUT6_1188 (
   .O(gates_201),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0110110000100010000110001110100011000000100011110110110011001010)  
) LUT6_1189 (
   .O(gates_556),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b1011010111100101111101101001101101011101001011011101111111111100)  
) LUT6_1190 (
   .O(gates_849),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b1000101101001001001010001100110101110110101111110100101101011111)  
) LUT6_1191 (
   .O(gates_311),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b0001111010000000100111010000100010111010110011100010110111010001)  
) LUT6_1192 (
   .O(gates_151),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1010010010101001001010100010101101101000101001000010110011010001)  
) LUT6_1193 (
   .O(gates_1357),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1001100011001100010010101000011110000010111011100100000111110010)  
) LUT6_1194 (
   .O(gates_1553),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1001101101110111110100000101111010001101110111001011010110101010)  
) LUT6_1195 (
   .O(gates_1264),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b1001010011000011100000011101100110111010010101001001010010000100)  
) LUT6_1196 (
   .O(gates_1078),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1111000000111011101000011001011101010111010001001110110000001011)  
) LUT6_1197 (
   .O(gates_132),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1111000100111101001100011110010000110101101011010011100111001101)  
) LUT6_1198 (
   .O(gates_832),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b1011111111100100111111111010001101000111110111110110010111110010)  
) LUT6_1199 (
   .O(gates_1262),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b0110101010011000001011011000100011001111100010110011011010011010)  
) LUT6_1200 (
   .O(gates_816),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b1101101110100111011010110000001110001110101110010011010101110100)  
) LUT6_1201 (
   .O(gates_1079),
   .I0(InputBits[239]),
   .I1(InputBits[236]),
   .I2(InputBits[55]),
   .I3(InputBits[569]),
   .I4(InputBits[415]),
   .I5(InputBits[166])
);
LUT6 #(
   .INIT(64'b1100110101100011110011101001111001010000111100101101110111001101)  
) LUT6_1202 (
   .O(gates_1366),
   .I0(InputBits[197]),
   .I1(InputBits[93]),
   .I2(InputBits[492]),
   .I3(InputBits[546]),
   .I4(InputBits[350]),
   .I5(InputBits[225])
);
LUT6 #(
   .INIT(64'b0001100110110001100101111011100100111101100011101000110110001110)  
) LUT6_1203 (
   .O(gates_698),
   .I0(InputBits[265]),
   .I1(InputBits[291]),
   .I2(InputBits[352]),
   .I3(InputBits[465]),
   .I4(InputBits[442]),
   .I5(InputBits[85])
);
LUT6 #(
   .INIT(64'b1111100100111101111101011000100001001010011100100100000001011100)  
) LUT6_1204 (
   .O(gates_1273),
   .I0(InputBits[178]),
   .I1(InputBits[443]),
   .I2(InputBits[174]),
   .I3(InputBits[564]),
   .I4(InputBits[9]),
   .I5(InputBits[275])
);
LUT6 #(
   .INIT(64'b0000110001110100100111011100010000010011100100001000111110110111)  
) LUT6_1205 (
   .O(gates_641),
   .I0(InputBits[544]),
   .I1(InputBits[559]),
   .I2(InputBits[26]),
   .I3(InputBits[7]),
   .I4(InputBits[374]),
   .I5(InputBits[369])
);
LUT6 #(
   .INIT(64'b1001010111001010001000100101010101011110010110111100100110111000)  
) LUT6_1206 (
   .O(gates_427),
   .I0(InputBits[376]),
   .I1(InputBits[266]),
   .I2(InputBits[488]),
   .I3(InputBits[461]),
   .I4(InputBits[308]),
   .I5(InputBits[101])
);
LUT6 #(
   .INIT(64'b0101101100110000101101101010001101111010011010100010100100000000)  
) LUT6_1207 (
   .O(gates_642),
   .I0(InputBits[398]),
   .I1(InputBits[41]),
   .I2(InputBits[332]),
   .I3(InputBits[503]),
   .I4(InputBits[246]),
   .I5(InputBits[499])
);
LUT6 #(
   .INIT(64'b0010111110100011001010000101000101111101000101011010000000001000)  
) LUT6_1208 (
   .O(gates_88),
   .I0(InputBits[184]),
   .I1(InputBits[529]),
   .I2(InputBits[211]),
   .I3(InputBits[8]),
   .I4(InputBits[296]),
   .I5(InputBits[298])
);
LUT6 #(
   .INIT(64'b0011111001010100101000110110101111100100001101111010110011011101)  
) LUT6_1209 (
   .O(gates_1151),
   .I0(InputBits[363]),
   .I1(InputBits[98]),
   .I2(InputBits[356]),
   .I3(InputBits[230]),
   .I4(InputBits[464]),
   .I5(InputBits[445])
);
LUT6 #(
   .INIT(64'b1110011101111100100110000010100010000001100100001000100010011110)  
) LUT6_1210 (
   .O(gates_999),
   .I0(InputBits[325]),
   .I1(InputBits[473]),
   .I2(InputBits[527]),
   .I3(InputBits[233]),
   .I4(InputBits[532]),
   .I5(InputBits[65])
);
LUT6 #(
   .INIT(64'b0001111010101000001010110110010101011000101001011011111001110101)  
) LUT6_1211 (
   .O(gates_1260),
   .I0(InputBits[509]),
   .I1(InputBits[571]),
   .I2(InputBits[107]),
   .I3(InputBits[51]),
   .I4(InputBits[419]),
   .I5(InputBits[34])
);
LUT6 #(
   .INIT(64'b1010001110111101000111001000100111110011010000100001111010110011)  
) LUT6_1212 (
   .O(gates_511),
   .I0(InputBits[242]),
   .I1(InputBits[278]),
   .I2(InputBits[190]),
   .I3(InputBits[506]),
   .I4(InputBits[303]),
   .I5(InputBits[73])
);
LUT6 #(
   .INIT(64'b0010011101011111101001100011001111110000000010101010100001111010)  
) LUT6_1213 (
   .O(gates_1196),
   .I0(InputBits[346]),
   .I1(InputBits[487]),
   .I2(InputBits[406]),
   .I3(InputBits[364]),
   .I4(InputBits[189]),
   .I5(InputBits[494])
);
LUT6 #(
   .INIT(64'b1100000100010111110111100111000010011101011001000100011111100010)  
) LUT6_1214 (
   .O(gates_812),
   .I0(InputBits[81]),
   .I1(InputBits[153]),
   .I2(InputBits[2]),
   .I3(InputBits[70]),
   .I4(InputBits[191]),
   .I5(InputBits[502])
);
LUT6 #(
   .INIT(64'b1011111000011001100111100010110011000001101111010100010110111110)  
) LUT6_1215 (
   .O(gates_704),
   .I0(InputBits[132]),
   .I1(InputBits[195]),
   .I2(InputBits[359]),
   .I3(InputBits[424]),
   .I4(InputBits[307]),
   .I5(InputBits[531])
);
LUT6 #(
   .INIT(64'b0010000001100011101001001101100000101000010100110000110010000000)  
) LUT6_1216 (
   .O(gates_1280),
   .I0(InputBits[348]),
   .I1(InputBits[439]),
   .I2(InputBits[551]),
   .I3(InputBits[342]),
   .I4(InputBits[400]),
   .I5(InputBits[60])
);
LUT6 #(
   .INIT(64'b0001101100101101100011100001111010100010101010110000111000010110)  
) LUT6_1217 (
   .O(gates_1075),
   .I0(InputBits[223]),
   .I1(InputBits[247]),
   .I2(InputBits[450]),
   .I3(InputBits[267]),
   .I4(InputBits[62]),
   .I5(InputBits[522])
);
LUT6 #(
   .INIT(64'b1001000001101111100000110100011010111000110101100101010111111101)  
) LUT6_1218 (
   .O(gates_1511),
   .I0(InputBits[128]),
   .I1(InputBits[386]),
   .I2(InputBits[57]),
   .I3(InputBits[537]),
   .I4(InputBits[138]),
   .I5(InputBits[29])
);
LUT6 #(
   .INIT(64'b0111011110101101001100111011010010010100100111110000110010010001)  
) LUT6_1219 (
   .O(gates_1189),
   .I0(InputBits[519]),
   .I1(InputBits[549]),
   .I2(InputBits[54]),
   .I3(InputBits[343]),
   .I4(InputBits[477]),
   .I5(InputBits[156])
);
LUT6 #(
   .INIT(64'b0000011110110000100011111000010100000101101101001100000000000000)  
) LUT6_1220 (
   .O(gates_288),
   .I0(InputBits[30]),
   .I1(InputBits[82]),
   .I2(InputBits[161]),
   .I3(InputBits[294]),
   .I4(InputBits[493]),
   .I5(InputBits[288])
);
LUT6 #(
   .INIT(64'b0111010000010010100010110011101110001100010100000111001001000010)  
) LUT6_1221 (
   .O(gates_830),
   .I0(InputBits[560]),
   .I1(InputBits[147]),
   .I2(InputBits[392]),
   .I3(InputBits[218]),
   .I4(InputBits[486]),
   .I5(InputBits[543])
);
LUT6 #(
   .INIT(64'b0110000111011111000110111000000100001010000011000100100110011110)  
) LUT6_1222 (
   .O(gates_1152),
   .I0(InputBits[123]),
   .I1(InputBits[423]),
   .I2(InputBits[212]),
   .I3(InputBits[295]),
   .I4(InputBits[129]),
   .I5(InputBits[312])
);
LUT6 #(
   .INIT(64'b1001100100111110101011001000100011110111011000101001011110011010)  
) LUT6_1223 (
   .O(gates_783),
   .I0(InputBits[431]),
   .I1(InputBits[357]),
   .I2(InputBits[169]),
   .I3(InputBits[451]),
   .I4(InputBits[505]),
   .I5(InputBits[270])
);
LUT6 #(
   .INIT(64'b0010110110011001110011010110101011100100011001011001101101100101)  
) LUT6_1224 (
   .O(gates_887),
   .I0(InputBits[305]),
   .I1(InputBits[448]),
   .I2(InputBits[286]),
   .I3(InputBits[420]),
   .I4(InputBits[414]),
   .I5(InputBits[192])
);
LUT6 #(
   .INIT(64'b0100010000001100011001011000111000011110101001110010101110100101)  
) LUT6_1225 (
   .O(gates_1004),
   .I0(InputBits[64]),
   .I1(InputBits[541]),
   .I2(InputBits[227]),
   .I3(InputBits[77]),
   .I4(InputBits[557]),
   .I5(InputBits[15])
);
LUT6 #(
   .INIT(64'b0110111111010010100100101011110010100101101100011111000000110011)  
) LUT6_1226 (
   .O(gates_909),
   .I0(InputBits[163]),
   .I1(InputBits[426]),
   .I2(InputBits[550]),
   .I3(InputBits[287]),
   .I4(InputBits[360]),
   .I5(InputBits[525])
);
LUT6 #(
   .INIT(64'b1000010010110010000110100011111000111011100001110110010010011011)  
) LUT6_1227 (
   .O(gates_73),
   .I0(InputBits[112]),
   .I1(InputBits[105]),
   .I2(InputBits[170]),
   .I3(InputBits[38]),
   .I4(InputBits[13]),
   .I5(InputBits[256])
);
LUT6 #(
   .INIT(64'b1110100010100100010001100000110100111111011010111111001001101010)  
) LUT6_1228 (
   .O(gates_1287),
   .I0(InputBits[371]),
   .I1(InputBits[449]),
   .I2(InputBits[28]),
   .I3(InputBits[45]),
   .I4(InputBits[530]),
   .I5(InputBits[413])
);
LUT6 #(
   .INIT(64'b1011000101110111001101111000100001010000111011101101100101101110)  
) LUT6_1229 (
   .O(gates_827),
   .I0(InputBits[299]),
   .I1(InputBits[164]),
   .I2(InputBits[338]),
   .I3(InputBits[199]),
   .I4(InputBits[508]),
   .I5(InputBits[50])
);
LUT6 #(
   .INIT(64'b1110111001000110110000011010001100000001001010100011001101010110)  
) LUT6_1230 (
   .O(gates_372),
   .I0(InputBits[124]),
   .I1(InputBits[251]),
   .I2(InputBits[315]),
   .I3(InputBits[556]),
   .I4(InputBits[304]),
   .I5(InputBits[395])
);
LUT6 #(
   .INIT(64'b0111011000101011011101011010011001000001010101111101001110110100)  
) LUT6_1231 (
   .O(gates_1407),
   .I0(InputBits[281]),
   .I1(InputBits[111]),
   .I2(InputBits[355]),
   .I3(InputBits[397]),
   .I4(InputBits[327]),
   .I5(InputBits[347])
);
LUT6 #(
   .INIT(64'b1110011111111000111000010111110100100001000010110110010001111010)  
) LUT6_1232 (
   .O(gates_774),
   .I0(InputBits[482]),
   .I1(InputBits[372]),
   .I2(InputBits[452]),
   .I3(InputBits[446]),
   .I4(InputBits[528]),
   .I5(InputBits[471])
);
LUT6 #(
   .INIT(64'b0001100101111100110010111001111011100111000110111100010001100011)  
) LUT6_1233 (
   .O(gates_419),
   .I0(InputBits[196]),
   .I1(InputBits[481]),
   .I2(InputBits[523]),
   .I3(InputBits[219]),
   .I4(InputBits[290]),
   .I5(InputBits[453])
);
LUT6 #(
   .INIT(64'b0110011011101101110111100100001000100101100001000111011000101110)  
) LUT6_1234 (
   .O(gates_974),
   .I0(InputBits[269]),
   .I1(InputBits[173]),
   .I2(InputBits[59]),
   .I3(InputBits[221]),
   .I4(InputBits[24]),
   .I5(InputBits[106])
);
LUT6 #(
   .INIT(64'b0110110100010100010010111100110110001101100100100100010011100111)  
) LUT6_1235 (
   .O(gates_596),
   .I0(InputBits[457]),
   .I1(InputBits[539]),
   .I2(InputBits[490]),
   .I3(InputBits[405]),
   .I4(InputBits[52]),
   .I5(InputBits[514])
);
LUT6 #(
   .INIT(64'b1101001101000001010010101111001101101100011101100010111111110000)  
) LUT6_1236 (
   .O(gates_988),
   .I0(InputBits[261]),
   .I1(InputBits[574]),
   .I2(InputBits[232]),
   .I3(InputBits[254]),
   .I4(InputBits[268]),
   .I5(InputBits[108])
);
LUT6 #(
   .INIT(64'b0011111010100110000101001011110100011110011101011010110111111011)  
) LUT6_1237 (
   .O(gates_1041),
   .I0(InputBits[120]),
   .I1(InputBits[339]),
   .I2(InputBits[497]),
   .I3(InputBits[323]),
   .I4(InputBits[538]),
   .I5(InputBits[437])
);
LUT6 #(
   .INIT(64'b1101110010110100001010111001010000111011110001110111011110111010)  
) LUT6_1238 (
   .O(gates_605),
   .I0(InputBits[297]),
   .I1(InputBits[507]),
   .I2(InputBits[326]),
   .I3(InputBits[403]),
   .I4(InputBits[257]),
   .I5(InputBits[263])
);
LUT6 #(
   .INIT(64'b0011010100000100011111111011011011110111111100111110001111000001)  
) LUT6_1239 (
   .O(gates_476),
   .I0(InputBits[244]),
   .I1(InputBits[575]),
   .I2(InputBits[23]),
   .I3(InputBits[340]),
   .I4(InputBits[383]),
   .I5(InputBits[545])
);
LUT6 #(
   .INIT(64'b0000110101100010001000001000110000010100101000101000000011111100)  
) LUT6_1240 (
   .O(gates_286),
   .I0(InputBits[411]),
   .I1(InputBits[479]),
   .I2(InputBits[572]),
   .I3(InputBits[231]),
   .I4(InputBits[100]),
   .I5(InputBits[292])
);
LUT6 #(
   .INIT(64'b1111110000110011000000000000010101110011100110010010111010111001)  
) LUT6_1241 (
   .O(gates_661),
   .I0(InputBits[289]),
   .I1(InputBits[167]),
   .I2(InputBits[21]),
   .I3(InputBits[150]),
   .I4(InputBits[384]),
   .I5(InputBits[116])
);
LUT6 #(
   .INIT(64'b0010111010000000111011011101110110010111110111111111101001011011)  
) LUT6_1242 (
   .O(gates_629),
   .I0(InputBits[249]),
   .I1(InputBits[160]),
   .I2(InputBits[136]),
   .I3(InputBits[19]),
   .I4(InputBits[427]),
   .I5(InputBits[351])
);
LUT6 #(
   .INIT(64'b1110101001111111111100110110010110100101101000000000000101000101)  
) LUT6_1243 (
   .O(gates_772),
   .I0(InputBits[353]),
   .I1(InputBits[32]),
   .I2(InputBits[122]),
   .I3(InputBits[388]),
   .I4(InputBits[272]),
   .I5(InputBits[521])
);
LUT6 #(
   .INIT(64'b1011011000000000010111000010101100010111011110010110111001101001)  
) LUT6_1244 (
   .O(gates_646),
   .I0(InputBits[217]),
   .I1(InputBits[110]),
   .I2(InputBits[317]),
   .I3(InputBits[165]),
   .I4(InputBits[252]),
   .I5(InputBits[78])
);
LUT6 #(
   .INIT(64'b1100000000000011111110011100111000111110100001111001101010000101)  
) LUT6_1245 (
   .O(gates_1307),
   .I0(InputBits[35]),
   .I1(InputBits[14]),
   .I2(InputBits[293]),
   .I3(InputBits[235]),
   .I4(InputBits[119]),
   .I5(InputBits[171])
);
LUT6 #(
   .INIT(64'b0001110010011010001000101111100011001001010011111100010101111010)  
) LUT6_1246 (
   .O(gates_236),
   .I0(InputBits[368]),
   .I1(InputBits[72]),
   .I2(InputBits[133]),
   .I3(InputBits[143]),
   .I4(InputBits[316]),
   .I5(InputBits[381])
);
LUT6 #(
   .INIT(64'b1111100110010000011110001111001111001000010011100111000001011101)  
) LUT6_1247 (
   .O(gates_1095),
   .I0(InputBits[109]),
   .I1(InputBits[175]),
   .I2(InputBits[558]),
   .I3(InputBits[536]),
   .I4(InputBits[66]),
   .I5(InputBits[389])
);
LUT6 #(
   .INIT(64'b1010011001000000000101111110110010010010001000101100110001011001)  
) LUT6_1248 (
   .O(gates_894),
   .I0(InputBits[205]),
   .I1(InputBits[151]),
   .I2(InputBits[126]),
   .I3(InputBits[157]),
   .I4(InputBits[186]),
   .I5(InputBits[336])
);
LUT6 #(
   .INIT(64'b0010000010110111000011110101000010111110001101111110111010110111)  
) LUT6_1249 (
   .O(gates_1093),
   .I0(InputBits[214]),
   .I1(InputBits[48]),
   .I2(InputBits[102]),
   .I3(InputBits[63]),
   .I4(InputBits[37]),
   .I5(InputBits[42])
);
LUT6 #(
   .INIT(64'b1100000110000010111101101101101111010100010101110100100001010110)  
) LUT6_1250 (
   .O(gates_1483),
   .I0(InputBits[429]),
   .I1(InputBits[80]),
   .I2(InputBits[94]),
   .I3(InputBits[180]),
   .I4(InputBits[412]),
   .I5(InputBits[567])
);
LUT6 #(
   .INIT(64'b1010111101110100000001101001001000110100011101001001001011101011)  
) LUT6_1251 (
   .O(gates_364),
   .I0(InputBits[277]),
   .I1(InputBits[540]),
   .I2(InputBits[79]),
   .I3(InputBits[517]),
   .I4(InputBits[425]),
   .I5(InputBits[271])
);
LUT6 #(
   .INIT(64'b0000011101011100011110001001010101111011110111101011100111000110)  
) LUT6_1252 (
   .O(gates_1437),
   .I0(InputBits[337]),
   .I1(InputBits[409]),
   .I2(InputBits[234]),
   .I3(InputBits[361]),
   .I4(InputBits[194]),
   .I5(InputBits[16])
);
LUT6 #(
   .INIT(64'b0011101010001000110100111001100001010111101000101000100100111011)  
) LUT6_1253 (
   .O(gates_706),
   .I0(InputBits[207]),
   .I1(InputBits[69]),
   .I2(InputBits[202]),
   .I3(InputBits[255]),
   .I4(InputBits[238]),
   .I5(InputBits[542])
);
LUT6 #(
   .INIT(64'b1100100010010001000110101100010001110011110110010110101000010100)  
) LUT6_1254 (
   .O(gates_1108),
   .I0(InputBits[430]),
   .I1(InputBits[90]),
   .I2(InputBits[158]),
   .I3(InputBits[380]),
   .I4(InputBits[436]),
   .I5(InputBits[228])
);
LUT6 #(
   .INIT(64'b0101101000001111101101000000001101101011100011011101001000011010)  
) LUT6_1255 (
   .O(gates_215),
   .I0(InputBits[365]),
   .I1(InputBits[320]),
   .I2(InputBits[279]),
   .I3(InputBits[334]),
   .I4(InputBits[113]),
   .I5(InputBits[306])
);
LUT6 #(
   .INIT(64'b0000000101011011001000010100010100110011011010011110011100101110)  
) LUT6_1256 (
   .O(gates_921),
   .I0(InputBits[302]),
   .I1(InputBits[422]),
   .I2(InputBits[135]),
   .I3(InputBits[408]),
   .I4(InputBits[321]),
   .I5(InputBits[43])
);
LUT6 #(
   .INIT(64'b1111100001101110110011101001111001010110111101000010110101100110)  
) LUT6_1257 (
   .O(gates_508),
   .I0(InputBits[56]),
   .I1(InputBits[210]),
   .I2(InputBits[565]),
   .I3(InputBits[309]),
   .I4(InputBits[285]),
   .I5(InputBits[282])
);
LUT6 #(
   .INIT(64'b0110110110111101100111110100001011010011101111110011011100001010)  
) LUT6_1258 (
   .O(gates_791),
   .I0(InputBits[440]),
   .I1(InputBits[391]),
   .I2(InputBits[476]),
   .I3(InputBits[68]),
   .I4(InputBits[524]),
   .I5(InputBits[382])
);
LUT6 #(
   .INIT(64'b1001101011011110000010110100101101010101001010010100100000000100)  
) LUT6_1259 (
   .O(gates_197),
   .I0(InputBits[435]),
   .I1(InputBits[177]),
   .I2(InputBits[548]),
   .I3(InputBits[259]),
   .I4(InputBits[146]),
   .I5(InputBits[203])
);
LUT6 #(
   .INIT(64'b0001011101011011101000000010011000100001011110001111001010100111)  
) LUT6_1260 (
   .O(gates_1519),
   .I0(InputBits[193]),
   .I1(InputBits[144]),
   .I2(InputBits[341]),
   .I3(InputBits[91]),
   .I4(InputBits[331]),
   .I5(InputBits[10])
);
LUT6 #(
   .INIT(64'b0100110000010011001000101011010011000011100100010001111111110110)  
) LUT6_1261 (
   .O(gates_483),
   .I0(InputBits[155]),
   .I1(InputBits[399]),
   .I2(InputBits[515]),
   .I3(InputBits[4]),
   .I4(InputBits[500]),
   .I5(InputBits[330])
);
LUT6 #(
   .INIT(64'b0001100010111001011111000101110000001110000101100110101000011100)  
) LUT6_1262 (
   .O(gates_1395),
   .I0(InputBits[300]),
   .I1(InputBits[573]),
   .I2(InputBits[208]),
   .I3(InputBits[462]),
   .I4(InputBits[159]),
   .I5(InputBits[39])
);
LUT6 #(
   .INIT(64'b0011001110110000000000111000001000111111010110101110001110000111)  
) LUT6_1263 (
   .O(gates_811),
   .I0(InputBits[71]),
   .I1(InputBits[393]),
   .I2(InputBits[313]),
   .I3(InputBits[318]),
   .I4(InputBits[83]),
   .I5(InputBits[53])
);
LUT6 #(
   .INIT(64'b1110101101111001101110101101111011000101100111110101011100101011)  
) LUT6_1264 (
   .O(gates_1243),
   .I0(InputBits[463]),
   .I1(InputBits[97]),
   .I2(InputBits[33]),
   .I3(InputBits[229]),
   .I4(InputBits[367]),
   .I5(InputBits[11])
);
LUT6 #(
   .INIT(64'b0000101010100100001011010101100011100011000001010001100001100010)  
) LUT6_1265 (
   .O(gates_301),
   .I0(InputBits[154]),
   .I1(InputBits[162]),
   .I2(InputBits[76]),
   .I3(InputBits[563]),
   .I4(InputBits[213]),
   .I5(InputBits[432])
);
LUT6 #(
   .INIT(64'b0000110110010010000010001110010111101110101000001111010000000011)  
) LUT6_1266 (
   .O(gates_259),
   .I0(InputBits[118]),
   .I1(InputBits[27]),
   .I2(InputBits[240]),
   .I3(InputBits[396]),
   .I4(InputBits[410]),
   .I5(InputBits[183])
);
LUT6 #(
   .INIT(64'b1001111111000010011001001011001000101110000001101101101110010001)  
) LUT6_1267 (
   .O(gates_191),
   .I0(InputBits[469]),
   .I1(InputBits[472]),
   .I2(InputBits[245]),
   .I3(InputBits[416]),
   .I4(InputBits[89]),
   .I5(InputBits[570])
);
LUT6 #(
   .INIT(64'b0100001101110001101000101010101001000101001100010010000110101011)  
) LUT6_1268 (
   .O(gates_963),
   .I0(InputBits[387]),
   .I1(InputBits[87]),
   .I2(InputBits[188]),
   .I3(InputBits[394]),
   .I4(InputBits[6]),
   .I5(InputBits[418])
);
LUT6 #(
   .INIT(64'b0010110111001011010001100000110001010010011110101100001000001010)  
) LUT6_1269 (
   .O(gates_97),
   .I0(InputBits[534]),
   .I1(InputBits[434]),
   .I2(InputBits[349]),
   .I3(InputBits[134]),
   .I4(InputBits[328]),
   .I5(InputBits[47])
);
LUT6 #(
   .INIT(64'b0001010001011000000101100000001001000011000111111111011101101000)  
) LUT6_1270 (
   .O(gates_21),
   .I0(InputBits[200]),
   .I1(InputBits[322]),
   .I2(InputBits[141]),
   .I3(InputBits[58]),
   .I4(InputBits[444]),
   .I5(InputBits[460])
);
LUT6 #(
   .INIT(64'b0101111110110101001000110100010101110010011101110001100101010001)  
) LUT6_1271 (
   .O(gates_1398),
   .I0(InputBits[49]),
   .I1(InputBits[276]),
   .I2(InputBits[84]),
   .I3(InputBits[566]),
   .I4(InputBits[385]),
   .I5(InputBits[402])
);
LUT6 #(
   .INIT(64'b1100011010100010101001110110101011000110011110000101101000101011)  
) LUT6_1272 (
   .O(gates_538),
   .I0(InputBits[504]),
   .I1(InputBits[520]),
   .I2(InputBits[216]),
   .I3(InputBits[455]),
   .I4(InputBits[140]),
   .I5(InputBits[407])
);
LUT6 #(
   .INIT(64'b1000100001000010110011011110011100111100100100010101011001010110)  
) LUT6_1273 (
   .O(gates_52),
   .I0(InputBits[362]),
   .I1(InputBits[344]),
   .I2(InputBits[370]),
   .I3(InputBits[152]),
   .I4(InputBits[1]),
   .I5(InputBits[280])
);
LUT6 #(
   .INIT(64'b1001011110010101001100001101001110111110011011011111010101001101)  
) LUT6_1274 (
   .O(gates_162),
   .I0(InputBits[489]),
   .I1(InputBits[139]),
   .I2(InputBits[335]),
   .I3(InputBits[562]),
   .I4(InputBits[67]),
   .I5(InputBits[149])
);
LUT6 #(
   .INIT(64'b1011111110010100100110011100111010110110100100000111111010111100)  
) LUT6_1275 (
   .O(gates_1510),
   .I0(InputBits[40]),
   .I1(InputBits[516]),
   .I2(InputBits[375]),
   .I3(InputBits[547]),
   .I4(InputBits[95]),
   .I5(InputBits[484])
);
LUT6 #(
   .INIT(64'b1010101011011111000010100100100110000110100111010010000100100001)  
) LUT6_1276 (
   .O(gates_1020),
   .I0(InputBits[220]),
   .I1(InputBits[86]),
   .I2(InputBits[458]),
   .I3(InputBits[185]),
   .I4(InputBits[17]),
   .I5(InputBits[273])
);
LUT6 #(
   .INIT(64'b1101110011100110001111001010000110110111110101010100101000111010)  
) LUT6_1277 (
   .O(gates_506),
   .I0(InputBits[510]),
   .I1(InputBits[474]),
   .I2(InputBits[366]),
   .I3(InputBits[31]),
   .I4(InputBits[428]),
   .I5(InputBits[241])
);
LUT6 #(
   .INIT(64'b0110101001100111011000101010100101000100001111111001000000110001)  
) LUT6_1278 (
   .O(gates_876),
   .I0(InputBits[553]),
   .I1(InputBits[253]),
   .I2(InputBits[358]),
   .I3(InputBits[378]),
   .I4(InputBits[433]),
   .I5(InputBits[518])
);
LUT6 #(
   .INIT(64'b1111011111111111010000000000010101100101001110111111001001100011)  
) LUT6_1279 (
   .O(gates_302),
   .I0(InputBits[44]),
   .I1(InputBits[512]),
   .I2(InputBits[243]),
   .I3(InputBits[46]),
   .I4(InputBits[470]),
   .I5(InputBits[417])
);
LUT6 #(
   .INIT(64'b1000110000001100010000101010001101100111010011110110100000001010)  
) LUT6_1280 (
   .O(gates_194),
   .I0(InputBits[513]),
   .I1(InputBits[25]),
   .I2(InputBits[404]),
   .I3(InputBits[130]),
   .I4(InputBits[274]),
   .I5(InputBits[262])
);
LUT6 #(
   .INIT(64'b0011001100101100001000110111110100011010110001000011010011000001)  
) LUT6_1281 (
   .O(gates_717),
   .I0(InputBits[117]),
   .I1(InputBits[495]),
   .I2(InputBits[438]),
   .I3(InputBits[103]),
   .I4(InputBits[576]),
   .I5(InputBits[483])
);
LUT6 #(
   .INIT(64'b0010001011010101101001011111001101000111110111111100100111001110)  
) LUT6_1282 (
   .O(gates_621),
   .I0(InputBits[127]),
   .I1(InputBits[283]),
   .I2(InputBits[379]),
   .I3(InputBits[554]),
   .I4(InputBits[480]),
   .I5(InputBits[345])
);
LUT6 #(
   .INIT(64'b1010111111000001010110010110001010001110110001011101101100110101)  
) LUT6_1283 (
   .O(gates_724),
   .I0(InputBits[250]),
   .I1(InputBits[18]),
   .I2(InputBits[260]),
   .I3(InputBits[137]),
   .I4(InputBits[314]),
   .I5(InputBits[485])
);
LUT6 #(
   .INIT(64'b1101100100100111010100010000111001110001101001001110100000111010)  
) LUT6_1284 (
   .O(gates_267),
   .I0(InputBits[226]),
   .I1(InputBits[74]),
   .I2(InputBits[478]),
   .I3(InputBits[466]),
   .I4(InputBits[176]),
   .I5(InputBits[526])
);
LUT6 #(
   .INIT(64'b0011010100100011011110010000111100011110101110100010110001000111)  
) LUT6_1285 (
   .O(gates_74),
   .I0(InputBits[181]),
   .I1(InputBits[459]),
   .I2(InputBits[114]),
   .I3(InputBits[561]),
   .I4(InputBits[201]),
   .I5(InputBits[264])
);
LUT6 #(
   .INIT(64'b0010000010101001110001111110001010011000101110000010110001100100)  
) LUT6_1286 (
   .O(gates_545),
   .I0(InputBits[142]),
   .I1(InputBits[22]),
   .I2(InputBits[187]),
   .I3(InputBits[310]),
   .I4(InputBits[168]),
   .I5(InputBits[5])
);
LUT6 #(
   .INIT(64'b1100100011101111100010000010101000001001001111010011101001111110)  
) LUT6_1287 (
   .O(gates_125),
   .I0(InputBits[311]),
   .I1(InputBits[377]),
   .I2(InputBits[20]),
   .I3(InputBits[96]),
   .I4(InputBits[552]),
   .I5(InputBits[131])
);
LUT6 #(
   .INIT(64'b1100100001011000111110111110001011111101100011101100001011011011)  
) LUT6_1288 (
   .O(gates_834),
   .I0(InputBits[454]),
   .I1(InputBits[115]),
   .I2(InputBits[533]),
   .I3(InputBits[182]),
   .I4(InputBits[198]),
   .I5(InputBits[3])
);
LUT6 #(
   .INIT(64'b1010010010001101100100101001010111110001111001010001010011011001)  
) LUT6_1289 (
   .O(gates_379),
   .I0(InputBits[104]),
   .I1(InputBits[475]),
   .I2(InputBits[447]),
   .I3(InputBits[209]),
   .I4(InputBits[172]),
   .I5(InputBits[204])
);
LUT6 #(
   .INIT(64'b1110000101000001101110010010000111101111100011101010111110001100)  
) LUT6_1290 (
   .O(gates_1006),
   .I0(InputBits[12]),
   .I1(InputBits[301]),
   .I2(InputBits[390]),
   .I3(InputBits[421]),
   .I4(InputBits[36]),
   .I5(InputBits[121])
);
LUT6 #(
   .INIT(64'b1010001100100101110110101010101100010011011101000011111011100001)  
) LUT6_1291 (
   .O(gates_654),
   .I0(InputBits[61]),
   .I1(InputBits[248]),
   .I2(InputBits[468]),
   .I3(InputBits[206]),
   .I4(InputBits[456]),
   .I5(InputBits[125])
);
LUT6 #(
   .INIT(64'b0101001101100000100100001010110011011100001100101010110001001101)  
) LUT6_1292 (
   .O(gates_1554),
   .I0(InputBits[501]),
   .I1(InputBits[88]),
   .I2(InputBits[148]),
   .I3(InputBits[555]),
   .I4(InputBits[258]),
   .I5(InputBits[491])
);
LUT6 #(
   .INIT(64'b1111011000000110100011100100111001010011101111111101000001000001)  
) LUT6_1293 (
   .O(gates_1085),
   .I0(InputBits[498]),
   .I1(InputBits[329]),
   .I2(InputBits[441]),
   .I3(InputBits[92]),
   .I4(InputBits[215]),
   .I5(InputBits[75])
);
LUT6 #(
   .INIT(64'b1010100111110001011100000010011010110010100011111110010101111101)  
) LUT6_1294 (
   .O(gates_292),
   .I0(InputBits[401]),
   .I1(InputBits[354]),
   .I2(InputBits[496]),
   .I3(InputBits[99]),
   .I4(InputBits[237]),
   .I5(InputBits[284])
);
LUT6 #(
   .INIT(64'b0011011101110010100100111110111110100000110101101110110110000101)  
) LUT6_1295 (
   .O(gates_557),
   .I0(InputBits[319]),
   .I1(InputBits[568]),
   .I2(InputBits[373]),
   .I3(InputBits[467]),
   .I4(InputBits[179]),
   .I5(InputBits[535])
);
LUT6 #(
   .INIT(64'b1000100101110111100111000010110101111100110111111111001011001001)  
) LUT6_1296 (
   .O(gates_82),
   .I0(InputBits[145]),
   .I1(InputBits[333]),
   .I2(InputBits[511]),
   .I3(InputBits[224]),
   .I4(InputBits[222]),
   .I5(InputBits[324])
);
LUT6 #(
   .INIT(64'b0100010110111101010100011001011000011000010000101101010110100011)  
) LUT6_1297 (
   .O(gates_81),
   .I0(gates_709),
   .I1(gates_1003),
   .I2(gates_780),
   .I3(gates_1412),
   .I4(gates_124),
   .I5(gates_29)
);
LUT6 #(
   .INIT(64'b1100001000111100101111010000111110100001000101110010011110010011)  
) LUT6_1298 (
   .O(gates_1150),
   .I0(gates_1266),
   .I1(gates_76),
   .I2(gates_86),
   .I3(gates_1415),
   .I4(gates_1250),
   .I5(gates_1173)
);
LUT6 #(
   .INIT(64'b0011011110111111010001101010001010101101100010110100100110111110)  
) LUT6_1299 (
   .O(gates_216),
   .I0(gates_1352),
   .I1(gates_588),
   .I2(gates_155),
   .I3(gates_309),
   .I4(gates_1451),
   .I5(gates_1051)
);
LUT6 #(
   .INIT(64'b1001001100101001110001011011000100110011110000100110111000000101)  
) LUT6_1300 (
   .O(gates_644),
   .I0(gates_20),
   .I1(gates_527),
   .I2(gates_205),
   .I3(gates_1153),
   .I4(gates_1210),
   .I5(gates_148)
);
LUT6 #(
   .INIT(64'b1001110001010001110011010010001100000011110111010111101101010000)  
) LUT6_1301 (
   .O(gates_733),
   .I0(gates_187),
   .I1(gates_1066),
   .I2(gates_1354),
   .I3(gates_606),
   .I4(gates_160),
   .I5(gates_1334)
);
LUT6 #(
   .INIT(64'b0101000100000001110000101011001110011100100011111000101000001001)  
) LUT6_1302 (
   .O(gates_720),
   .I0(gates_1447),
   .I1(gates_1247),
   .I2(gates_656),
   .I3(gates_854),
   .I4(gates_80),
   .I5(gates_1127)
);
LUT6 #(
   .INIT(64'b0110100010011010101100010011101000000111110010110010011001111111)  
) LUT6_1303 (
   .O(gates_31),
   .I0(gates_671),
   .I1(gates_315),
   .I2(gates_226),
   .I3(gates_785),
   .I4(gates_298),
   .I5(gates_1207)
);
LUT6 #(
   .INIT(64'b1101101011100101100001110011011111111101100011101100110001011001)  
) LUT6_1304 (
   .O(gates_130),
   .I0(gates_1359),
   .I1(gates_547),
   .I2(gates_1479),
   .I3(gates_1100),
   .I4(gates_478),
   .I5(gates_69)
);
LUT6 #(
   .INIT(64'b0110101010100000111101100010101101000010001011001111100011010101)  
) LUT6_1305 (
   .O(gates_346),
   .I0(gates_1133),
   .I1(gates_1436),
   .I2(gates_270),
   .I3(gates_409),
   .I4(gates_330),
   .I5(gates_435)
);
LUT6 #(
   .INIT(64'b0110011000111101011110100010101101000110001010010001101111011001)  
) LUT6_1306 (
   .O(gates_1217),
   .I0(gates_745),
   .I1(gates_636),
   .I2(gates_183),
   .I3(gates_27),
   .I4(gates_1289),
   .I5(gates_240)
);
LUT6 #(
   .INIT(64'b0111100101011011010110000000110101111011111100011011101000110000)  
) LUT6_1307 (
   .O(gates_447),
   .I0(gates_1249),
   .I1(gates_149),
   .I2(gates_1098),
   .I3(gates_1272),
   .I4(gates_1312),
   .I5(gates_1208)
);
LUT6 #(
   .INIT(64'b0001100000100100000100111011101011001110111100101010100010000011)  
) LUT6_1308 (
   .O(gates_199),
   .I0(gates_1043),
   .I1(gates_1503),
   .I2(gates_649),
   .I3(gates_874),
   .I4(gates_888),
   .I5(gates_687)
);
LUT6 #(
   .INIT(64'b1111100110100111100110000001111101010010010101001011101011001001)  
) LUT6_1309 (
   .O(gates_1110),
   .I0(gates_1472),
   .I1(gates_1146),
   .I2(gates_180),
   .I3(gates_136),
   .I4(gates_586),
   .I5(gates_1425)
);
LUT6 #(
   .INIT(64'b1000010101011111000011000110000110101000000110011001011011101000)  
) LUT6_1310 (
   .O(gates_853),
   .I0(gates_1199),
   .I1(gates_233),
   .I2(gates_246),
   .I3(gates_456),
   .I4(gates_998),
   .I5(gates_530)
);
LUT6 #(
   .INIT(64'b0110011101111110101001101000100110001001011010101110001100010001)  
) LUT6_1311 (
   .O(gates_562),
   .I0(gates_765),
   .I1(gates_581),
   .I2(gates_1327),
   .I3(gates_1406),
   .I4(gates_711),
   .I5(gates_863)
);
LUT6 #(
   .INIT(64'b0101101000000000110010001100101101101101101101110111111110011000)  
) LUT6_1312 (
   .O(gates_410),
   .I0(gates_1476),
   .I1(gates_1304),
   .I2(gates_554),
   .I3(gates_1530),
   .I4(gates_960),
   .I5(gates_403)
);
LUT6 #(
   .INIT(64'b0001110010110010000010010111111110111110001110110111010011101000)  
) LUT6_1313 (
   .O(gates_1031),
   .I0(gates_1337),
   .I1(gates_1209),
   .I2(gates_1388),
   .I3(gates_1259),
   .I4(gates_1362),
   .I5(gates_806)
);
LUT6 #(
   .INIT(64'b1000001010101111001000001010001011100110000001101010010011100001)  
) LUT6_1314 (
   .O(gates_1061),
   .I0(gates_1387),
   .I1(gates_294),
   .I2(gates_1096),
   .I3(gates_702),
   .I4(gates_207),
   .I5(gates_775)
);
LUT6 #(
   .INIT(64'b0100110100010110100010111011000100011110011000001111011100001010)  
) LUT6_1315 (
   .O(gates_1339),
   .I0(gates_381),
   .I1(gates_432),
   .I2(gates_164),
   .I3(gates_1375),
   .I4(gates_371),
   .I5(gates_243)
);
LUT6 #(
   .INIT(64'b0010000100011101011111101101001011111110111110001000000001001000)  
) LUT6_1316 (
   .O(gates_218),
   .I0(gates_523),
   .I1(gates_261),
   .I2(gates_555),
   .I3(gates_912),
   .I4(gates_1302),
   .I5(gates_408)
);
LUT6 #(
   .INIT(64'b1000010110111110101110101011101010111110110111110010110100110101)  
) LUT6_1317 (
   .O(gates_929),
   .I0(gates_582),
   .I1(gates_12),
   .I2(gates_917),
   .I3(gates_55),
   .I4(gates_147),
   .I5(gates_971)
);
LUT6 #(
   .INIT(64'b0111000110101011011110011110001001000011000111001001011101010100)  
) LUT6_1318 (
   .O(gates_110),
   .I0(gates_672),
   .I1(gates_313),
   .I2(gates_116),
   .I3(gates_119),
   .I4(gates_166),
   .I5(gates_499)
);
LUT6 #(
   .INIT(64'b1011000111010101010100101001011000101100011101001000110111000000)  
) LUT6_1319 (
   .O(gates_1131),
   .I0(gates_1507),
   .I1(gates_297),
   .I2(gates_282),
   .I3(gates_157),
   .I4(gates_1397),
   .I5(gates_747)
);
LUT6 #(
   .INIT(64'b1110111111011011101101011100001110001001100000010110001111110100)  
) LUT6_1320 (
   .O(gates_1068),
   .I0(gates_682),
   .I1(gates_1462),
   .I2(gates_673),
   .I3(gates_1309),
   .I4(gates_993),
   .I5(gates_61)
);
LUT6 #(
   .INIT(64'b0000100011100011101000011100001110000000100000110110000011011111)  
) LUT6_1321 (
   .O(gates_601),
   .I0(gates_455),
   .I1(gates_1058),
   .I2(gates_1411),
   .I3(gates_571),
   .I4(gates_897),
   .I5(gates_1251)
);
LUT6 #(
   .INIT(64'b1010100010010011001001001100100101001101110001100100111000111110)  
) LUT6_1322 (
   .O(gates_1067),
   .I0(gates_1092),
   .I1(gates_1416),
   .I2(gates_263),
   .I3(gates_884),
   .I4(gates_319),
   .I5(gates_1267)
);
LUT6 #(
   .INIT(64'b0010010110101100011100111010101011000010101000000110011011010001)  
) LUT6_1323 (
   .O(gates_1114),
   .I0(gates_904),
   .I1(gates_327),
   .I2(gates_1271),
   .I3(gates_678),
   .I4(gates_1215),
   .I5(gates_1294)
);
LUT6 #(
   .INIT(64'b0000100110011010100001001000100110001010101000000111110101001111)  
) LUT6_1324 (
   .O(gates_628),
   .I0(gates_1385),
   .I1(gates_1118),
   .I2(gates_1522),
   .I3(gates_722),
   .I4(gates_735),
   .I5(gates_1290)
);
LUT6 #(
   .INIT(64'b0111101001101011011010100011110011111001100000101010011111010101)  
) LUT6_1325 (
   .O(gates_1132),
   .I0(gates_13),
   .I1(gates_230),
   .I2(gates_359),
   .I3(gates_1489),
   .I4(gates_326),
   .I5(gates_1493)
);
LUT6 #(
   .INIT(64'b0100101110001010101101101000011000011000000011001000110010111101)  
) LUT6_1326 (
   .O(gates_920),
   .I0(gates_1030),
   .I1(gates_501),
   .I2(gates_595),
   .I3(gates_669),
   .I4(gates_428),
   .I5(gates_16)
);
LUT6 #(
   .INIT(64'b0101101110111100000011001000111100101001110111100001001110110000)  
) LUT6_1327 (
   .O(gates_1012),
   .I0(gates_195),
   .I1(gates_1514),
   .I2(gates_1161),
   .I3(gates_1028),
   .I4(gates_1303),
   .I5(gates_474)
);
LUT6 #(
   .INIT(64'b0101100110111011000111101010011000101010011011101101000011010110)  
) LUT6_1328 (
   .O(gates_946),
   .I0(gates_1527),
   .I1(gates_1147),
   .I2(gates_50),
   .I3(gates_105),
   .I4(gates_632),
   .I5(gates_387)
);
LUT6 #(
   .INIT(64'b1110111101101111000010101101011011111000011000010101000011100110)  
) LUT6_1329 (
   .O(gates_1408),
   .I0(gates_1433),
   .I1(gates_1305),
   .I2(gates_1163),
   .I3(gates_1046),
   .I4(gates_725),
   .I5(gates_289)
);
LUT6 #(
   .INIT(64'b0001100100101111010110101010110100101001001001111001111100111000)  
) LUT6_1330 (
   .O(gates_500),
   .I0(gates_391),
   .I1(gates_522),
   .I2(gates_56),
   .I3(gates_1370),
   .I4(gates_962),
   .I5(gates_287)
);
LUT6 #(
   .INIT(64'b0011111100111011001110001010110011000000001100110111011000011001)  
) LUT6_1331 (
   .O(gates_1257),
   .I0(gates_1206),
   .I1(gates_740),
   .I2(gates_1072),
   .I3(gates_700),
   .I4(gates_949),
   .I5(gates_668)
);
LUT6 #(
   .INIT(64'b0001000111010000001011000011010010101010110010101001000001010010)  
) LUT6_1332 (
   .O(gates_266),
   .I0(gates_177),
   .I1(gates_1306),
   .I2(gates_1320),
   .I3(gates_503),
   .I4(gates_93),
   .I5(gates_1383)
);
LUT6 #(
   .INIT(64'b1111010010101110111001111101001010011101100101011111111000100101)  
) LUT6_1333 (
   .O(gates_663),
   .I0(gates_997),
   .I1(gates_1341),
   .I2(gates_19),
   .I3(gates_926),
   .I4(gates_879),
   .I5(gates_314)
);
LUT6 #(
   .INIT(64'b1111100110111001100111011100111100011101000000101111100001110001)  
) LUT6_1334 (
   .O(gates_731),
   .I0(gates_1548),
   .I1(gates_1116),
   .I2(gates_652),
   .I3(gates_422),
   .I4(gates_938),
   .I5(gates_1018)
);
LUT6 #(
   .INIT(64'b1101111111101011010101101001010101000011000011000100111010110011)  
) LUT6_1335 (
   .O(gates_271),
   .I0(gates_1245),
   .I1(gates_1549),
   .I2(gates_249),
   .I3(gates_14),
   .I4(gates_987),
   .I5(gates_457)
);
LUT6 #(
   .INIT(64'b1110111100000010101010010001010111011001001100100110011111101010)  
) LUT6_1336 (
   .O(gates_1525),
   .I0(gates_1317),
   .I1(gates_188),
   .I2(gates_881),
   .I3(gates_57),
   .I4(gates_186),
   .I5(gates_639)
);
LUT6 #(
   .INIT(64'b1110010101001100100100111011011001110110010010000100101111000010)  
) LUT6_1337 (
   .O(gates_258),
   .I0(gates_349),
   .I1(gates_750),
   .I2(gates_984),
   .I3(gates_730),
   .I4(gates_1380),
   .I5(gates_316)
);
LUT6 #(
   .INIT(64'b0010011001100101000011010110100011010111010100110010100100010010)  
) LUT6_1338 (
   .O(gates_789),
   .I0(gates_1457),
   .I1(gates_442),
   .I2(gates_1135),
   .I3(gates_625),
   .I4(gates_1461),
   .I5(gates_1089)
);
LUT6 #(
   .INIT(64'b0010011000100100100010100010000101111011111111100111011100111100)  
) LUT6_1339 (
   .O(gates_104),
   .I0(gates_450),
   .I1(gates_693),
   .I2(gates_1277),
   .I3(gates_1402),
   .I4(gates_411),
   .I5(gates_792)
);
LUT6 #(
   .INIT(64'b1100000110001110111111100101100100101101110110010100001010100110)  
) LUT6_1340 (
   .O(gates_845),
   .I0(gates_1367),
   .I1(gates_470),
   .I2(gates_1177),
   .I3(gates_1237),
   .I4(gates_531),
   .I5(gates_793)
);
LUT6 #(
   .INIT(64'b0001001100010110010001010001010000101101110000000101101101001001)  
) LUT6_1341 (
   .O(gates_802),
   .I0(gates_1346),
   .I1(gates_118),
   .I2(gates_942),
   .I3(gates_659),
   .I4(gates_798),
   .I5(gates_1270)
);
LUT6 #(
   .INIT(64'b1100001111011110100000110011101100001110100011110110001111110100)  
) LUT6_1342 (
   .O(gates_174),
   .I0(gates_824),
   .I1(gates_665),
   .I2(gates_386),
   .I3(gates_208),
   .I4(gates_1498),
   .I5(gates_406)
);
LUT6 #(
   .INIT(64'b0101100100110111100100100011010001010111100110011001101100101000)  
) LUT6_1343 (
   .O(gates_964),
   .I0(gates_587),
   .I1(gates_647),
   .I2(gates_1145),
   .I3(gates_536),
   .I4(gates_200),
   .I5(gates_404)
);
LUT6 #(
   .INIT(64'b0001100011000110101011101000000101100000100100001100001010011111)  
) LUT6_1344 (
   .O(gates_1221),
   .I0(gates_1403),
   .I1(gates_1170),
   .I2(gates_1418),
   .I3(gates_902),
   .I4(gates_357),
   .I5(gates_460)
);
LUT6 #(
   .INIT(64'b1011011000110000000111111010111001000110100000001101011001100010)  
) LUT6_1345 (
   .O(gates_737),
   .I0(gates_1299),
   .I1(gates_212),
   .I2(gates_710),
   .I3(gates_440),
   .I4(gates_648),
   .I5(gates_444)
);
LUT6 #(
   .INIT(64'b0110100110100111101001111000001001101011100010101100101100011110)  
) LUT6_1346 (
   .O(gates_1442),
   .I0(gates_1474),
   .I1(gates_269),
   .I2(gates_940),
   .I3(gates_1296),
   .I4(gates_414),
   .I5(gates_719)
);
LUT6 #(
   .INIT(64'b0010100001110011011011000100010100110110000001100100010110000001)  
) LUT6_1347 (
   .O(gates_486),
   .I0(gates_1232),
   .I1(gates_895),
   .I2(gates_2),
   .I3(gates_680),
   .I4(gates_1495),
   .I5(gates_189)
);
LUT6 #(
   .INIT(64'b0100011111100100111011010011111100001010100011010110100101110001)  
) LUT6_1348 (
   .O(gates_573),
   .I0(gates_924),
   .I1(gates_217),
   .I2(gates_48),
   .I3(gates_1038),
   .I4(gates_677),
   .I5(gates_941)
);
LUT6 #(
   .INIT(64'b0101001110010101111001000110001110011110010000011010111000010101)  
) LUT6_1349 (
   .O(gates_398),
   .I0(gates_951),
   .I1(gates_1045),
   .I2(gates_1355),
   .I3(gates_1534),
   .I4(gates_1450),
   .I5(gates_512)
);
LUT6 #(
   .INIT(64'b0011011001010010010111101001011111010111011101011110000000100000)  
) LUT6_1350 (
   .O(gates_10),
   .I0(gates_1252),
   .I1(gates_1537),
   .I2(gates_1478),
   .I3(gates_1228),
   .I4(gates_137),
   .I5(gates_223)
);
LUT6 #(
   .INIT(64'b1110100011100010010100100110101001110100110001001101100011100100)  
) LUT6_1351 (
   .O(gates_1513),
   .I0(gates_1231),
   .I1(gates_161),
   .I2(gates_63),
   .I3(gates_58),
   .I4(gates_510),
   .I5(gates_265)
);
LUT6 #(
   .INIT(64'b0000111100111100011111100010110010110100000000000111111101000001)  
) LUT6_1352 (
   .O(gates_1014),
   .I0(gates_836),
   .I1(gates_1547),
   .I2(gates_4),
   .I3(gates_1081),
   .I4(gates_1326),
   .I5(gates_485)
);
LUT6 #(
   .INIT(64'b0010111111000001000000000010110100111101010110010110000001000100)  
) LUT6_1353 (
   .O(gates_53),
   .I0(gates_622),
   .I1(gates_275),
   .I2(gates_752),
   .I3(gates_850),
   .I4(gates_462),
   .I5(gates_84)
);
LUT6 #(
   .INIT(64'b0010000011111011101110111000110001010000111000011010100001111100)  
) LUT6_1354 (
   .O(gates_1253),
   .I0(gates_906),
   .I1(gates_1042),
   .I2(gates_544),
   .I3(gates_548),
   .I4(gates_489),
   .I5(gates_1369)
);
LUT6 #(
   .INIT(64'b1001011101000110110101110010101010100111110110011011110001110110)  
) LUT6_1355 (
   .O(gates_1368),
   .I0(gates_1318),
   .I1(gates_128),
   .I2(gates_256),
   .I3(gates_1053),
   .I4(gates_401),
   .I5(gates_1330)
);
LUT6 #(
   .INIT(64'b0011111011000101110011011000111111011100011101000001100001010000)  
) LUT6_1356 (
   .O(gates_1162),
   .I0(gates_362),
   .I1(gates_1444),
   .I2(gates_1134),
   .I3(gates_866),
   .I4(gates_708),
   .I5(gates_823)
);
LUT6 #(
   .INIT(64'b0110000011100010011111111110110010110111001010111101010000010101)  
) LUT6_1357 (
   .O(gates_219),
   .I0(gates_799),
   .I1(gates_103),
   .I2(gates_1496),
   .I3(gates_341),
   .I4(gates_449),
   .I5(gates_1499)
);
LUT6 #(
   .INIT(64'b0001111010011000000011000100100011101111111101011110000010001100)  
) LUT6_1358 (
   .O(gates_71),
   .I0(gates_9),
   .I1(gates_848),
   .I2(gates_504),
   .I3(gates_412),
   .I4(gates_616),
   .I5(gates_1463)
);
LUT6 #(
   .INIT(64'b0100101101111111101000011110000110101010101110111011110011011101)  
) LUT6_1359 (
   .O(gates_604),
   .I0(gates_1344),
   .I1(gates_279),
   .I2(gates_1090),
   .I3(gates_1233),
   .I4(gates_1176),
   .I5(gates_1242)
);
LUT6 #(
   .INIT(64'b0111101000111001010100010110010000000010101010101111000101100011)  
) LUT6_1360 (
   .O(gates_910),
   .I0(gates_736),
   .I1(gates_840),
   .I2(gates_953),
   .I3(gates_870),
   .I4(gates_959),
   .I5(gates_1192)
);
LUT6 #(
   .INIT(64'b1110010001100011101001010110100001110001011000110011011000110100)  
) LUT6_1361 (
   .O(gates_472),
   .I0(gates_376),
   .I1(gates_1469),
   .I2(gates_1545),
   .I3(gates_1102),
   .I4(gates_1099),
   .I5(gates_1288)
);
LUT6 #(
   .INIT(64'b0111110101010001010111010110100001011111100101000101001111011100)  
) LUT6_1362 (
   .O(gates_1319),
   .I0(gates_248),
   .I1(gates_1504),
   .I2(gates_108),
   .I3(gates_333),
   .I4(gates_1185),
   .I5(gates_607)
);
LUT6 #(
   .INIT(64'b0110100000001100101101111111101011101011001011100111111010110011)  
) LUT6_1363 (
   .O(gates_925),
   .I0(gates_90),
   .I1(gates_363),
   .I2(gates_885),
   .I3(gates_96),
   .I4(gates_1160),
   .I5(gates_1165)
);
LUT6 #(
   .INIT(64'b0101110111100001111101100000010101011110000000010110110011111101)  
) LUT6_1364 (
   .O(gates_1227),
   .I0(gates_1060),
   .I1(gates_575),
   .I2(gates_1222),
   .I3(gates_322),
   .I4(gates_1284),
   .I5(gates_968)
);
LUT6 #(
   .INIT(64'b1000100001100111110101111110000000110100001101101100000000111011)  
) LUT6_1365 (
   .O(gates_707),
   .I0(gates_209),
   .I1(gates_835),
   .I2(gates_1512),
   .I3(gates_25),
   .I4(gates_934),
   .I5(gates_1526)
);
LUT6 #(
   .INIT(64'b1010010000101000110101100110100001000001111100000000111101010100)  
) LUT6_1366 (
   .O(gates_397),
   .I0(gates_585),
   .I1(gates_291),
   .I2(gates_609),
   .I3(gates_1009),
   .I4(gates_766),
   .I5(gates_1332)
);
LUT6 #(
   .INIT(64'b0101101010010111011111101000111111001101101101111100011110011101)  
) LUT6_1367 (
   .O(gates_1521),
   .I0(gates_1027),
   .I1(gates_340),
   .I2(gates_334),
   .I3(gates_1347),
   .I4(gates_1427),
   .I5(gates_117)
);
LUT6 #(
   .INIT(64'b0100010101000001011111001000101111001100011011100100110011011100)  
) LUT6_1368 (
   .O(gates_1301),
   .I0(gates_681),
   .I1(gates_1382),
   .I2(gates_880),
   .I3(gates_467),
   .I4(gates_982),
   .I5(gates_173)
);
LUT6 #(
   .INIT(64'b1011100010101000010110100011011001101100001100110011010110011111)  
) LUT6_1369 (
   .O(gates_407),
   .I0(gates_1482),
   .I1(gates_425),
   .I2(gates_549),
   .I3(gates_570),
   .I4(gates_153),
   .I5(gates_620)
);
LUT6 #(
   .INIT(64'b0100001011010110111000111100111000011111010011100101011010010000)  
) LUT6_1370 (
   .O(gates_1117),
   .I0(gates_1389),
   .I1(gates_1532),
   .I2(gates_5),
   .I3(gates_804),
   .I4(gates_1084),
   .I5(gates_1298)
);
LUT6 #(
   .INIT(64'b1001101010101100101100101110111001001001010110110011001001111100)  
) LUT6_1371 (
   .O(gates_1179),
   .I0(gates_1115),
   .I1(gates_583),
   .I2(gates_936),
   .I3(gates_862),
   .I4(gates_1248),
   .I5(gates_916)
);
LUT6 #(
   .INIT(64'b0101101111110000011111111110010111111011101100001111010110011001)  
) LUT6_1372 (
   .O(gates_684),
   .I0(gates_892),
   .I1(gates_1175),
   .I2(gates_1508),
   .I3(gates_631),
   .I4(gates_1438),
   .I5(gates_1539)
);
LUT6 #(
   .INIT(64'b0010101001010011010100100110010001111001000110100000010010011100)  
) LUT6_1373 (
   .O(gates_662),
   .I0(gates_1393),
   .I1(gates_1432),
   .I2(gates_382),
   .I3(gates_1443),
   .I4(gates_805),
   .I5(gates_762)
);
LUT6 #(
   .INIT(64'b0101110011100010010101000101010111011001111011010011011011100101)  
) LUT6_1374 (
   .O(gates_1047),
   .I0(gates_507),
   .I1(gates_537),
   .I2(gates_262),
   .I3(gates_1188),
   .I4(gates_1157),
   .I5(gates_78)
);
LUT6 #(
   .INIT(64'b0111100111110101110010110111001001010100111010010010000101110000)  
) LUT6_1375 (
   .O(gates_634),
   .I0(gates_1446),
   .I1(gates_563),
   .I2(gates_491),
   .I3(gates_380),
   .I4(gates_42),
   .I5(gates_808)
);
LUT6 #(
   .INIT(64'b0101000100000110010101000101010101011101010010001110110100101111)  
) LUT6_1376 (
   .O(gates_1471),
   .I0(gates_141),
   .I1(gates_600),
   .I2(gates_224),
   .I3(gates_1225),
   .I4(gates_592),
   .I5(gates_239)
);
LUT6 #(
   .INIT(64'b0110001001100011011110001111100101010001110110101010111010001110)  
) LUT6_1377 (
   .O(gates_821),
   .I0(gates_1541),
   .I1(gates_299),
   .I2(gates_374),
   .I3(gates_1465),
   .I4(gates_274),
   .I5(gates_308)
);
LUT6 #(
   .INIT(64'b0010001100010010100010001011110100101110000010000001110011101100)  
) LUT6_1378 (
   .O(gates_593),
   .I0(gates_1137),
   .I1(gates_914),
   .I2(gates_1070),
   .I3(gates_847),
   .I4(gates_1401),
   .I5(gates_945)
);
LUT6 #(
   .INIT(64'b1101010101100001000110011101100000000111101101100101000011101000)  
) LUT6_1379 (
   .O(gates_991),
   .I0(gates_172),
   .I1(gates_293),
   .I2(gates_40),
   .I3(gates_1529),
   .I4(gates_858),
   .I5(gates_1052)
);
LUT6 #(
   .INIT(64'b1001000000011011110100000111110111101101111011010000111111011111)  
) LUT6_1380 (
   .O(gates_794),
   .I0(gates_728),
   .I1(gates_869),
   .I2(gates_1220),
   .I3(gates_332),
   .I4(gates_72),
   .I5(gates_1417)
);
LUT6 #(
   .INIT(64'b1101001000001110110111011000011011001110111101100001010100101101)  
) LUT6_1381 (
   .O(gates_751),
   .I0(gates_828),
   .I1(gates_46),
   .I2(gates_1219),
   .I3(gates_1279),
   .I4(gates_932),
   .I5(gates_1293)
);
LUT6 #(
   .INIT(64'b1101001111100001110110001101000101110101101101011010100000110100)  
) LUT6_1382 (
   .O(gates_418),
   .I0(gates_115),
   .I1(gates_1104),
   .I2(gates_1077),
   .I3(gates_520),
   .I4(gates_244),
   .I5(gates_1536)
);
LUT6 #(
   .INIT(64'b1010110011011011001000001111100010101001111000000100101001011010)  
) LUT6_1383 (
   .O(gates_339),
   .I0(gates_703),
   .I1(gates_106),
   .I2(gates_1459),
   .I3(gates_1343),
   .I4(gates_324),
   .I5(gates_1286)
);
LUT6 #(
   .INIT(64'b0010100010110110110000011110001011111001011001100000001001000111)  
) LUT6_1384 (
   .O(gates_1141),
   .I0(gates_1458),
   .I1(gates_1128),
   .I2(gates_323),
   .I3(gates_102),
   .I4(gates_516),
   .I5(gates_1156)
);
LUT6 #(
   .INIT(64'b1101010011101000101000000110111000100110010111101011100101010000)  
) LUT6_1385 (
   .O(gates_1216),
   .I0(gates_1390),
   .I1(gates_214),
   .I2(gates_1148),
   .I3(gates_713),
   .I4(gates_667),
   .I5(gates_167)
);
LUT6 #(
   .INIT(64'b0101100010101111010111000001100111101011011001000110000010001010)  
) LUT6_1386 (
   .O(gates_434),
   .I0(gates_1353),
   .I1(gates_815),
   .I2(gates_825),
   .I3(gates_871),
   .I4(gates_580),
   .I5(gates_966)
);
LUT6 #(
   .INIT(64'b1110001101011001100101000011010010000010010010010100110100100010)  
) LUT6_1387 (
   .O(gates_475),
   .I0(gates_769),
   .I1(gates_1358),
   .I2(gates_886),
   .I3(gates_961),
   .I4(gates_461),
   .I5(gates_135)
);
LUT6 #(
   .INIT(64'b0000011111110011001001101110000100011101101010001101010111001000)  
) LUT6_1388 (
   .O(gates_599),
   .I0(gates_1360),
   .I1(gates_487),
   .I2(gates_1502),
   .I3(gates_1204),
   .I4(gates_1183),
   .I5(gates_1056)
);
LUT6 #(
   .INIT(64'b0101011111010111101001010101101100100110000000100001100111000101)  
) LUT6_1389 (
   .O(gates_202),
   .I0(gates_1239),
   .I1(gates_185),
   .I2(gates_1139),
   .I3(gates_225),
   .I4(gates_1105),
   .I5(gates_1048)
);
LUT6 #(
   .INIT(64'b0110011110110100010000111110111011111111001100000010101110011001)  
) LUT6_1390 (
   .O(gates_776),
   .I0(gates_1240),
   .I1(gates_1340),
   .I2(gates_1230),
   .I3(gates_715),
   .I4(gates_889),
   .I5(gates_1282)
);
LUT6 #(
   .INIT(64'b1111100010110001010110000100011010111010111000111101100110101100)  
) LUT6_1391 (
   .O(gates_1011),
   .I0(gates_152),
   .I1(gates_87),
   .I2(gates_1445),
   .I3(gates_238),
   .I4(gates_851),
   .I5(gates_561)
);
LUT6 #(
   .INIT(64'b1001010010111010000001111010110001100000111000111110000101011101)  
) LUT6_1392 (
   .O(gates_685),
   .I0(gates_62),
   .I1(gates_618),
   .I2(gates_159),
   .I3(gates_443),
   .I4(gates_416),
   .I5(gates_1313)
);
LUT6 #(
   .INIT(64'b1111011101110010111000100100010101111001001000011010100101001101)  
) LUT6_1393 (
   .O(gates_1454),
   .I0(gates_1325),
   .I1(gates_643),
   .I2(gates_70),
   .I3(gates_1292),
   .I4(gates_329),
   .I5(gates_782)
);
LUT6 #(
   .INIT(64'b1100111101000000000010111100110001011010101000110001001000110010)  
) LUT6_1394 (
   .O(gates_619),
   .I0(gates_613),
   .I1(gates_1324),
   .I2(gates_60),
   .I3(gates_145),
   .I4(gates_498),
   .I5(gates_1180)
);
LUT6 #(
   .INIT(64'b0001100110000100010000111001000011011101001000111110110111001110)  
) LUT6_1395 (
   .O(gates_594),
   .I0(gates_1364),
   .I1(gates_203),
   .I2(gates_420),
   .I3(gates_488),
   .I4(gates_1399),
   .I5(gates_85)
);
LUT6 #(
   .INIT(64'b0010011010011000101100111000011000010100111101011110101110101001)  
) LUT6_1396 (
   .O(gates_1452),
   .I0(gates_952),
   .I1(gates_181),
   .I2(gates_1186),
   .I3(gates_666),
   .I4(gates_1119),
   .I5(gates_281)
);
LUT6 #(
   .INIT(64'b0111101111011101110110001101110111110100111110100011111010000010)  
) LUT6_1397 (
   .O(gates_295),
   .I0(gates_896),
   .I1(gates_1328),
   .I2(gates_121),
   .I3(gates_1255),
   .I4(gates_655),
   .I5(gates_112)
);
LUT6 #(
   .INIT(64'b0111110111000111001000001110110111111111111011011100011001000100)  
) LUT6_1398 (
   .O(gates_347),
   .I0(gates_519),
   .I1(gates_690),
   .I2(gates_670),
   .I3(gates_471),
   .I4(gates_1002),
   .I5(gates_441)
);
LUT6 #(
   .INIT(64'b1100000010101110011011101011111000000101011111001011101000000001)  
) LUT6_1399 (
   .O(gates_787),
   .I0(gates_675),
   .I1(gates_905),
   .I2(gates_1087),
   .I3(gates_572),
   .I4(gates_1342),
   .I5(gates_957)
);
LUT6 #(
   .INIT(64'b0100010010001011111110101010110101010010100100110001100111000100)  
) LUT6_1400 (
   .O(gates_564),
   .I0(gates_973),
   .I1(gates_254),
   .I2(gates_514),
   .I3(gates_415),
   .I4(gates_640),
   .I5(gates_304)
);
LUT6 #(
   .INIT(64'b0110011110000001000110111111010010110111001101000111101000100001)  
) LUT6_1401 (
   .O(gates_1254),
   .I0(gates_421),
   .I1(gates_1083),
   .I2(gates_1063),
   .I3(gates_1026),
   .I4(gates_901),
   .I5(gates_723)
);
LUT6 #(
   .INIT(64'b1000101010100010011011011000111101010101101100111101101000011001)  
) LUT6_1402 (
   .O(gates_1174),
   .I0(gates_893),
   .I1(gates_1551),
   .I2(gates_228),
   .I3(gates_1315),
   .I4(gates_1201),
   .I5(gates_231)
);
LUT6 #(
   .INIT(64'b0100111011010001000101011101001011010000110101111110001011011110)  
) LUT6_1403 (
   .O(gates_559),
   .I0(gates_1297),
   .I1(gates_41),
   .I2(gates_477),
   .I3(gates_610),
   .I4(gates_464),
   .I5(gates_343)
);
LUT6 #(
   .INIT(64'b0001100000010100111101000110000110001001101100111010011100011100)  
) LUT6_1404 (
   .O(gates_868),
   .I0(gates_578),
   .I1(gates_1466),
   .I2(gates_1490),
   .I3(gates_624),
   .I4(gates_345),
   .I5(gates_1550)
);
LUT6 #(
   .INIT(64'b0111010001100110110000001001110010110110100010110101110101001000)  
) LUT6_1405 (
   .O(gates_1055),
   .I0(gates_852),
   .I1(gates_686),
   .I2(gates_8),
   .I3(gates_1381),
   .I4(gates_738),
   .I5(gates_683)
);
LUT6 #(
   .INIT(64'b0011010000110010011110110110011110011110010111010110010011001111)  
) LUT6_1406 (
   .O(gates_918),
   .I0(gates_542),
   .I1(gates_990),
   .I2(gates_95),
   .I3(gates_1125),
   .I4(gates_676),
   .I5(gates_944)
);
LUT6 #(
   .INIT(64'b0010111001110000101001101101010001010000010101011111100010011111)  
) LUT6_1407 (
   .O(gates_695),
   .I0(gates_277),
   .I1(gates_935),
   .I2(gates_1485),
   .I3(gates_890),
   .I4(gates_176),
   .I5(gates_729)
);
LUT6 #(
   .INIT(64'b1001001011100101100000000101001111110011011110101100101000000100)  
) LUT6_1408 (
   .O(gates_232),
   .I0(gates_196),
   .I1(gates_1391),
   .I2(gates_1376),
   .I3(gates_844),
   .I4(gates_1517),
   .I5(gates_7)
);
LUT6 #(
   .INIT(64'b0111101000111111000001100001001001010000101001111010011010010000)  
) LUT6_1409 (
   .O(gates_877),
   .I0(gates_1464),
   .I1(gates_335),
   .I2(gates_1138),
   .I3(gates_1500),
   .I4(gates_1223),
   .I5(gates_426)
);
LUT6 #(
   .INIT(64'b0101101001000111000111011101011101010010110000101100111100110001)  
) LUT6_1410 (
   .O(gates_742),
   .I0(gates_831),
   .I1(gates_493),
   .I2(gates_350),
   .I3(gates_479),
   .I4(gates_726),
   .I5(gates_1349)
);
LUT6 #(
   .INIT(64'b1011100010000010110100000100001110010110101101000001011000101011)  
) LUT6_1411 (
   .O(gates_611),
   .I0(gates_567),
   .I1(gates_99),
   .I2(gates_306),
   .I3(gates_1420),
   .I4(gates_405),
   .I5(gates_37)
);
LUT6 #(
   .INIT(64'b0000010110001110100110010111110110110000001101000101110110110110)  
) LUT6_1412 (
   .O(gates_296),
   .I0(gates_143),
   .I1(gates_490),
   .I2(gates_744),
   .I3(gates_651),
   .I4(gates_1338),
   .I5(gates_518)
);
LUT6 #(
   .INIT(64'b1001100011100110001011001101101001000110001001110011010100011010)  
) LUT6_1413 (
   .O(gates_211),
   .I0(gates_579),
   .I1(gates_1316),
   .I2(gates_1308),
   .I3(gates_1421),
   .I4(gates_975),
   .I5(gates_437)
);
LUT6 #(
   .INIT(64'b0110111000111010000111110010001010110100000110010111010101001010)  
) LUT6_1414 (
   .O(gates_284),
   .I0(gates_867),
   .I1(gates_303),
   .I2(gates_977),
   .I3(gates_290),
   .I4(gates_1405),
   .I5(gates_727)
);
LUT6 #(
   .INIT(64'b0111100111100111110001000111010001100001101000011110011011110011)  
) LUT6_1415 (
   .O(gates_1311),
   .I0(gates_1033),
   .I1(gates_192),
   .I2(gates_480),
   .I3(gates_553),
   .I4(gates_356),
   .I5(gates_1172)
);
LUT6 #(
   .INIT(64'b1111101100110101000111010110111001011000011000110010000000010010)  
) LUT6_1416 (
   .O(gates_400),
   .I0(gates_569),
   .I1(gates_247),
   .I2(gates_1295),
   .I3(gates_59),
   .I4(gates_1032),
   .I5(gates_861)
);
LUT6 #(
   .INIT(64'b0101000110000100100010111100001011111110111000011101111100101100)  
) LUT6_1417 (
   .O(gates_67),
   .I0(gates_826),
   .I1(gates_1285),
   .I2(gates_761),
   .I3(gates_1136),
   .I4(gates_1213),
   .I5(gates_385)
);
LUT6 #(
   .INIT(64'b1001111010010000011100011001101110101100000100100001001111010111)  
) LUT6_1418 (
   .O(gates_755),
   .I0(gates_320),
   .I1(gates_251),
   .I2(gates_781),
   .I3(gates_842),
   .I4(gates_505),
   .I5(gates_922)
);
LUT6 #(
   .INIT(64'b1010110101110001010011111011101100011110111111110001111000000001)  
) LUT6_1419 (
   .O(gates_777),
   .I0(gates_1091),
   .I1(gates_1212),
   .I2(gates_34),
   .I3(gates_978),
   .I4(gates_1178),
   .I5(gates_283)
);
LUT6 #(
   .INIT(64'b1101100010001101110101111010101001100010101110100100000011110001)  
) LUT6_1420 (
   .O(gates_1515),
   .I0(gates_377),
   .I1(gates_378),
   .I2(gates_541),
   .I3(gates_384),
   .I4(gates_229),
   .I5(gates_699)
);
LUT6 #(
   .INIT(64'b0010111100010001011000011111100101110001001000101111100001110001)  
) LUT6_1421 (
   .O(gates_1487),
   .I0(gates_1361),
   .I1(gates_1074),
   .I2(gates_833),
   .I3(gates_1034),
   .I4(gates_1468),
   .I5(gates_252)
);
LUT6 #(
   .INIT(64'b1010101001100010000100100011011010001101101011001111100010101011)  
) LUT6_1422 (
   .O(gates_660),
   .I0(gates_1182),
   .I1(gates_560),
   .I2(gates_28),
   .I3(gates_768),
   .I4(gates_1203),
   .I5(gates_64)
);
LUT6 #(
   .INIT(64'b1101010111110110110011100010111011011010111000000001111010100101)  
) LUT6_1423 (
   .O(gates_1276),
   .I0(gates_838),
   .I1(gates_35),
   .I2(gates_1054),
   .I3(gates_937),
   .I4(gates_1211),
   .I5(gates_342)
);
LUT6 #(
   .INIT(64'b1000110111010010100100111100100010011011111101011001000100110000)  
) LUT6_1424 (
   .O(gates_524),
   .I0(gates_1473),
   .I1(gates_111),
   .I2(gates_1477),
   .I3(gates_468),
   .I4(gates_608),
   .I5(gates_1435)
);
LUT6 #(
   .INIT(64'b0111011100100010111101001111111001111000111001100011101011111011)  
) LUT6_1425 (
   .O(gates_758),
   .I0(gates_1467),
   .I1(gates_1029),
   .I2(gates_1200),
   .I3(gates_1394),
   .I4(gates_1130),
   .I5(gates_1120)
);
LUT6 #(
   .INIT(64'b1000000000100010111001000010110100010111010011111001101010111010)  
) LUT6_1426 (
   .O(gates_650),
   .I0(gates_171),
   .I1(gates_1065),
   .I2(gates_767),
   .I3(gates_494),
   .I4(gates_144),
   .I5(gates_127)
);
LUT6 #(
   .INIT(64'b0001111010110011111110111100100101001011101101000110010000000010)  
) LUT6_1427 (
   .O(gates_1191),
   .I0(gates_701),
   .I1(gates_1181),
   .I2(gates_165),
   .I3(gates_392),
   .I4(gates_17),
   .I5(gates_565)
);
LUT6 #(
   .INIT(64'b1101110111101111100010011100000101001000011110011010001010000000)  
) LUT6_1428 (
   .O(gates_989),
   .I0(gates_748),
   .I1(gates_1440),
   .I2(gates_841),
   .I3(gates_156),
   .I4(gates_550),
   .I5(gates_198)
);
LUT6 #(
   .INIT(64'b1011111110010000101000010010001010001111000001101011101011011001)  
) LUT6_1429 (
   .O(gates_645),
   .I0(gates_1101),
   .I1(gates_864),
   .I2(gates_1449),
   .I3(gates_1005),
   .I4(gates_126),
   .I5(gates_1226)
);
LUT6 #(
   .INIT(64'b1010100101010000101000011110111001101010011010101010101000000110)  
) LUT6_1430 (
   .O(gates_431),
   .I0(gates_369),
   .I1(gates_1414),
   .I2(gates_1198),
   .I3(gates_43),
   .I4(gates_1314),
   .I5(gates_1535)
);
LUT6 #(
   .INIT(64'b1111100011011110111101011010101010111101001001100000011011110011)  
) LUT6_1431 (
   .O(gates_528),
   .I0(gates_446),
   .I1(gates_1523),
   .I2(gates_336),
   .I3(gates_109),
   .I4(gates_433),
   .I5(gates_1121)
);
LUT6 #(
   .INIT(64'b0000011011001100100100111100110110100000101010100001110010110101)  
) LUT6_1432 (
   .O(gates_354),
   .I0(gates_994),
   .I1(gates_178),
   .I2(gates_691),
   .I3(gates_795),
   .I4(gates_697),
   .I5(gates_796)
);
LUT6 #(
   .INIT(64'b0010011010101101011010100011001011011100010001101001101101001100)  
) LUT6_1433 (
   .O(gates_92),
   .I0(gates_163),
   .I1(gates_513),
   .I2(gates_626),
   .I3(gates_355),
   .I4(gates_801),
   .I5(gates_1039)
);
LUT6 #(
   .INIT(64'b0000011011101011000010001111011010000111011110010011111011000000)  
) LUT6_1434 (
   .O(gates_1419),
   .I0(gates_94),
   .I1(gates_142),
   .I2(gates_6),
   .I3(gates_1448),
   .I4(gates_331),
   .I5(gates_930)
);
LUT6 #(
   .INIT(64'b1100111101010001100001111101110111011001011111000100010111011001)  
) LUT6_1435 (
   .O(gates_466),
   .I0(gates_206),
   .I1(gates_394),
   .I2(gates_1424),
   .I3(gates_1335),
   .I4(gates_1010),
   .I5(gates_430)
);
LUT6 #(
   .INIT(64'b0010110000001100010011111111111010100011100111111010011101000001)  
) LUT6_1436 (
   .O(gates_1050),
   .I0(gates_746),
   .I1(gates_694),
   .I2(gates_1516),
   .I3(gates_1122),
   .I4(gates_985),
   .I5(gates_497)
);
LUT6 #(
   .INIT(64'b1011100101101110111011011110110010000000110000111110101001111110)  
) LUT6_1437 (
   .O(gates_338),
   .I0(gates_1241),
   .I1(gates_469),
   .I2(gates_972),
   .I3(gates_257),
   .I4(gates_1193),
   .I5(gates_1017)
);
LUT6 #(
   .INIT(64'b1111000111000010110101000101010000110101001111001100001110111010)  
) LUT6_1438 (
   .O(gates_633),
   .I0(gates_15),
   .I1(gates_908),
   .I2(gates_182),
   .I3(gates_948),
   .I4(gates_822),
   .I5(gates_1506)
);
LUT6 #(
   .INIT(64'b0011010111010110000000011011010000101001011110111011101110110110)  
) LUT6_1439 (
   .O(gates_590),
   .I0(gates_465),
   .I1(gates_1430),
   .I2(gates_857),
   .I3(gates_448),
   .I4(gates_1106),
   .I5(gates_114)
);
LUT6 #(
   .INIT(64'b1110100110101001001101000110100000110110010101011010110101110001)  
) LUT6_1440 (
   .O(gates_1094),
   .I0(gates_1455),
   .I1(gates_98),
   .I2(gates_344),
   .I3(gates_241),
   .I4(gates_264),
   .I5(gates_1481)
);
LUT6 #(
   .INIT(64'b0101111100101110001100001101101101101000100111110011001000111010)  
) LUT6_1441 (
   .O(gates_540),
   .I0(gates_635),
   .I1(gates_1409),
   .I2(gates_872),
   .I3(gates_552),
   .I4(gates_24),
   .I5(gates_1528)
);
LUT6 #(
   .INIT(64'b1011110001110011100100100000010101100011100100110000001011110101)  
) LUT6_1442 (
   .O(gates_515),
   .I0(gates_310),
   .I1(gates_979),
   .I2(gates_533),
   .I3(gates_1143),
   .I4(gates_366),
   .I5(gates_1379)
);
LUT6 #(
   .INIT(64'b1011110011111110000101100101110001000011010011101011100111110000)  
) LUT6_1443 (
   .O(gates_529),
   .I0(gates_445),
   .I1(gates_919),
   .I2(gates_1404),
   .I3(gates_1123),
   .I4(gates_150),
   .I5(gates_939)
);
LUT6 #(
   .INIT(64'b0110101011111111100110111110111011101000010101011100011011001111)  
) LUT6_1444 (
   .O(gates_454),
   .I0(gates_1013),
   .I1(gates_1235),
   .I2(gates_1229),
   .I3(gates_1126),
   .I4(gates_1190),
   .I5(gates_300)
);
LUT6 #(
   .INIT(64'b1011001001111101001010000101000100101011010000101111011011100011)  
) LUT6_1445 (
   .O(gates_1501),
   .I0(gates_969),
   .I1(gates_696),
   .I2(gates_786),
   .I3(gates_318),
   .I4(gates_873),
   .I5(gates_741)
);
LUT6 #(
   .INIT(64'b1011001111001111001100101000100010001100101100111101111001011100)  
) LUT6_1446 (
   .O(gates_139),
   .I0(gates_1080),
   .I1(gates_521),
   .I2(gates_168),
   .I3(gates_1470),
   .I4(gates_1275),
   .I5(gates_1168)
);
LUT6 #(
   .INIT(64'b1100111111010011001011101010001000000010100101010100010000011010)  
) LUT6_1447 (
   .O(gates_1073),
   .I0(gates_688),
   .I1(gates_1480),
   .I2(gates_612),
   .I3(gates_245),
   .I4(gates_1413),
   .I5(gates_417)
);
LUT6 #(
   .INIT(64'b1001000001111011100100001011110010001111001001110110101001010111)  
) LUT6_1448 (
   .O(gates_623),
   .I0(gates_819),
   .I1(gates_692),
   .I2(gates_1088),
   .I3(gates_603),
   .I4(gates_473),
   .I5(gates_679)
);
LUT6 #(
   .INIT(64'b0001110010101011000100101101111110011100101010111001110001100001)  
) LUT6_1449 (
   .O(gates_1076),
   .I0(gates_1202),
   .I1(gates_809),
   .I2(gates_1187),
   .I3(gates_1274),
   .I4(gates_1484),
   .I5(gates_928)
);
LUT6 #(
   .INIT(64'b0110000100000001000011101000100000100100101100001001000101100111)  
) LUT6_1450 (
   .O(gates_49),
   .I0(gates_627),
   .I1(gates_1169),
   .I2(gates_1423),
   .I3(gates_1059),
   .I4(gates_358),
   .I5(gates_763)
);
LUT6 #(
   .INIT(64'b0010000100100111001100010111000100000100011010000001001000010010)  
) LUT6_1451 (
   .O(gates_285),
   .I0(gates_365),
   .I1(gates_773),
   .I2(gates_829),
   .I3(gates_734),
   .I4(gates_123),
   .I5(gates_75)
);
LUT6 #(
   .INIT(64'b1101011111111100100001010000010001011001101000111011111110111101)  
) LUT6_1452 (
   .O(gates_1234),
   .I0(gates_995),
   .I1(gates_253),
   .I2(gates_131),
   .I3(gates_1205),
   .I4(gates_1356),
   .I5(gates_1372)
);
LUT6 #(
   .INIT(64'b1010000000101011001001000100111000010000000011010101110000000111)  
) LUT6_1453 (
   .O(gates_502),
   .I0(gates_1497),
   .I1(gates_1439),
   .I2(gates_818),
   .I3(gates_1144),
   .I4(gates_184),
   .I5(gates_907)
);
LUT6 #(
   .INIT(64'b0010111011010010110001011100010000110101011001001000000001101000)  
) LUT6_1454 (
   .O(gates_803),
   .I0(gates_1486),
   .I1(gates_1336),
   .I2(gates_788),
   .I3(gates_771),
   .I4(gates_23),
   .I5(gates_1112)
);
LUT6 #(
   .INIT(64'b0111001001110010000110111100010101110000101010111110101101011111)  
) LUT6_1455 (
   .O(gates_1238),
   .I0(gates_1124),
   .I1(gates_1000),
   .I2(gates_875),
   .I3(gates_757),
   .I4(gates_817),
   .I5(gates_784)
);
LUT6 #(
   .INIT(64'b0001101111010101101111100000010011001010101111101001000001111000)  
) LUT6_1456 (
   .O(gates_54),
   .I0(gates_1023),
   .I1(gates_1460),
   .I2(gates_1386),
   .I3(gates_986),
   .I4(gates_89),
   .I5(gates_760)
);
LUT6 #(
   .INIT(64'b1001110011100001010010011000011110000010001000110011110000000101)  
) LUT6_1457 (
   .O(gates_551),
   .I0(gates_1429),
   .I1(gates_589),
   .I2(gates_878),
   .I3(gates_630),
   .I4(gates_1377),
   .I5(gates_360)
);
LUT6 #(
   .INIT(64'b0101111111110110010100010001000100001110111111101110110001011110)  
) LUT6_1458 (
   .O(gates_429),
   .I0(gates_1392),
   .I1(gates_1164),
   .I2(gates_534),
   .I3(gates_967),
   .I4(gates_1396),
   .I5(gates_1246)
);
LUT6 #(
   .INIT(64'b0010010010111101001001110100010011001100001110011000111111001010)  
) LUT6_1459 (
   .O(gates_865),
   .I0(gates_154),
   .I1(gates_1552),
   .I2(gates_1494),
   .I3(gates_1086),
   .I4(gates_674),
   .I5(gates_1524)
);
LUT6 #(
   .INIT(64'b1001111101110100110100110000111000000011100000011001010111010000)  
) LUT6_1460 (
   .O(gates_526),
   .I0(gates_615),
   .I1(gates_1149),
   .I2(gates_234),
   .I3(gates_1129),
   .I4(gates_1140),
   .I5(gates_1348)
);
LUT6 #(
   .INIT(64'b0011110101100000110100010101101010101011100011001110110010110101)  
) LUT6_1461 (
   .O(gates_1434),
   .I0(gates_44),
   .I1(gates_1378),
   .I2(gates_402),
   .I3(gates_325),
   .I4(gates_1456),
   .I5(gates_1453)
);
LUT6 #(
   .INIT(64'b1101100011100011011011111010100100100100000111000001110101010001)  
) LUT6_1462 (
   .O(gates_535),
   .I0(gates_1049),
   .I1(gates_965),
   .I2(gates_1218),
   .I3(gates_1107),
   .I4(gates_26),
   .I5(gates_911)
);
LUT6 #(
   .INIT(64'b0010100011100110110011010101001111011100001100111101111110101110)  
) LUT6_1463 (
   .O(gates_927),
   .I0(gates_749),
   .I1(gates_1),
   .I2(gates_543),
   .I3(gates_227),
   .I4(gates_321),
   .I5(gates_1322)
);
LUT6 #(
   .INIT(64'b1010001100000010011001101010101000000011011001110101010111101001)  
) LUT6_1464 (
   .O(gates_813),
   .I0(gates_482),
   .I1(gates_770),
   .I2(gates_492),
   .I3(gates_413),
   .I4(gates_1384),
   .I5(gates_438)
);
LUT6 #(
   .INIT(64'b1100010011000100110110001100100001111011111101011101111001111010)  
) LUT6_1465 (
   .O(gates_1103),
   .I0(gates_898),
   .I1(gates_1329),
   .I2(gates_146),
   .I3(gates_1321),
   .I4(gates_891),
   .I5(gates_1410)
);
LUT6 #(
   .INIT(64'b1101010110011000101111111110000111101100011000010100001101011000)  
) LUT6_1466 (
   .O(gates_33),
   .I0(gates_388),
   .I1(gates_1269),
   .I2(gates_954),
   .I3(gates_1323),
   .I4(gates_947),
   .I5(gates_950)
);
LUT6 #(
   .INIT(64'b1001101101101001100011011111110010001000011101000001000111011111)  
) LUT6_1467 (
   .O(gates_352),
   .I0(gates_900),
   .I1(gates_204),
   .I2(gates_1431),
   .I3(gates_846),
   .I4(gates_814),
   .I5(gates_370)
);
LUT6 #(
   .INIT(64'b1011001111111100111011001011101111101011111110100100011000010001)  
) LUT6_1468 (
   .O(gates_1016),
   .I0(gates_574),
   .I1(gates_272),
   .I2(gates_1224),
   .I3(gates_577),
   .I4(gates_237),
   .I5(gates_213)
);
LUT6 #(
   .INIT(64'b1001110100011100111001001010000011111101100100000000001111110100)  
) LUT6_1469 (
   .O(gates_602),
   .I0(gates_732),
   .I1(gates_1167),
   .I2(gates_1441),
   .I3(gates_120),
   .I4(gates_250),
   .I5(gates_1044)
);
LUT6 #(
   .INIT(64'b0001100100010001010100010100100101001100010000110011110000001001)  
) LUT6_1470 (
   .O(gates_931),
   .I0(gates_1426),
   .I1(gates_255),
   .I2(gates_190),
   .I3(gates_395),
   .I4(gates_1509),
   .I5(gates_807)
);
LUT6 #(
   .INIT(64'b1101100000010000001111001000101011110101100001110101100010010001)  
) LUT6_1471 (
   .O(gates_353),
   .I0(gates_1064),
   .I1(gates_235),
   .I2(gates_1142),
   .I3(gates_1491),
   .I4(gates_882),
   .I5(gates_712)
);
LUT6 #(
   .INIT(64'b1000111101100100011100001010110101101111001001011110100000011111)  
) LUT6_1472 (
   .O(gates_436),
   .I0(gates_532),
   .I1(gates_367),
   .I2(gates_170),
   .I3(gates_140),
   .I4(gates_179),
   .I5(gates_280)
);
LUT6 #(
   .INIT(64'b0101011111101000111001011111000111010011011010111100100010100110)  
) LUT6_1473 (
   .O(gates_1261),
   .I0(gates_65),
   .I1(gates_481),
   .I2(gates_1001),
   .I3(gates_638),
   .I4(gates_375),
   .I5(gates_855)
);
LUT6 #(
   .INIT(64'b0001110101000001100110110111100010111110000111010000001111101101)  
) LUT6_1474 (
   .O(gates_1371),
   .I0(gates_260),
   .I1(gates_1518),
   .I2(gates_859),
   .I3(gates_79),
   .I4(gates_1007),
   .I5(gates_495)
);
LUT6 #(
   .INIT(64'b1100101101111000001010001010001110000111111010100101110000111000)  
) LUT6_1475 (
   .O(gates_373),
   .I0(gates_718),
   .I1(gates_1022),
   .I2(gates_923),
   .I3(gates_1278),
   .I4(gates_361),
   .I5(gates_129)
);
LUT6 #(
   .INIT(64'b0000011000010100111100011100100000010110100010011100000010111010)  
) LUT6_1476 (
   .O(gates_764),
   .I0(gates_66),
   .I1(gates_657),
   .I2(gates_1184),
   .I3(gates_32),
   .I4(gates_653),
   .I5(gates_1008)
);
LUT6 #(
   .INIT(64'b0111001000111101011110000100101110111010000100110011111110000000)  
) LUT6_1477 (
   .O(gates_337),
   .I0(gates_453),
   .I1(gates_100),
   .I2(gates_36),
   .I3(gates_980),
   .I4(gates_614),
   .I5(gates_790)
);
LUT6 #(
   .INIT(64'b1111101101011101011011001011111001110111001011001001011000110110)  
) LUT6_1478 (
   .O(gates_837),
   .I0(gates_800),
   .I1(gates_278),
   .I2(gates_1345),
   .I3(gates_45),
   .I4(gates_1214),
   .I5(gates_38)
);
LUT6 #(
   .INIT(64'b1010011000100011001101100000001010010000001110001101110001100000)  
) LUT6_1479 (
   .O(gates_899),
   .I0(gates_399),
   .I1(gates_943),
   .I2(gates_1071),
   .I3(gates_820),
   .I4(gates_759),
   .I5(gates_1546)
);
LUT6 #(
   .INIT(64'b1000001011010111000011000111001011011111010111110111110100001100)  
) LUT6_1480 (
   .O(gates_1040),
   .I0(gates_1166),
   .I1(gates_1109),
   .I2(gates_509),
   .I3(gates_1374),
   .I4(gates_568),
   .I5(gates_743)
);
LUT6 #(
   .INIT(64'b1011001010000000111100011100011111001110001001000110011101011001)  
) LUT6_1481 (
   .O(gates_517),
   .I0(gates_753),
   .I1(gates_222),
   .I2(gates_393),
   .I3(gates_1019),
   .I4(gates_539),
   .I5(gates_451)
);
LUT6 #(
   .INIT(64'b0001001001110010111110100110111010101011111101100100101011101110)  
) LUT6_1482 (
   .O(gates_983),
   .I0(gates_1159),
   .I1(gates_689),
   .I2(gates_351),
   .I3(gates_133),
   .I4(gates_396),
   .I5(gates_1057)
);
LUT6 #(
   .INIT(64'b0101101000111001011110101111000010100000100111111000001101111110)  
) LUT6_1483 (
   .O(gates_1015),
   .I0(gates_1171),
   .I1(gates_996),
   .I2(gates_1350),
   .I3(gates_1236),
   .I4(gates_1037),
   .I5(gates_933)
);
LUT6 #(
   .INIT(64'b0011000100001110111001100000110111000110111100000000100010101001)  
) LUT6_1484 (
   .O(gates_439),
   .I0(gates_122),
   .I1(gates_1111),
   .I2(gates_598),
   .I3(gates_797),
   .I4(gates_220),
   .I5(gates_317)
);
LUT6 #(
   .INIT(64'b0111110010001001010111101001110110011110100011110110010010111101)  
) LUT6_1485 (
   .O(gates_221),
   .I0(gates_1300),
   .I1(gates_739),
   .I2(gates_307),
   .I3(gates_810),
   .I4(gates_970),
   .I5(gates_390)
);
LUT6 #(
   .INIT(64'b1111101001000011001000010101100110011001011101100001010100010110)  
) LUT6_1486 (
   .O(gates_754),
   .I0(gates_22),
   .I1(gates_591),
   .I2(gates_1194),
   .I3(gates_1492),
   .I4(gates_383),
   .I5(gates_778)
);
LUT6 #(
   .INIT(64'b1011010101110001011111000101100110111000111011001000000000010000)  
) LUT6_1487 (
   .O(gates_423),
   .I0(gates_496),
   .I1(gates_1197),
   .I2(gates_566),
   .I3(gates_11),
   .I4(gates_955),
   .I5(gates_1263)
);
LUT6 #(
   .INIT(64'b0001111101011110111100100000111100100001011101001101011000010111)  
) LUT6_1488 (
   .O(gates_883),
   .I0(gates_107),
   .I1(gates_1400),
   .I2(gates_1268),
   .I3(gates_664),
   .I4(gates_459),
   .I5(gates_169)
);
LUT6 #(
   .INIT(64'b1010011001110110111011101111000001001101110110001000000110011101)  
) LUT6_1489 (
   .O(gates_83),
   .I0(gates_424),
   .I1(gates_839),
   .I2(gates_1195),
   .I3(gates_617),
   .I4(gates_305),
   .I5(gates_756)
);
LUT6 #(
   .INIT(64'b1000000011000110000011011100011110100111001001101100101111011011)  
) LUT6_1490 (
   .O(gates_47),
   .I0(gates_1555),
   .I1(gates_1113),
   .I2(gates_1082),
   .I3(gates_597),
   .I4(gates_276),
   .I5(gates_463)
);
LUT6 #(
   .INIT(64'b1101101010001000101001110001100100100101101011001101111001001100)  
) LUT6_1491 (
   .O(gates_1333),
   .I0(gates_913),
   .I1(gates_484),
   .I2(gates_1365),
   .I3(gates_1021),
   .I4(gates_1310),
   .I5(gates_1331)
);
LUT6 #(
   .INIT(64'b1010110110000110010100001001110110101110010010000010010011110011)  
) LUT6_1492 (
   .O(gates_210),
   .I0(gates_1543),
   .I1(gates_705),
   .I2(gates_1154),
   .I3(gates_1258),
   .I4(gates_1373),
   .I5(gates_389)
);
LUT6 #(
   .INIT(64'b0100001001101010101111101010111001100101101111001110000001111100)  
) LUT6_1493 (
   .O(gates_101),
   .I0(gates_268),
   .I1(gates_584),
   .I2(gates_68),
   .I3(gates_1158),
   .I4(gates_1036),
   .I5(gates_328)
);
LUT6 #(
   .INIT(64'b0101010000110011010010111110110011111100100011011110000110110111)  
) LUT6_1494 (
   .O(gates_193),
   .I0(gates_201),
   .I1(gates_3),
   .I2(gates_30),
   .I3(gates_1062),
   .I4(gates_1538),
   .I5(gates_1069)
);
LUT6 #(
   .INIT(64'b1100001001010010101001100000001010010001010010110101000001010010)  
) LUT6_1495 (
   .O(gates_368),
   .I0(gates_1553),
   .I1(gates_1357),
   .I2(gates_151),
   .I3(gates_311),
   .I4(gates_849),
   .I5(gates_556)
);
LUT6 #(
   .INIT(64'b0011001111101100101100101111111001111010010100100001000010000110)  
) LUT6_1496 (
   .O(gates_158),
   .I0(gates_816),
   .I1(gates_1262),
   .I2(gates_832),
   .I3(gates_132),
   .I4(gates_1078),
   .I5(gates_1264)
);
LUT6 #(
   .INIT(64'b1101011001101101100110101100001111110000011101011000101100000110)  
) LUT6_1497 (
   .O(gates_714),
   .I0(gates_427),
   .I1(gates_641),
   .I2(gates_1273),
   .I3(gates_698),
   .I4(gates_1366),
   .I5(gates_1079)
);
LUT6 #(
   .INIT(64'b1101000011001001000011111101011001101111000111101101111101000101)  
) LUT6_1498 (
   .O(gates_348),
   .I0(gates_511),
   .I1(gates_1260),
   .I2(gates_999),
   .I3(gates_1151),
   .I4(gates_88),
   .I5(gates_642)
);
LUT6 #(
   .INIT(64'b1110101010101011101000101111001000110001000110100010001110001011)  
) LUT6_1499 (
   .O(gates_1351),
   .I0(gates_1511),
   .I1(gates_1075),
   .I2(gates_1280),
   .I3(gates_704),
   .I4(gates_812),
   .I5(gates_1196)
);
LUT6 #(
   .INIT(64'b0110011101001101110111110110100101111001000100000101011001101110)  
) LUT6_1500 (
   .O(gates_716),
   .I0(gates_887),
   .I1(gates_783),
   .I2(gates_1152),
   .I3(gates_830),
   .I4(gates_288),
   .I5(gates_1189)
);
LUT6 #(
   .INIT(64'b0000011010010100111110100001001101110010110010010000110011001110)  
) LUT6_1501 (
   .O(gates_77),
   .I0(gates_372),
   .I1(gates_827),
   .I2(gates_1287),
   .I3(gates_73),
   .I4(gates_909),
   .I5(gates_1004)
);
LUT6 #(
   .INIT(64'b0110010110100001010000001000110011110110010100000011111100111001)  
) LUT6_1502 (
   .O(gates_1531),
   .I0(gates_988),
   .I1(gates_596),
   .I2(gates_974),
   .I3(gates_419),
   .I4(gates_774),
   .I5(gates_1407)
);
LUT6 #(
   .INIT(64'b1011111100010011101100110100110101111000100101011111001100001010)  
) LUT6_1503 (
   .O(gates_1520),
   .I0(gates_629),
   .I1(gates_661),
   .I2(gates_286),
   .I3(gates_476),
   .I4(gates_605),
   .I5(gates_1041)
);
LUT6 #(
   .INIT(64'b0100000110111011011011000101001010111101100100101001000100101110)  
) LUT6_1504 (
   .O(gates_1281),
   .I0(gates_894),
   .I1(gates_1095),
   .I2(gates_236),
   .I3(gates_1307),
   .I4(gates_646),
   .I5(gates_772)
);
LUT6 #(
   .INIT(64'b1110000101111110101010010110100100001111000101011110000001010000)  
) LUT6_1505 (
   .O(gates_992),
   .I0(gates_1108),
   .I1(gates_706),
   .I2(gates_1437),
   .I3(gates_364),
   .I4(gates_1483),
   .I5(gates_1093)
);
LUT6 #(
   .INIT(64'b1100110010010111111111101000000000011110010110000011101000000100)  
) LUT6_1506 (
   .O(gates_51),
   .I0(gates_1519),
   .I1(gates_197),
   .I2(gates_791),
   .I3(gates_508),
   .I4(gates_921),
   .I5(gates_215)
);
LUT6 #(
   .INIT(64'b0001110000010111101000001111100111111011010101010000101010000110)  
) LUT6_1507 (
   .O(gates_458),
   .I0(gates_259),
   .I1(gates_301),
   .I2(gates_1243),
   .I3(gates_811),
   .I4(gates_1395),
   .I5(gates_483)
);
LUT6 #(
   .INIT(64'b1111101000100000100010011001100111100010111010001111100010000101)  
) LUT6_1508 (
   .O(gates_1024),
   .I0(gates_538),
   .I1(gates_1398),
   .I2(gates_21),
   .I3(gates_97),
   .I4(gates_963),
   .I5(gates_191)
);
LUT6 #(
   .INIT(64'b1010000101001001110011001010010010001111000110100000011101010111)  
) LUT6_1509 (
   .O(gates_546),
   .I0(gates_876),
   .I1(gates_506),
   .I2(gates_1020),
   .I3(gates_1510),
   .I4(gates_162),
   .I5(gates_52)
);
LUT6 #(
   .INIT(64'b1001111001111110101001000011011110111111100000100011110111010000)  
) LUT6_1510 (
   .O(gates_903),
   .I0(gates_267),
   .I1(gates_724),
   .I2(gates_621),
   .I3(gates_717),
   .I4(gates_194),
   .I5(gates_302)
);
LUT6 #(
   .INIT(64'b1011101011001100110010111111000001010010111110111010011010010010)  
) LUT6_1511 (
   .O(gates_558),
   .I0(gates_1006),
   .I1(gates_379),
   .I2(gates_834),
   .I3(gates_125),
   .I4(gates_545),
   .I5(gates_74)
);
LUT6 #(
   .INIT(64'b1101100011000111111000001111100111010011100111000010111101011001)  
) LUT6_1512 (
   .O(gates_134),
   .I0(gates_82),
   .I1(gates_557),
   .I2(gates_292),
   .I3(gates_1085),
   .I4(gates_1554),
   .I5(gates_654)
);
LUT6 #(
   .INIT(64'b0100000000101001110110110001101110011101110111100000110101000110)  
) LUT6_1513 (
   .O(gates_1035),
   .I0(gates_720),
   .I1(gates_733),
   .I2(gates_644),
   .I3(gates_216),
   .I4(gates_1150),
   .I5(gates_81)
);
LUT6 #(
   .INIT(64'b1001100111101001101111110001110100100100100111010101111111011011)  
) LUT6_1514 (
   .O(gates_91),
   .I0(gates_199),
   .I1(gates_447),
   .I2(gates_1217),
   .I3(gates_346),
   .I4(gates_130),
   .I5(gates_31)
);
LUT6 #(
   .INIT(64'b0101100110011000001111010010010000000100100011001010011000100001)  
) LUT6_1515 (
   .O(gates_1505),
   .I0(gates_1061),
   .I1(gates_1031),
   .I2(gates_410),
   .I3(gates_562),
   .I4(gates_853),
   .I5(gates_1110)
);
LUT6 #(
   .INIT(64'b1001001100001001001001011001100000100100011011010010111101101011)  
) LUT6_1516 (
   .O(gates_452),
   .I0(gates_1068),
   .I1(gates_1131),
   .I2(gates_110),
   .I3(gates_929),
   .I4(gates_218),
   .I5(gates_1339)
);
LUT6 #(
   .INIT(64'b0110000011010111111001000100010010000100001010010110001111101010)  
) LUT6_1517 (
   .O(gates_1488),
   .I0(gates_920),
   .I1(gates_1132),
   .I2(gates_628),
   .I3(gates_1114),
   .I4(gates_1067),
   .I5(gates_601)
);
LUT6 #(
   .INIT(64'b1111111001110001011111000101000100001110111110001001011101010001)  
) LUT6_1518 (
   .O(gates_576),
   .I0(gates_266),
   .I1(gates_1257),
   .I2(gates_500),
   .I3(gates_1408),
   .I4(gates_946),
   .I5(gates_1012)
);
LUT6 #(
   .INIT(64'b1001111100110001100100101001010101101101001110100011110110011011)  
) LUT6_1519 (
   .O(gates_1542),
   .I0(gates_789),
   .I1(gates_258),
   .I2(gates_1525),
   .I3(gates_271),
   .I4(gates_731),
   .I5(gates_663)
);
LUT6 #(
   .INIT(64'b0010101110000001110011100000011110111100010110111010110001010000)  
) LUT6_1520 (
   .O(gates_779),
   .I0(gates_1221),
   .I1(gates_964),
   .I2(gates_174),
   .I3(gates_802),
   .I4(gates_845),
   .I5(gates_104)
);
LUT6 #(
   .INIT(64'b1111100000100011110010001011101000010110000100110100001101000101)  
) LUT6_1521 (
   .O(gates_1155),
   .I0(gates_10),
   .I1(gates_398),
   .I2(gates_573),
   .I3(gates_486),
   .I4(gates_1442),
   .I5(gates_737)
);
LUT6 #(
   .INIT(64'b1101010101010000100001001111110111110011110011101100000110011010)  
) LUT6_1522 (
   .O(gates_1097),
   .I0(gates_1162),
   .I1(gates_1368),
   .I2(gates_1253),
   .I3(gates_53),
   .I4(gates_1014),
   .I5(gates_1513)
);
LUT6 #(
   .INIT(64'b1110000010000010111100011011111000001110101011001001110111000010)  
) LUT6_1523 (
   .O(gates_658),
   .I0(gates_1319),
   .I1(gates_472),
   .I2(gates_910),
   .I3(gates_604),
   .I4(gates_71),
   .I5(gates_219)
);
LUT6 #(
   .INIT(64'b1101011111110001010110110000100001111011111111001011101110101010)  
) LUT6_1524 (
   .O(gates_525),
   .I0(gates_1301),
   .I1(gates_1521),
   .I2(gates_397),
   .I3(gates_707),
   .I4(gates_1227),
   .I5(gates_925)
);
LUT6 #(
   .INIT(64'b0111100110001110011000100011101011100010100101010000011010010100)  
) LUT6_1525 (
   .O(gates_956),
   .I0(gates_1047),
   .I1(gates_662),
   .I2(gates_684),
   .I3(gates_1179),
   .I4(gates_1117),
   .I5(gates_407)
);
LUT6 #(
   .INIT(64'b0000100100001101011001000110111110001101100111011110111111000110)  
) LUT6_1526 (
   .O(gates_1475),
   .I0(gates_794),
   .I1(gates_991),
   .I2(gates_593),
   .I3(gates_821),
   .I4(gates_1471),
   .I5(gates_634)
);
LUT6 #(
   .INIT(64'b0111101100111111011111010001100000000000000111110100111000001011)  
) LUT6_1527 (
   .O(gates_856),
   .I0(gates_434),
   .I1(gates_1216),
   .I2(gates_1141),
   .I3(gates_339),
   .I4(gates_418),
   .I5(gates_751)
);
LUT6 #(
   .INIT(64'b0001110101110101111111110101000001101001111011111111010110011100)  
) LUT6_1528 (
   .O(gates_976),
   .I0(gates_685),
   .I1(gates_1011),
   .I2(gates_776),
   .I3(gates_202),
   .I4(gates_599),
   .I5(gates_475)
);
LUT6 #(
   .INIT(64'b0010111010000100101110000001111110110110100000000011011000111100)  
) LUT6_1529 (
   .O(gates_1265),
   .I0(gates_347),
   .I1(gates_295),
   .I2(gates_1452),
   .I3(gates_594),
   .I4(gates_619),
   .I5(gates_1454)
);
LUT6 #(
   .INIT(64'b1111000000110010000000101100011000000010010011010100110111101001)  
) LUT6_1530 (
   .O(gates_1544),
   .I0(gates_868),
   .I1(gates_559),
   .I2(gates_1174),
   .I3(gates_1254),
   .I4(gates_564),
   .I5(gates_787)
);
LUT6 #(
   .INIT(64'b1100011000011100000001101000010110000111001111011000001011011010)  
) LUT6_1531 (
   .O(gates_1283),
   .I0(gates_742),
   .I1(gates_877),
   .I2(gates_232),
   .I3(gates_695),
   .I4(gates_918),
   .I5(gates_1055)
);
LUT6 #(
   .INIT(64'b1110111111111010100001000111111001001110001100000100011011110010)  
) LUT6_1532 (
   .O(gates_1363),
   .I0(gates_400),
   .I1(gates_1311),
   .I2(gates_284),
   .I3(gates_211),
   .I4(gates_296),
   .I5(gates_611)
);
LUT6 #(
   .INIT(64'b1000001000101000100000110000000001111111000101101000100100101001)  
) LUT6_1533 (
   .O(gates_915),
   .I0(gates_660),
   .I1(gates_1487),
   .I2(gates_1515),
   .I3(gates_777),
   .I4(gates_755),
   .I5(gates_67)
);
LUT6 #(
   .INIT(64'b1110111100100110001111011100010110110000011111011011000111001010)  
) LUT6_1534 (
   .O(gates_843),
   .I0(gates_989),
   .I1(gates_1191),
   .I2(gates_650),
   .I3(gates_758),
   .I4(gates_524),
   .I5(gates_1276)
);
LUT6 #(
   .INIT(64'b0010000101010011000000000110111100111110101100011010011011001010)  
) LUT6_1535 (
   .O(gates_273),
   .I0(gates_1419),
   .I1(gates_92),
   .I2(gates_354),
   .I3(gates_528),
   .I4(gates_431),
   .I5(gates_645)
);
LUT6 #(
   .INIT(64'b1001010101010001111110111011001101110100001001011111010011100000)  
) LUT6_1536 (
   .O(gates_242),
   .I0(gates_1094),
   .I1(gates_590),
   .I2(gates_633),
   .I3(gates_338),
   .I4(gates_1050),
   .I5(gates_466)
);
LUT6 #(
   .INIT(64'b0000100011100011100011011101010100001000100100001110011100101001)  
) LUT6_1537 (
   .O(gates_1244),
   .I0(gates_139),
   .I1(gates_1501),
   .I2(gates_454),
   .I3(gates_529),
   .I4(gates_515),
   .I5(gates_540)
);
LUT6 #(
   .INIT(64'b1111010000000101011010111010000000000001110010111100011100101010)  
) LUT6_1538 (
   .O(gates_637),
   .I0(gates_1234),
   .I1(gates_285),
   .I2(gates_49),
   .I3(gates_1076),
   .I4(gates_623),
   .I5(gates_1073)
);
LUT6 #(
   .INIT(64'b1101111011001101000100111011100110100001111111001111011000001001)  
) LUT6_1539 (
   .O(gates_721),
   .I0(gates_429),
   .I1(gates_551),
   .I2(gates_54),
   .I3(gates_1238),
   .I4(gates_803),
   .I5(gates_502)
);
LUT6 #(
   .INIT(64'b0010110011110100110010101111111100100101001111100111010101111110)  
) LUT6_1540 (
   .O(gates_18),
   .I0(gates_813),
   .I1(gates_927),
   .I2(gates_535),
   .I3(gates_1434),
   .I4(gates_526),
   .I5(gates_865)
);
LUT6 #(
   .INIT(64'b1010001001001001011110101011001111101101101011000101011001010111)  
) LUT6_1541 (
   .O(gates_958),
   .I0(gates_931),
   .I1(gates_602),
   .I2(gates_1016),
   .I3(gates_352),
   .I4(gates_33),
   .I5(gates_1103)
);
LUT6 #(
   .INIT(64'b0110101010110010111100111100110111101000001011011000011111110100)  
) LUT6_1542 (
   .O(gates_113),
   .I0(gates_764),
   .I1(gates_373),
   .I2(gates_1371),
   .I3(gates_1261),
   .I4(gates_436),
   .I5(gates_353)
);
LUT6 #(
   .INIT(64'b1001010101110110011000101101010001111001100101001010011010111011)  
) LUT6_1543 (
   .O(gates_1025),
   .I0(gates_983),
   .I1(gates_517),
   .I2(gates_1040),
   .I3(gates_899),
   .I4(gates_837),
   .I5(gates_337)
);
LUT6 #(
   .INIT(64'b0101101000000111111001111011011110011001110101101000111101100111)  
) LUT6_1544 (
   .O(gates_1291),
   .I0(gates_883),
   .I1(gates_423),
   .I2(gates_754),
   .I3(gates_221),
   .I4(gates_439),
   .I5(gates_1015)
);
LUT6 #(
   .INIT(64'b0000000101101100100100010110110001010110000101110011011101110100)  
) LUT6_1545 (
   .O(gates_1428),
   .I0(gates_193),
   .I1(gates_101),
   .I2(gates_210),
   .I3(gates_1333),
   .I4(gates_47),
   .I5(gates_83)
);
LUT6 #(
   .INIT(64'b1100100000011100111101001011010000000000110110111101111100000001)  
) LUT6_1546 (
   .O(gates_1540),
   .I0(gates_716),
   .I1(gates_1351),
   .I2(gates_348),
   .I3(gates_714),
   .I4(gates_158),
   .I5(gates_368)
);
LUT6 #(
   .INIT(64'b1011100111001110001010011011100010110011100100101010101101111001)  
) LUT6_1547 (
   .O(gates_1533),
   .I0(gates_51),
   .I1(gates_992),
   .I2(gates_1281),
   .I3(gates_1520),
   .I4(gates_1531),
   .I5(gates_77)
);
LUT6 #(
   .INIT(64'b1001001110111110001101001100010010010000101100000000100101011101)  
) LUT6_1548 (
   .O(gates_312),
   .I0(gates_134),
   .I1(gates_558),
   .I2(gates_903),
   .I3(gates_546),
   .I4(gates_1024),
   .I5(gates_458)
);
LUT6 #(
   .INIT(64'b0100010011101011011100011000010110011000110011110100001010011111)  
) LUT6_1549 (
   .O(gates_39),
   .I0(gates_576),
   .I1(gates_1488),
   .I2(gates_452),
   .I3(gates_1505),
   .I4(gates_91),
   .I5(gates_1035)
);
LUT6 #(
   .INIT(64'b1101011100101100111101111100101000011011100111001000101111101000)  
) LUT6_1550 (
   .O(gates_860),
   .I0(gates_525),
   .I1(gates_658),
   .I2(gates_1097),
   .I3(gates_1155),
   .I4(gates_779),
   .I5(gates_1542)
);
LUT6 #(
   .INIT(64'b0110001100101000000010010101001100100100000110101110101001010111)  
) LUT6_1551 (
   .O(gates_138),
   .I0(gates_1544),
   .I1(gates_1265),
   .I2(gates_976),
   .I3(gates_856),
   .I4(gates_1475),
   .I5(gates_956)
);
LUT6 #(
   .INIT(64'b0111101100101111101100000010110011100100110101010101111111111010)  
) LUT6_1552 (
   .O(gates_981),
   .I0(gates_242),
   .I1(gates_273),
   .I2(gates_843),
   .I3(gates_915),
   .I4(gates_1363),
   .I5(gates_1283)
);
LUT6 #(
   .INIT(64'b1001001111111010001101011010100111010000010100110101010101001000)  
) LUT6_1553 (
   .O(gates_1256),
   .I0(gates_113),
   .I1(gates_958),
   .I2(gates_18),
   .I3(gates_721),
   .I4(gates_637),
   .I5(gates_1244)
);
LUT6 #(
   .INIT(64'b0110000000100110001100001011011101101111111100000010111011010001)  
) LUT6_1554 (
   .O(gates_175),
   .I0(gates_312),
   .I1(gates_1533),
   .I2(gates_1540),
   .I3(gates_1428),
   .I4(gates_1291),
   .I5(gates_1025)
);
LUT6 #(
   .INIT(64'b1000001100101011100110110111011011000101001110001100011101000101)  
) LUT6_1555 (
   .O(gates_1422),
   .I0(gates_175),
   .I1(gates_1256),
   .I2(gates_981),
   .I3(gates_138),
   .I4(gates_860),
   .I5(gates_39)
);



endmodule